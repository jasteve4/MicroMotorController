magic
tech gf180mcuC
magscale 1 5
timestamp 1670300988
<< obsm1 >>
rect 672 1538 89320 70198
<< metal2 >>
rect 2128 0 2184 400
rect 4032 0 4088 400
rect 5936 0 5992 400
rect 7840 0 7896 400
rect 9744 0 9800 400
rect 11648 0 11704 400
rect 13552 0 13608 400
rect 15456 0 15512 400
rect 17360 0 17416 400
rect 19264 0 19320 400
rect 21168 0 21224 400
rect 23072 0 23128 400
rect 24976 0 25032 400
rect 26880 0 26936 400
rect 28784 0 28840 400
rect 30688 0 30744 400
rect 32592 0 32648 400
rect 34496 0 34552 400
rect 36400 0 36456 400
rect 38304 0 38360 400
rect 40208 0 40264 400
rect 42112 0 42168 400
rect 44016 0 44072 400
rect 45920 0 45976 400
rect 47824 0 47880 400
rect 49728 0 49784 400
rect 51632 0 51688 400
rect 53536 0 53592 400
rect 55440 0 55496 400
rect 57344 0 57400 400
rect 59248 0 59304 400
rect 61152 0 61208 400
rect 63056 0 63112 400
rect 64960 0 65016 400
rect 66864 0 66920 400
rect 68768 0 68824 400
rect 70672 0 70728 400
rect 72576 0 72632 400
rect 74480 0 74536 400
rect 76384 0 76440 400
rect 78288 0 78344 400
rect 80192 0 80248 400
rect 82096 0 82152 400
rect 84000 0 84056 400
rect 85904 0 85960 400
rect 87808 0 87864 400
<< obsm2 >>
rect 798 430 89474 70187
rect 798 289 2098 430
rect 2214 289 4002 430
rect 4118 289 5906 430
rect 6022 289 7810 430
rect 7926 289 9714 430
rect 9830 289 11618 430
rect 11734 289 13522 430
rect 13638 289 15426 430
rect 15542 289 17330 430
rect 17446 289 19234 430
rect 19350 289 21138 430
rect 21254 289 23042 430
rect 23158 289 24946 430
rect 25062 289 26850 430
rect 26966 289 28754 430
rect 28870 289 30658 430
rect 30774 289 32562 430
rect 32678 289 34466 430
rect 34582 289 36370 430
rect 36486 289 38274 430
rect 38390 289 40178 430
rect 40294 289 42082 430
rect 42198 289 43986 430
rect 44102 289 45890 430
rect 46006 289 47794 430
rect 47910 289 49698 430
rect 49814 289 51602 430
rect 51718 289 53506 430
rect 53622 289 55410 430
rect 55526 289 57314 430
rect 57430 289 59218 430
rect 59334 289 61122 430
rect 61238 289 63026 430
rect 63142 289 64930 430
rect 65046 289 66834 430
rect 66950 289 68738 430
rect 68854 289 70642 430
rect 70758 289 72546 430
rect 72662 289 74450 430
rect 74566 289 76354 430
rect 76470 289 78258 430
rect 78374 289 80162 430
rect 80278 289 82066 430
rect 82182 289 83970 430
rect 84086 289 85874 430
rect 85990 289 87778 430
rect 87894 289 89474 430
<< obsm3 >>
rect 793 294 89479 70182
<< metal4 >>
rect 1092 1538 1252 70198
rect 5592 1538 5752 70198
rect 10092 1538 10252 70198
rect 14592 1538 14752 70198
rect 19092 1538 19252 70198
rect 23592 1538 23752 70198
rect 28092 1538 28252 70198
rect 32592 1538 32752 70198
rect 37092 1538 37252 70198
rect 41592 1538 41752 70198
rect 46092 1538 46252 70198
rect 50592 1538 50752 70198
rect 55092 1538 55252 70198
rect 59592 1538 59752 70198
rect 64092 1538 64252 70198
rect 68592 1538 68752 70198
rect 73092 1538 73252 70198
rect 77592 1538 77752 70198
rect 82092 1538 82252 70198
rect 86592 1538 86752 70198
<< obsm4 >>
rect 5502 1508 5562 68143
rect 5782 1508 10062 68143
rect 10282 1508 14562 68143
rect 14782 1508 19062 68143
rect 19282 1508 23562 68143
rect 23782 1508 28062 68143
rect 28282 1508 32562 68143
rect 32782 1508 37062 68143
rect 37282 1508 41562 68143
rect 41782 1508 46062 68143
rect 46282 1508 50562 68143
rect 50782 1508 55062 68143
rect 55282 1508 59562 68143
rect 59782 1508 64062 68143
rect 64282 1508 68562 68143
rect 68782 1508 73062 68143
rect 73282 1508 77562 68143
rect 77782 1508 82062 68143
rect 82282 1508 86562 68143
rect 86782 1508 88466 68143
rect 5502 457 88466 1508
<< labels >>
rlabel metal2 s 68768 0 68824 400 6 clock
port 1 nsew signal input
rlabel metal2 s 70672 0 70728 400 6 clock_a
port 2 nsew signal input
rlabel metal2 s 57344 0 57400 400 6 col_select_a[0]
port 3 nsew signal input
rlabel metal2 s 59248 0 59304 400 6 col_select_a[1]
port 4 nsew signal input
rlabel metal2 s 61152 0 61208 400 6 col_select_a[2]
port 5 nsew signal input
rlabel metal2 s 63056 0 63112 400 6 col_select_a[3]
port 6 nsew signal input
rlabel metal2 s 64960 0 65016 400 6 col_select_a[4]
port 7 nsew signal input
rlabel metal2 s 66864 0 66920 400 6 col_select_a[5]
port 8 nsew signal input
rlabel metal2 s 5936 0 5992 400 6 data_in_a[0]
port 9 nsew signal input
rlabel metal2 s 24976 0 25032 400 6 data_in_a[10]
port 10 nsew signal input
rlabel metal2 s 26880 0 26936 400 6 data_in_a[11]
port 11 nsew signal input
rlabel metal2 s 28784 0 28840 400 6 data_in_a[12]
port 12 nsew signal input
rlabel metal2 s 30688 0 30744 400 6 data_in_a[13]
port 13 nsew signal input
rlabel metal2 s 32592 0 32648 400 6 data_in_a[14]
port 14 nsew signal input
rlabel metal2 s 34496 0 34552 400 6 data_in_a[15]
port 15 nsew signal input
rlabel metal2 s 7840 0 7896 400 6 data_in_a[1]
port 16 nsew signal input
rlabel metal2 s 9744 0 9800 400 6 data_in_a[2]
port 17 nsew signal input
rlabel metal2 s 11648 0 11704 400 6 data_in_a[3]
port 18 nsew signal input
rlabel metal2 s 13552 0 13608 400 6 data_in_a[4]
port 19 nsew signal input
rlabel metal2 s 15456 0 15512 400 6 data_in_a[5]
port 20 nsew signal input
rlabel metal2 s 17360 0 17416 400 6 data_in_a[6]
port 21 nsew signal input
rlabel metal2 s 19264 0 19320 400 6 data_in_a[7]
port 22 nsew signal input
rlabel metal2 s 21168 0 21224 400 6 data_in_a[8]
port 23 nsew signal input
rlabel metal2 s 23072 0 23128 400 6 data_in_a[9]
port 24 nsew signal input
rlabel metal2 s 2128 0 2184 400 6 driver_io[0]
port 25 nsew signal output
rlabel metal2 s 4032 0 4088 400 6 driver_io[1]
port 26 nsew signal output
rlabel metal2 s 87808 0 87864 400 6 inverter_select_a
port 27 nsew signal input
rlabel metal2 s 36400 0 36456 400 6 mem_address_a[0]
port 28 nsew signal input
rlabel metal2 s 38304 0 38360 400 6 mem_address_a[1]
port 29 nsew signal input
rlabel metal2 s 40208 0 40264 400 6 mem_address_a[2]
port 30 nsew signal input
rlabel metal2 s 42112 0 42168 400 6 mem_address_a[3]
port 31 nsew signal input
rlabel metal2 s 44016 0 44072 400 6 mem_address_a[4]
port 32 nsew signal input
rlabel metal2 s 45920 0 45976 400 6 mem_address_a[5]
port 33 nsew signal input
rlabel metal2 s 47824 0 47880 400 6 mem_address_a[6]
port 34 nsew signal input
rlabel metal2 s 49728 0 49784 400 6 mem_address_a[7]
port 35 nsew signal input
rlabel metal2 s 51632 0 51688 400 6 mem_address_a[8]
port 36 nsew signal input
rlabel metal2 s 53536 0 53592 400 6 mem_address_a[9]
port 37 nsew signal input
rlabel metal2 s 55440 0 55496 400 6 mem_write_n_a
port 38 nsew signal input
rlabel metal2 s 85904 0 85960 400 6 output_active_a
port 39 nsew signal input
rlabel metal2 s 84000 0 84056 400 6 row_col_select_a
port 40 nsew signal input
rlabel metal2 s 72576 0 72632 400 6 row_select_a[0]
port 41 nsew signal input
rlabel metal2 s 74480 0 74536 400 6 row_select_a[1]
port 42 nsew signal input
rlabel metal2 s 76384 0 76440 400 6 row_select_a[2]
port 43 nsew signal input
rlabel metal2 s 78288 0 78344 400 6 row_select_a[3]
port 44 nsew signal input
rlabel metal2 s 80192 0 80248 400 6 row_select_a[4]
port 45 nsew signal input
rlabel metal2 s 82096 0 82152 400 6 row_select_a[5]
port 46 nsew signal input
rlabel metal4 s 1092 1538 1252 70198 6 vdd
port 47 nsew power bidirectional
rlabel metal4 s 10092 1538 10252 70198 6 vdd
port 47 nsew power bidirectional
rlabel metal4 s 19092 1538 19252 70198 6 vdd
port 47 nsew power bidirectional
rlabel metal4 s 28092 1538 28252 70198 6 vdd
port 47 nsew power bidirectional
rlabel metal4 s 37092 1538 37252 70198 6 vdd
port 47 nsew power bidirectional
rlabel metal4 s 46092 1538 46252 70198 6 vdd
port 47 nsew power bidirectional
rlabel metal4 s 55092 1538 55252 70198 6 vdd
port 47 nsew power bidirectional
rlabel metal4 s 64092 1538 64252 70198 6 vdd
port 47 nsew power bidirectional
rlabel metal4 s 73092 1538 73252 70198 6 vdd
port 47 nsew power bidirectional
rlabel metal4 s 82092 1538 82252 70198 6 vdd
port 47 nsew power bidirectional
rlabel metal4 s 5592 1538 5752 70198 6 vss
port 48 nsew ground bidirectional
rlabel metal4 s 14592 1538 14752 70198 6 vss
port 48 nsew ground bidirectional
rlabel metal4 s 23592 1538 23752 70198 6 vss
port 48 nsew ground bidirectional
rlabel metal4 s 32592 1538 32752 70198 6 vss
port 48 nsew ground bidirectional
rlabel metal4 s 41592 1538 41752 70198 6 vss
port 48 nsew ground bidirectional
rlabel metal4 s 50592 1538 50752 70198 6 vss
port 48 nsew ground bidirectional
rlabel metal4 s 59592 1538 59752 70198 6 vss
port 48 nsew ground bidirectional
rlabel metal4 s 68592 1538 68752 70198 6 vss
port 48 nsew ground bidirectional
rlabel metal4 s 77592 1538 77752 70198 6 vss
port 48 nsew ground bidirectional
rlabel metal4 s 86592 1538 86752 70198 6 vss
port 48 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 90000 72000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 17958882
string GDS_FILE /home/jasteve4/Documents/MicroMotorController/openlane/driver_core/runs/22_12_05_23_26/results/signoff/driver_core.magic.gds
string GDS_START 274444
<< end >>


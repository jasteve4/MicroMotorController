magic
tech gf180mcuC
magscale 1 5
timestamp 1670279604
<< obsm1 >>
rect 672 1538 89320 70198
<< metal2 >>
rect 2100 -480 2212 240
rect 4004 -480 4116 240
rect 5908 -480 6020 240
rect 7812 -480 7924 240
rect 9716 -480 9828 240
rect 11620 -480 11732 240
rect 13524 -480 13636 240
rect 15428 -480 15540 240
rect 17332 -480 17444 240
rect 19236 -480 19348 240
rect 21140 -480 21252 240
rect 23044 -480 23156 240
rect 24948 -480 25060 240
rect 26852 -480 26964 240
rect 28756 -480 28868 240
rect 30660 -480 30772 240
rect 32564 -480 32676 240
rect 34468 -480 34580 240
rect 36372 -480 36484 240
rect 38276 -480 38388 240
rect 40180 -480 40292 240
rect 42084 -480 42196 240
rect 43988 -480 44100 240
rect 45892 -480 46004 240
rect 47796 -480 47908 240
rect 49700 -480 49812 240
rect 51604 -480 51716 240
rect 53508 -480 53620 240
rect 55412 -480 55524 240
rect 57316 -480 57428 240
rect 59220 -480 59332 240
rect 61124 -480 61236 240
rect 63028 -480 63140 240
rect 64932 -480 65044 240
rect 66836 -480 66948 240
rect 68740 -480 68852 240
rect 70644 -480 70756 240
rect 72548 -480 72660 240
rect 74452 -480 74564 240
rect 76356 -480 76468 240
rect 78260 -480 78372 240
rect 80164 -480 80276 240
rect 82068 -480 82180 240
rect 83972 -480 84084 240
rect 85876 -480 85988 240
rect 87780 -480 87892 240
<< obsm2 >>
rect 966 270 89194 70187
rect 966 177 2070 270
rect 2242 177 3974 270
rect 4146 177 5878 270
rect 6050 177 7782 270
rect 7954 177 9686 270
rect 9858 177 11590 270
rect 11762 177 13494 270
rect 13666 177 15398 270
rect 15570 177 17302 270
rect 17474 177 19206 270
rect 19378 177 21110 270
rect 21282 177 23014 270
rect 23186 177 24918 270
rect 25090 177 26822 270
rect 26994 177 28726 270
rect 28898 177 30630 270
rect 30802 177 32534 270
rect 32706 177 34438 270
rect 34610 177 36342 270
rect 36514 177 38246 270
rect 38418 177 40150 270
rect 40322 177 42054 270
rect 42226 177 43958 270
rect 44130 177 45862 270
rect 46034 177 47766 270
rect 47938 177 49670 270
rect 49842 177 51574 270
rect 51746 177 53478 270
rect 53650 177 55382 270
rect 55554 177 57286 270
rect 57458 177 59190 270
rect 59362 177 61094 270
rect 61266 177 62998 270
rect 63170 177 64902 270
rect 65074 177 66806 270
rect 66978 177 68710 270
rect 68882 177 70614 270
rect 70786 177 72518 270
rect 72690 177 74422 270
rect 74594 177 76326 270
rect 76498 177 78230 270
rect 78402 177 80134 270
rect 80306 177 82038 270
rect 82210 177 83942 270
rect 84114 177 85846 270
rect 86018 177 87750 270
rect 87922 177 89194 270
<< obsm3 >>
rect 961 182 89199 70182
<< metal4 >>
rect 1017 1538 1327 70198
rect 2877 1538 3187 70198
rect 19017 1538 19327 70198
rect 20877 1538 21187 70198
rect 37017 1538 37327 70198
rect 38877 1538 39187 70198
rect 55017 1538 55327 70198
rect 56877 1538 57187 70198
rect 73017 1538 73327 70198
rect 74877 1538 75187 70198
<< obsm4 >>
rect 3262 1508 18987 65959
rect 19357 1508 20847 65959
rect 21217 1508 36987 65959
rect 37357 1508 38847 65959
rect 39217 1508 54987 65959
rect 55357 1508 56847 65959
rect 57217 1508 72987 65959
rect 73357 1508 74847 65959
rect 75217 1508 86562 65959
rect 3262 457 86562 1508
<< labels >>
rlabel metal2 s 68740 -480 68852 240 8 clock
port 1 nsew signal input
rlabel metal2 s 70644 -480 70756 240 8 clock_a
port 2 nsew signal input
rlabel metal2 s 57316 -480 57428 240 8 col_select_a[0]
port 3 nsew signal input
rlabel metal2 s 59220 -480 59332 240 8 col_select_a[1]
port 4 nsew signal input
rlabel metal2 s 61124 -480 61236 240 8 col_select_a[2]
port 5 nsew signal input
rlabel metal2 s 63028 -480 63140 240 8 col_select_a[3]
port 6 nsew signal input
rlabel metal2 s 64932 -480 65044 240 8 col_select_a[4]
port 7 nsew signal input
rlabel metal2 s 66836 -480 66948 240 8 col_select_a[5]
port 8 nsew signal input
rlabel metal2 s 5908 -480 6020 240 8 data_in_a[0]
port 9 nsew signal input
rlabel metal2 s 24948 -480 25060 240 8 data_in_a[10]
port 10 nsew signal input
rlabel metal2 s 26852 -480 26964 240 8 data_in_a[11]
port 11 nsew signal input
rlabel metal2 s 28756 -480 28868 240 8 data_in_a[12]
port 12 nsew signal input
rlabel metal2 s 30660 -480 30772 240 8 data_in_a[13]
port 13 nsew signal input
rlabel metal2 s 32564 -480 32676 240 8 data_in_a[14]
port 14 nsew signal input
rlabel metal2 s 34468 -480 34580 240 8 data_in_a[15]
port 15 nsew signal input
rlabel metal2 s 7812 -480 7924 240 8 data_in_a[1]
port 16 nsew signal input
rlabel metal2 s 9716 -480 9828 240 8 data_in_a[2]
port 17 nsew signal input
rlabel metal2 s 11620 -480 11732 240 8 data_in_a[3]
port 18 nsew signal input
rlabel metal2 s 13524 -480 13636 240 8 data_in_a[4]
port 19 nsew signal input
rlabel metal2 s 15428 -480 15540 240 8 data_in_a[5]
port 20 nsew signal input
rlabel metal2 s 17332 -480 17444 240 8 data_in_a[6]
port 21 nsew signal input
rlabel metal2 s 19236 -480 19348 240 8 data_in_a[7]
port 22 nsew signal input
rlabel metal2 s 21140 -480 21252 240 8 data_in_a[8]
port 23 nsew signal input
rlabel metal2 s 23044 -480 23156 240 8 data_in_a[9]
port 24 nsew signal input
rlabel metal2 s 2100 -480 2212 240 8 driver_io[0]
port 25 nsew signal output
rlabel metal2 s 4004 -480 4116 240 8 driver_io[1]
port 26 nsew signal output
rlabel metal2 s 87780 -480 87892 240 8 inverter_select_a
port 27 nsew signal input
rlabel metal2 s 36372 -480 36484 240 8 mem_address_a[0]
port 28 nsew signal input
rlabel metal2 s 38276 -480 38388 240 8 mem_address_a[1]
port 29 nsew signal input
rlabel metal2 s 40180 -480 40292 240 8 mem_address_a[2]
port 30 nsew signal input
rlabel metal2 s 42084 -480 42196 240 8 mem_address_a[3]
port 31 nsew signal input
rlabel metal2 s 43988 -480 44100 240 8 mem_address_a[4]
port 32 nsew signal input
rlabel metal2 s 45892 -480 46004 240 8 mem_address_a[5]
port 33 nsew signal input
rlabel metal2 s 47796 -480 47908 240 8 mem_address_a[6]
port 34 nsew signal input
rlabel metal2 s 49700 -480 49812 240 8 mem_address_a[7]
port 35 nsew signal input
rlabel metal2 s 51604 -480 51716 240 8 mem_address_a[8]
port 36 nsew signal input
rlabel metal2 s 53508 -480 53620 240 8 mem_address_a[9]
port 37 nsew signal input
rlabel metal2 s 55412 -480 55524 240 8 mem_write_n_a
port 38 nsew signal input
rlabel metal2 s 85876 -480 85988 240 8 output_active_a
port 39 nsew signal input
rlabel metal2 s 83972 -480 84084 240 8 row_col_select_a
port 40 nsew signal input
rlabel metal2 s 72548 -480 72660 240 8 row_select_a[0]
port 41 nsew signal input
rlabel metal2 s 74452 -480 74564 240 8 row_select_a[1]
port 42 nsew signal input
rlabel metal2 s 76356 -480 76468 240 8 row_select_a[2]
port 43 nsew signal input
rlabel metal2 s 78260 -480 78372 240 8 row_select_a[3]
port 44 nsew signal input
rlabel metal2 s 80164 -480 80276 240 8 row_select_a[4]
port 45 nsew signal input
rlabel metal2 s 82068 -480 82180 240 8 row_select_a[5]
port 46 nsew signal input
rlabel metal4 s 1017 1538 1327 70198 6 vccd1
port 47 nsew power bidirectional
rlabel metal4 s 19017 1538 19327 70198 6 vccd1
port 47 nsew power bidirectional
rlabel metal4 s 37017 1538 37327 70198 6 vccd1
port 47 nsew power bidirectional
rlabel metal4 s 55017 1538 55327 70198 6 vccd1
port 47 nsew power bidirectional
rlabel metal4 s 73017 1538 73327 70198 6 vccd1
port 47 nsew power bidirectional
rlabel metal4 s 2877 1538 3187 70198 6 vssd1
port 48 nsew ground bidirectional
rlabel metal4 s 20877 1538 21187 70198 6 vssd1
port 48 nsew ground bidirectional
rlabel metal4 s 38877 1538 39187 70198 6 vssd1
port 48 nsew ground bidirectional
rlabel metal4 s 56877 1538 57187 70198 6 vssd1
port 48 nsew ground bidirectional
rlabel metal4 s 74877 1538 75187 70198 6 vssd1
port 48 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 90000 72000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 17836706
string GDS_FILE /home/jasteve4/Documents/MicroMotorController/openlane/driver_core/runs/22_12_05_17_30/results/signoff/driver_core.magic.gds
string GDS_START 275842
<< end >>


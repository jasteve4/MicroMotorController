* NGSPICE file created from driver_core.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VSS
.ends

.subckt driver_core clock clock_a col_select_a[0] col_select_a[1] col_select_a[2]
+ col_select_a[3] col_select_a[4] col_select_a[5] data_in_a[0] data_in_a[10] data_in_a[11]
+ data_in_a[12] data_in_a[13] data_in_a[14] data_in_a[15] data_in_a[1] data_in_a[2]
+ data_in_a[3] data_in_a[4] data_in_a[5] data_in_a[6] data_in_a[7] data_in_a[8] data_in_a[9]
+ driver_io[0] driver_io[1] inverter_select_a mem_address_a[0] mem_address_a[1] mem_address_a[2]
+ mem_address_a[3] mem_address_a[4] mem_address_a[5] mem_address_a[6] mem_address_a[7]
+ mem_address_a[8] mem_address_a[9] mem_write_n_a output_active_a row_col_select_a
+ row_select_a[0] row_select_a[1] row_select_a[2] row_select_a[3] row_select_a[4]
+ row_select_a[5] vdd vss
XFILLER_132_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07383__I _02618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11705__I1 u2.mem\[181\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09671_ _04550_ _00582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06883_ _02338_ _02345_ _02362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__06337__A2 _01834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08582__I0 _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12595__CLK clknet_leaf_112_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08622_ _03885_ _00198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09304__S _04323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08553_ _03834_ _03845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_78_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07298__B1 _02591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07504_ u2.mem\[40\]\[7\] _02789_ _02790_ u2.mem\[30\]\[7\] _02976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_35_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08484_ _03797_ u2.mem\[9\]\[0\] _03799_ _03800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_1_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07435_ _02568_ _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10841__A1 _03982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07301__A4 _02776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10249__I _04604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07366_ _02579_ _02841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_350_clock clknet_5_4_0_clock clknet_leaf_350_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_52_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09105_ _04199_ _00367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06317_ u2.mem\[158\]\[3\] _01728_ _01729_ u2.mem\[151\]\[3\] _01731_ u2.mem\[193\]\[3\]
+ _01821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_163_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07297_ u2.mem\[23\]\[3\] _02682_ _02683_ u2.mem\[22\]\[3\] _02773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_136_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09036_ _04152_ _00345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07470__B1 _02884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06248_ u2.mem\[184\]\[1\] _01626_ _01753_ _01754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06462__I _01914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_365_clock clknet_5_4_0_clock clknet_leaf_365_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06179_ _01563_ _01677_ _01587_ _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_172_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06025__A1 _01516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07222__B1 _02634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13370__CLK clknet_leaf_375_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06576__A2 _02060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10712__I _05195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09938_ _04689_ u2.mem\[42\]\[3\] _04719_ _04723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_120_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12938__CLK clknet_leaf_148_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09869_ _04605_ u2.mem\[40\]\[12\] _04676_ _04677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06328__A2 _01712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08573__I0 _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11900_ _05927_ _05942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_133_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12880_ _00759_ clknet_5_24_0_clock u2.mem\[47\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_303_clock clknet_5_20_0_clock clknet_leaf_303_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11831_ _05870_ u2.mem\[189\]\[2\] _05896_ _05899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07289__B1 _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11762_ _04248_ _05847_ _05856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09013__I data_in_trans\[3\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13501_ _01380_ clknet_leaf_354_clock u2.mem\[187\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10713_ _05194_ u2.mem\[61\]\[0\] _05196_ _05197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12318__CLK clknet_leaf_185_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11880__I0 u2.mem\[192\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11693_ _05794_ u2.mem\[180\]\[3\] _05810_ _05814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_318_clock clknet_5_17_0_clock clknet_leaf_318_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_13_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13432_ _01311_ clknet_leaf_350_clock u2.mem\[175\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08852__I _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10644_ _05156_ _00949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11632__I0 _05756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13363_ _01242_ clknet_leaf_374_clock u2.mem\[164\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10575_ _05114_ _00922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07056__A3 _02503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12314_ _00193_ clknet_leaf_116_clock u2.mem\[11\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13294_ _01173_ clknet_leaf_383_clock u2.mem\[152\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11919__S _05950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12245_ _00124_ clknet_leaf_74_clock u2.mem\[7\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08005__A2 _03464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07213__B1 _02690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11935__I1 u2.mem\[193\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12176_ _00055_ clknet_leaf_233_clock u2.mem\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11718__I _03661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08299__I _03674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11127_ _05457_ _01131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_142_clock_I clknet_5_13_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11058_ _05384_ u2.mem\[141\]\[1\] _05413_ _05415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07516__A1 u2.mem\[58\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10009_ _04685_ u2.mem\[44\]\[1\] _04762_ _04764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_64_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08316__I0 _03688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10069__I _04591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11871__I0 _05915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13243__CLK clknet_leaf_289_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07220_ _02674_ _02681_ _02688_ _02697_ _02698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_20_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07151_ u2.mem\[5\]\[0\] _02627_ _02629_ u2.mem\[38\]\[0\] _02630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_leaf_67_clock_I clknet_5_9_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09292__I1 u2.mem\[27\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07378__I _02605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06102_ _01547_ _01608_ _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_121_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09794__S _04633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07082_ _02448_ _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06255__B2 u2.mem\[188\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13393__CLK clknet_leaf_327_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11829__S _05896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06033_ _01528_ _01540_ _01541_ _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_173_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11926__I1 u2.mem\[193\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08203__S _03608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07984_ u2.mem\[17\]\[15\] _03312_ _03313_ u2.mem\[24\]\[15\] _03448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_101_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09723_ data_in_trans\[6\].data_sync _04585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06935_ _01551_ _02016_ _02414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11564__S _05731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09654_ _04496_ u2.mem\[35\]\[14\] _04537_ _04540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06866_ _02339_ _02344_ _02345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07841__I _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08605_ _03874_ _00192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09585_ _04500_ _04501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06797_ u2.mem\[164\]\[4\] _02050_ _02053_ u2.mem\[178\]\[4\] _02278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_58_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06730__A2 _02043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09969__S _04740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08536_ _03797_ u2.mem\[10\]\[0\] _03835_ _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_344_clock_I clknet_5_7_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08467_ _03789_ _00139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10908__S _05319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07286__A3 _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07418_ _02520_ _02892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08672__I _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08398_ _03746_ _00113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07349_ _02793_ _02805_ _02814_ _02823_ _02824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__11614__I0 _05754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08235__A2 mem_address_trans\[3\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06246__A1 u2.mem\[171\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07443__B1 _02916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10360_ _04978_ _00843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06246__B2 u2.mem\[157\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06192__I _01698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07994__A1 _01980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06797__A2 _02050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11739__S _05840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09019_ _04138_ _04139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10291_ _04913_ u2.mem\[50\]\[12\] _04938_ _04939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10643__S _05152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12760__CLK clknet_leaf_52_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12030_ row_select_trans\[2\].A clknet_leaf_303_clock row_select_trans\[2\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11917__I1 u2.mem\[193\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06549__A2 _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09008__I data_in_trans\[2\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13116__CLK clknet_leaf_276_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12932_ _00811_ clknet_leaf_64_clock u2.mem\[50\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_242_clock clknet_5_25_0_clock clknet_leaf_242_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12863_ _00742_ clknet_leaf_154_clock u2.mem\[46\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12140__CLK clknet_leaf_225_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06721__A2 _01995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11814_ _05889_ _01386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12794_ _00673_ clknet_leaf_338_clock u2.mem\[41\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11745_ _05837_ u2.mem\[183\]\[5\] _05839_ _05846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_257_clock clknet_5_19_0_clock clknet_leaf_257_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_144_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09678__I _04543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07682__B1 _03083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12290__CLK clknet_leaf_179_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11676_ _05792_ u2.mem\[179\]\[2\] _05801_ _05804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13415_ _01294_ clknet_leaf_357_clock u2.mem\[172\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10617__I _05130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10627_ _05121_ u2.mem\[58\]\[12\] _05146_ _05147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07198__I _02568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09274__I1 u2.mem\[26\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13346_ _01225_ clknet_leaf_3_clock u2.mem\[161\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10558_ _05102_ _00917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06788__A2 _02267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13277_ _01156_ clknet_leaf_8_clock u2.mem\[149\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10489_ _05050_ _05061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_12228_ _00107_ clknet_leaf_73_clock u2.mem\[6\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07737__A1 _03190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07147__B _02474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12159_ _00038_ clknet_leaf_236_clock u2.mem\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08958__S _04097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_293_clock_I clknet_5_21_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06720_ _02179_ _02190_ _02194_ _02203_ _02204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_110_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06651_ _02119_ _02044_ _02136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_37_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09789__S _04628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09370_ _04363_ _00468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08693__S _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06582_ _02045_ _02018_ _02067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_17_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12633__CLK clknet_leaf_115_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08321_ _03658_ _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_36_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08252_ _03559_ u2.mem\[4\]\[6\] _03639_ _03642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07673__B1 _03142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08492__I _03670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07203_ _02677_ _02678_ _02679_ _02680_ _02681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_119_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08183_ _03599_ _00045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10527__I _05072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07134_ u2.mem\[8\]\[0\] _02610_ _02612_ u2.mem\[4\]\[0\] _02613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_14_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11221__A1 _05354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06779__A2 _02042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07065_ _02543_ _02544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12013__CLK clknet_2_3__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06016_ u2.driver_mem\[5\] _01517_ _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__13139__CLK clknet_leaf_34_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08776__I0 _03938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11524__A2 _05690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10583__I0 _05119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input36_I row_col_select_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06400__A1 u2.mem\[144\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06400__B2 u2.mem\[182\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07967_ u2.mem\[44\]\[15\] _02514_ _02518_ u2.mem\[42\]\[15\] _03431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_114_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12163__CLK clknet_leaf_79_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11294__S _05558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13289__CLK clknet_leaf_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09706_ _04130_ _04572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06918_ _02396_ _02397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07898_ u2.mem\[17\]\[13\] _03312_ _03313_ u2.mem\[24\]\[13\] _03364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07571__I _02482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09637_ _04530_ _00568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06849_ u2.mem\[154\]\[5\] _02225_ _02226_ u2.mem\[162\]\[5\] _02328_ _02329_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_15_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07900__B2 u2.mem\[19\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06187__I _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09568_ _04163_ _04489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08519_ _03823_ u2.mem\[9\]\[11\] _03817_ _03824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_93_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11835__I0 _05874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09499_ _04445_ _00515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11530_ _05712_ _01279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07664__B1 _03133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06915__I _02362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11461_ _05667_ _05668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13200_ _01079_ clknet_leaf_291_clock u2.mem\[136\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06219__A1 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10412_ _05014_ u2.mem\[53\]\[9\] _05012_ _05015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11392_ _05295_ _05606_ _05624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_104_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13131_ _01010_ clknet_leaf_261_clock u2.mem\[63\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10343_ _04891_ u2.mem\[52\]\[2\] _04966_ _04969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_124_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10274_ _04929_ _00806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13062_ _00941_ clknet_leaf_30_clock u2.mem\[58\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07982__A4 _03445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08767__I0 _03929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12013_ net28 clknet_2_3__leaf_clock_a mem_address_trans\[4\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10574__I0 _05112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07195__A2 _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_181_clock clknet_5_27_0_clock clknet_leaf_181_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_15_clock_I clknet_5_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08519__I0 _03823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12656__CLK clknet_leaf_235_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12915_ _00794_ clknet_leaf_87_clock u2.mem\[49\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06155__C2 u2.mem\[181\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06097__I _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_196_clock clknet_5_31_0_clock clknet_leaf_196_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_146_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12846_ _00725_ clknet_leaf_214_clock u2.mem\[45\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09402__S _04385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10629__I1 u2.mem\[58\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12777_ _00656_ clknet_leaf_147_clock u2.mem\[40\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10548__S _05095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11728_ _05835_ u2.mem\[182\]\[4\] _05826_ _05836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_159_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09201__I _04135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10347__I _04965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11659_ _05792_ u2.mem\[178\]\[2\] _05788_ _05793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06046__B _01552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12036__CLK clknet_leaf_303_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13329_ _01208_ clknet_leaf_1_clock u2.mem\[158\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_134_clock clknet_5_15_0_clock clknet_leaf_134_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_118_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08758__I0 _03920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12186__CLK clknet_leaf_59_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10082__I _04604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08870_ _04044_ u2.mem\[17\]\[13\] _04042_ _04045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_123_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07186__A2 _02661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07821_ u2.mem\[43\]\[12\] _03286_ _03287_ u2.mem\[20\]\[12\] _03288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_149_clock clknet_5_13_0_clock clknet_leaf_149_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_85_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10810__I _05252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07752_ u2.mem\[53\]\[11\] _03041_ _03042_ u2.mem\[56\]\[11\] _03220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06703_ _02101_ _02187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07683_ u2.mem\[18\]\[9\] _03085_ _03086_ u2.mem\[19\]\[9\] _03153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07489__A3 _02960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08930__I0 _04026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09422_ _04399_ _00484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06697__A1 u2.mem\[167\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06697__B2 u2.mem\[183\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06634_ _02027_ _02017_ _02119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09353_ _04352_ _00462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11817__I0 _05870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06565_ _02031_ _02041_ _02050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_90_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06449__A1 _01878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08304_ _03678_ _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06449__B2 _01944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09284_ _04311_ _04250_ _04312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06496_ _01981_ _01927_ _01982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_166_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09111__I _04202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08235_ _03630_ mem_address_trans\[3\].data_sync _03631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09238__I1 u2.mem\[25\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07661__A3 _03121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08166_ _03584_ _03590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_101_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07117_ _02595_ _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12529__CLK clknet_leaf_178_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08097_ _03540_ _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_49_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08610__A2 _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09982__S _04745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07048_ _02418_ _02433_ _02434_ _02454_ _02527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__06621__A1 u2.mem\[188\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06621__B2 u2.mem\[175\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08749__I0 _03911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07177__A2 _02652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07716__A4 _03184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08999_ _04121_ _04122_ _04123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_189_clock_I clknet_5_30_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10961_ _05354_ _05317_ _05355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_112_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11752__S _05849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08921__I0 _04017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12700_ _00579_ clknet_leaf_222_clock u2.mem\[36\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06688__A1 u2.mem\[151\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06688__B2 u2.mem\[158\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10892_ _05309_ _05310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09222__S _04270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12631_ _00510_ clknet_leaf_113_clock u2.mem\[31\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11808__I0 _05876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_241_clock_I clknet_5_25_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12059__CLK clknet_2_1__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12562_ _00441_ clknet_leaf_160_clock u2.mem\[27\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09021__I _04123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11513_ _05668_ u2.mem\[169\]\[1\] _05700_ _05702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12493_ _00372_ clknet_leaf_197_clock u2.mem\[23\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_51_clock clknet_5_13_0_clock clknet_leaf_51_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11444_ _05627_ u2.mem\[165\]\[1\] _05655_ _05657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_172_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11199__S _05502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13454__CLK clknet_leaf_320_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11375_ _05595_ u2.mem\[160\]\[5\] _05607_ _05614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13114_ _00993_ clknet_leaf_45_clock u2.mem\[61\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10326_ _04958_ _00829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_66_clock clknet_5_9_0_clock clknet_leaf_66_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13045_ _00924_ clknet_leaf_28_clock u2.mem\[57\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10257_ _04918_ u2.mem\[49\]\[14\] _04914_ _04919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10831__S _05268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10188_ _04873_ _00776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10172__A1 _03982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11662__S _05788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06679__A1 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07876__B1 _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09132__S _04213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07340__A2 _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12829_ _00708_ clknet_leaf_203_clock u2.mem\[44\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11461__I _05667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06350_ _01849_ _01850_ _01851_ _01852_ _01853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_163_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07628__B1 _03057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06281_ u2.mem\[175\]\[2\] _01602_ _01632_ u2.mem\[188\]\[2\] _01786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_72_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_19_clock clknet_5_2_0_clock clknet_leaf_19_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_129_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08020_ mem_address_trans\[0\].data_sync _03481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_141_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07386__I _02611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06603__A1 _01992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09971_ _04685_ u2.mem\[43\]\[1\] _04740_ _04742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11837__S _05895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08922_ _04076_ _00307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07159__A2 _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08853_ _04014_ _04033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_131_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06367__B1 _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_190_clock_I clknet_5_30_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07804_ _03262_ _03265_ _03268_ _03270_ _03271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_61_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12971__CLK clknet_leaf_266_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08784_ _03987_ _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05996_ u2.select_mem_col\[0\] _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_73_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07735_ u2.mem\[6\]\[10\] _03160_ _03161_ u2.mem\[47\]\[10\] _03204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08945__I _04073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07666_ u2.mem\[37\]\[9\] _03062_ _03063_ u2.mem\[59\]\[9\] _03136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_168_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12201__CLK clknet_leaf_42_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07331__A2 _02647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13327__CLK clknet_leaf_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06134__A3 _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09405_ _04387_ u2.mem\[29\]\[13\] _04385_ _04388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06617_ u2.mem\[187\]\[0\] _02100_ _02101_ u2.mem\[192\]\[0\] _02102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_90_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07597_ _02558_ _03068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09336_ _04263_ u2.mem\[28\]\[5\] _04341_ _04343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06548_ _02032_ _02010_ _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09267_ _04272_ u2.mem\[26\]\[9\] _04300_ _04302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10916__S _05318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06479_ _01966_ _01955_ _01967_ _01968_ _01460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08218_ _03620_ _00059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06842__A1 u2.mem\[145\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06842__B2 u2.mem\[168\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09198_ _04131_ _04256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08149_ _03578_ _00032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11160_ _05468_ u2.mem\[147\]\[3\] _05475_ _05479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10111_ _04828_ _00744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11091_ _05436_ _01116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06070__A2 _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09395__I0 _04380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10042_ _04564_ _04782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06373__A3 _01862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11993_ _00005_ clknet_leaf_334_clock u2.mem\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11482__S _05683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10944_ _04130_ _05342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10875_ _05298_ _01038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12614_ _00493_ clknet_leaf_92_clock u2.mem\[30\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08791__S _03990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12545_ _00424_ clknet_leaf_178_clock u2.mem\[26\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10826__S _05263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06833__A1 u2.mem\[180\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08590__I _03855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12476_ _00355_ clknet_leaf_195_clock u2.mem\[22\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06833__B2 u2.mem\[172\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12844__CLK clknet_leaf_215_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11427_ _05646_ _05647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07389__A2 _02859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11358_ _05603_ _01216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10309_ _04943_ _04949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10561__S _05104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11289_ _05561_ _01189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09127__S _04208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13028_ _00907_ clknet_leaf_67_clock u2.mem\[56\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11193__I0 _05472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07010__A1 _02455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12224__CLK clknet_leaf_241_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07561__A2 _03030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07520_ u2.mem\[49\]\[7\] _02817_ _02818_ u2.mem\[46\]\[7\] _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_169_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07451_ u2.mem\[39\]\[5\] _02857_ _02858_ u2.mem\[48\]\[5\] _02925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_90_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07864__A3 _03321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06402_ u2.mem\[170\]\[5\] _01686_ _01688_ u2.mem\[156\]\[5\] _01904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11248__I1 u2.mem\[152\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07382_ _02616_ _02857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09310__I0 _04276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09121_ _04140_ u2.mem\[23\]\[4\] _04208_ _04209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07077__A1 u2.mem\[61\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06333_ u2.mem\[191\]\[3\] _01682_ _01684_ u2.mem\[179\]\[3\] _01837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_leaf_137_clock_I clknet_5_14_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06285__C1 u2.mem\[165\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09052_ _04164_ u2.mem\[21\]\[11\] _04155_ _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06264_ _01763_ _01764_ _01769_ _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06824__A1 _01844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08003_ u2.active_mem\[8\] _03458_ _03459_ u2.active_mem\[9\] _03466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06195_ _01561_ _01563_ _01580_ _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_85_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09954_ _04705_ u2.mem\[42\]\[10\] _04729_ _04732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08905_ _04065_ _00301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09885_ _04572_ _04687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08836_ _03670_ _04021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08767_ _03929_ u2.mem\[15\]\[11\] _03972_ _03976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06760__B1 _02177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11636__A1 _05285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07718_ u2.mem\[60\]\[10\] _03059_ _03060_ u2.mem\[62\]\[10\] _03187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08675__I _03687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08698_ _03717_ _03936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07304__A2 _02610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07649_ u2.mem\[53\]\[9\] _03041_ _03042_ u2.mem\[56\]\[9\] _03119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_15_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06409__B _01910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10660_ _05165_ _00956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09301__I0 _04267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09500__S _04443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09319_ _04285_ u2.mem\[27\]\[15\] _04328_ _04332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07068__A1 _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10591_ _05125_ _00927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12330_ _00209_ clknet_leaf_136_clock u2.mem\[12\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06815__A1 u2.mem\[194\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12261_ _00140_ clknet_leaf_23_clock u2.mem\[8\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11212_ _05512_ _01161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12192_ _00071_ clknet_leaf_253_clock u2.mem\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_162_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11143_ _05345_ _05468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_339_clock_I clknet_5_7_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07240__B2 u2.mem\[20\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12247__CLK clknet_leaf_56_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07791__A2 _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11074_ _05424_ u2.mem\[142\]\[1\] _05422_ _05425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11175__I0 _05468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10025_ _04700_ u2.mem\[44\]\[8\] _04772_ _04773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10922__I0 _05294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12397__CLK clknet_leaf_193_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06751__B1 _02152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11478__I1 u2.mem\[166\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11976_ _05218_ u2.mem\[194\]\[10\] _05985_ _05986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_17_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09540__I0 _04469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10927_ _05330_ _01058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10858_ _05194_ u2.mem\[129\]\[0\] _05287_ _05288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07059__A1 _02463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13577_ _01456_ clknet_leaf_35_clock u2.mem\[194\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10789_ _05220_ u2.mem\[62\]\[11\] _05242_ _05246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06806__A1 u2.mem\[180\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12528_ _00407_ clknet_leaf_189_clock u2.mem\[25\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06806__B2 u2.mem\[172\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12459_ _00338_ clknet_leaf_188_clock u2.mem\[21\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13022__CLK clknet_leaf_272_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11387__S _05615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07231__A1 _02704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10291__S _04938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06034__A2 _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07782__A2 _03017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13172__CLK clknet_leaf_278_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06951_ _02428_ _02405_ _02429_ _02430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_80_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09670_ _04473_ u2.mem\[36\]\[4\] _04549_ _04550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08696__S _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06882_ _02360_ _02361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07534__A2 _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_63_clock_I clknet_5_9_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08621_ _03807_ u2.mem\[12\]\[4\] _03884_ _03885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11914__I _05949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08552_ _03844_ _00169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08495__I _03674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07503_ u2.mem\[32\]\[7\] _02786_ _02787_ u2.mem\[2\]\[7\] _02975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_78_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07298__A1 u2.mem\[17\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08483_ _03798_ _03799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_35_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07434_ _02566_ _02908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07365_ u2.mem\[9\]\[4\] _02838_ _02839_ u2.mem\[25\]\[4\] _02840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_4_15_0_clock clknet_3_7_0_clock clknet_4_15_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_149_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10466__S _05045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_288_clock_I clknet_5_20_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09104_ _04171_ u2.mem\[22\]\[13\] _04197_ _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06316_ u2.mem\[177\]\[3\] _01734_ _01646_ u2.mem\[165\]\[3\] u2.mem\[163\]\[3\]
+ _01643_ _01820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_149_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06743__I _02127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07296_ _02768_ _02769_ _02770_ _02771_ _02772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_11_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09035_ _04151_ u2.mem\[21\]\[7\] _04141_ _04152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06247_ _01553_ _01753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06178_ u2.mem\[191\]\[0\] _01682_ _01684_ u2.mem\[179\]\[0\] _01685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__13515__CLK clknet_leaf_347_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_340_clock_I clknet_5_7_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08270__I0 _03577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07574__I _02489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07773__A2 _03082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09937_ _04722_ _00676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09868_ _04660_ _04676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08819_ _04008_ _00272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09799_ _04636_ _00624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06733__B1 _02177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11830_ _05898_ _01393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06918__I _02396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11761_ _05855_ _01367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11760__S _05848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13500_ _01379_ clknet_leaf_331_clock u2.mem\[186\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10712_ _05195_ _05196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11692_ _05813_ _01340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11880__I1 _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13431_ _01310_ clknet_leaf_350_clock u2.mem\[175\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10643_ _05101_ u2.mem\[59\]\[3\] _05152_ _05156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13362_ _01241_ clknet_leaf_368_clock u2.mem\[163\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11632__I1 u2.mem\[176\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10574_ _05112_ u2.mem\[57\]\[8\] _05113_ _05114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07056__A4 _02534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12313_ _00192_ clknet_leaf_116_clock u2.mem\[11\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07461__A1 u2.mem\[40\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07461__B2 u2.mem\[30\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13293_ _01172_ clknet_leaf_384_clock u2.mem\[152\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12244_ _00123_ clknet_leaf_73_clock u2.mem\[7\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13195__CLK clknet_leaf_294_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06016__A2 _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08261__I0 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12175_ _00054_ clknet_leaf_236_clock u2.mem\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07213__B2 u2.mem\[38\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11000__S _05372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07764__A2 _03137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11126_ _05428_ u2.mem\[145\]\[3\] _05453_ _05457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_150_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11057_ _05414_ _01104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09405__S _04385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10008_ _04763_ _00706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06724__B1 _02068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09204__I _04139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08316__I1 u2.mem\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11959_ _05976_ _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11871__I1 u2.mem\[191\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10286__S _04933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07150_ _02628_ _02629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12412__CLK clknet_leaf_192_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13538__CLK clknet_leaf_34_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06101_ _01584_ _01559_ _01608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07081_ _02446_ _02560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_173_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06032_ u2.select_mem_row\[3\] u2.select_mem_col\[3\] _01515_ _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08252__I0 _03559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07755__A2 _03122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07983_ u2.mem\[23\]\[15\] _02594_ _02596_ u2.mem\[22\]\[15\] _03447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09722_ _04584_ _00599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06934_ _02388_ _02413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09653_ _04539_ _00575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06865_ _02340_ _02341_ _02342_ _02343_ _02344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08604_ _03830_ u2.mem\[11\]\[14\] _03871_ _03874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09584_ _03583_ _04441_ _04500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06191__A1 _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06796_ _02273_ _02274_ _02275_ _02276_ _02277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_58_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08535_ _03834_ _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_82_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11311__I0 _05556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11580__S _05739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08466_ _03697_ u2.mem\[8\]\[9\] _03787_ _03789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07286__A4 _02761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07417_ u2.mem\[44\]\[5\] _02889_ _02890_ u2.mem\[42\]\[5\] _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08397_ _03722_ u2.mem\[6\]\[15\] _03742_ _03746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12092__CLK clknet_leaf_304_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06473__I _01913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07348_ _02815_ _02816_ _02819_ _02822_ _02823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_13_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07038__A4 _02485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06246__A2 _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07443__A1 u2.mem\[23\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07443__B2 u2.mem\[22\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07279_ u2.mem\[58\]\[3\] _02487_ _02490_ u2.mem\[36\]\[3\] _02755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10924__S _05327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12905__CLK clknet_leaf_52_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09784__I _04617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09018_ data_in_trans\[4\].data_sync _04138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10290_ _04922_ _04938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08243__I0 _03550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07746__A2 _03033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09991__I0 _04705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07210__A4 _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09225__S _04270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12931_ _00810_ clknet_leaf_65_clock u2.mem\[50\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12862_ _00741_ clknet_leaf_204_clock u2.mem\[46\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09024__I data_in_trans\[5\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11813_ _05864_ u2.mem\[188\]\[0\] _05888_ _05889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12793_ _00672_ clknet_leaf_340_clock u2.mem\[41\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11490__S _05682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11744_ _05845_ _01360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12435__CLK clknet_leaf_102_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11675_ _05803_ _01333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_169_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13414_ _01293_ clknet_leaf_357_clock u2.mem\[172\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_11_clock_I clknet_5_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10626_ _05130_ _05146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_122_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06237__A2 _01741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13345_ _01224_ clknet_leaf_3_clock u2.mem\[161\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12585__CLK clknet_leaf_117_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10557_ _05101_ u2.mem\[57\]\[3\] _05095_ _05102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13276_ _01155_ clknet_leaf_8_clock u2.mem\[149\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10488_ _05060_ _00889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11369__I0 _05589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12227_ _00106_ clknet_leaf_68_clock u2.mem\[6\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07737__A2 _03195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09982__I0 _04696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12158_ _00037_ clknet_leaf_219_clock u2.mem\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07147__C _02562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_236_clock_I clknet_5_25_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11665__S _05787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11109_ _05447_ _01123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12089_ net35 clknet_2_2__leaf_clock_a output_active_trans.A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09734__I0 _04592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11464__I _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11541__I0 _05719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06558__I _02042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06650_ u2.mem\[194\]\[0\] _02133_ _02134_ u2.mem\[190\]\[0\] _02135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07370__B1 _02683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06581_ _02065_ _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_364_clock clknet_5_4_0_clock clknet_leaf_364_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08320_ _03691_ _03692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13360__CLK clknet_leaf_371_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08251_ _03641_ _00071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07673__A1 u2.mem\[26\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12928__CLK clknet_leaf_243_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07202_ u2.mem\[28\]\[1\] _02580_ _02582_ u2.mem\[31\]\[1\] _02680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_144_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08182_ _03570_ u2.mem\[2\]\[11\] _03595_ _03599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_379_clock clknet_5_0_0_clock clknet_leaf_379_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_105_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07133_ _02611_ _02612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08473__I0 _03709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07976__A2 _02548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07064_ _02408_ _02515_ _02516_ _02406_ _02543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xclkbuf_leaf_302_clock clknet_5_21_0_clock clknet_leaf_302_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06015_ u2.driver_mem\[6\] _01522_ _01523_ _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_47_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07728__A2 _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09973__I0 _04687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06400__A2 _01670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07966_ _03426_ _03427_ _03428_ _03429_ _03430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xclkbuf_leaf_317_clock clknet_5_16_0_clock clknet_leaf_317_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07852__I _02605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09705_ _04571_ _00595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09725__I0 _04586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06917_ _02387_ _02389_ _02393_ _02395_ _02396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_114_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06951__A3 _02429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input29_I mem_address_a[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07897_ u2.mem\[23\]\[13\] _02594_ _02596_ u2.mem\[22\]\[13\] _03363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11532__I0 _05713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09636_ _04478_ u2.mem\[35\]\[6\] _04527_ _04530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06848_ _02325_ _02326_ _02327_ _02328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_55_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06468__I _01927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08884__S _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12458__CLK clknet_leaf_135_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09567_ _04488_ _00540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06779_ u2.mem\[180\]\[3\] _02042_ _02012_ u2.mem\[172\]\[3\] _02261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10099__I0 _04786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08518_ _03704_ _03823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07113__B1 _02591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09498_ _04360_ u2.mem\[32\]\[1\] _04443_ _04445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11835__I1 u2.mem\[189\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08449_ _03779_ _00131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06467__A2 _01929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07664__A1 u2.mem\[61\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11460_ _03495_ _05667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_185_clock_I clknet_5_30_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10411_ _03695_ _05014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08464__I0 _03692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11391_ _05499_ _05623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07967__A2 _02514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13130_ _01009_ clknet_5_6_0_clock u2.mem\[62\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10342_ _04968_ _00835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06931__I _02409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13061_ _00940_ clknet_leaf_29_clock u2.mem\[58\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10273_ _04895_ u2.mem\[50\]\[4\] _04928_ _04929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09019__I _04138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12012_ mem_address_trans\[3\].A clknet_leaf_315_clock mem_address_trans\[3\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07719__A2 _03062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13233__CLK clknet_leaf_303_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12914_ _00793_ clknet_leaf_163_clock u2.mem\[49\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06155__B2 u2.mem\[155\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13383__CLK clknet_leaf_318_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12845_ _00724_ clknet_leaf_214_clock u2.mem\[45\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10829__S _05268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12776_ _00655_ clknet_leaf_58_clock u2.mem\[40\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07104__B1 _02582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11727_ _03673_ _05835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06458__A2 _01946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11658_ _05670_ _05792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07670__A4 _03139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10609_ _05103_ u2.mem\[58\]\[4\] _05136_ _05137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08455__I0 _03675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10564__S _05104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11589_ _05746_ u2.mem\[174\]\[0\] _05748_ _05749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13328_ _01207_ clknet_leaf_1_clock u2.mem\[158\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08080__A1 _03527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13259_ _01138_ clknet_leaf_311_clock u2.mem\[146\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07820_ _02507_ _03287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07672__I _02568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12600__CLK clknet_leaf_115_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07751_ u2.mem\[54\]\[11\] _03116_ _03117_ u2.mem\[55\]\[11\] _03219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_78_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06702_ _02100_ _02186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07682_ u2.mem\[52\]\[9\] _03082_ _03083_ u2.mem\[21\]\[9\] _03152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06146__A1 _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09421_ _04362_ u2.mem\[30\]\[2\] _04396_ _04399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06633_ u2.mem\[144\]\[0\] _02115_ _02117_ u2.mem\[182\]\[0\] _02118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_64_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06697__A2 _02058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07894__B2 u2.mem\[25\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12750__CLK clknet_leaf_271_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09352_ _04278_ u2.mem\[28\]\[12\] _04351_ _04352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06564_ _02021_ _02040_ _02048_ _02049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11817__I1 u2.mem\[188\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08303_ _03509_ _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06449__A2 _01938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09283_ _04310_ _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06495_ u2.mem\[192\]\[15\] _01981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_166_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08234_ mem_address_trans\[2\].data_sync _03630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_165_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13106__CLK clknet_leaf_330_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07661__A4 _03130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08165_ _03589_ _00037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08446__I0 _03656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10474__S _05051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_241_clock clknet_5_25_0_clock clknet_leaf_241_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_147_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07116_ _02587_ _02588_ _02497_ _02589_ _02595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_107_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08096_ _03478_ _03539_ _03540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_69_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08610__A3 _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12130__CLK clknet_leaf_35_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07047_ u2.mem\[14\]\[0\] _02521_ _02525_ u2.mem\[12\]\[0\] _02526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__13256__CLK clknet_leaf_287_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_256_clock clknet_5_19_0_clock clknet_leaf_256_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_173_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08678__I _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08998_ _03987_ _04122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06385__A1 _01883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07582__I _02504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07949_ _03410_ _03411_ _03412_ _03413_ _03414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_29_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11505__I0 _05677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06198__I _01704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10960_ _03750_ _05354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_60_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07885__A1 _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09619_ _04498_ u2.mem\[34\]\[15\] _04516_ _04520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10891_ _04072_ _05276_ _05309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_71_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12630_ _00509_ clknet_leaf_95_clock u2.mem\[31\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06926__I _02404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11808__I1 u2.mem\[187\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11998__CLK clknet_5_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12561_ _00440_ clknet_leaf_161_clock u2.mem\[27\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10492__I0 _05014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11512_ _05701_ _01272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12492_ _00371_ clknet_leaf_197_clock u2.mem\[23\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08437__I0 _03718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11443_ _05656_ _01248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06860__A2 _01989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_209_clock clknet_5_28_0_clock clknet_leaf_209_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11197__A1 _04179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10244__I0 _04909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06661__I _02145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08062__A1 _01951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11374_ _05613_ _01222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13113_ _00992_ clknet_leaf_39_clock u2.mem\[61\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10325_ _04911_ u2.mem\[51\]\[11\] _04954_ _04958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08789__S _03990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13044_ _00923_ clknet_leaf_33_clock u2.mem\[57\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10256_ _04611_ _04918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10187_ _04797_ u2.mem\[48\]\[6\] _04870_ _04873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_66_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10172__A2 _04863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12773__CLK clknet_leaf_76_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12828_ _00707_ clknet_leaf_203_clock u2.mem\[44\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12003__CLK clknet_leaf_41_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07891__A4 _03356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07628__A1 _01954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08676__I0 _03920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12759_ _00638_ clknet_leaf_53_clock u2.mem\[39\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10483__I0 _05005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06280_ u2.mem\[187\]\[2\] _01634_ _01637_ u2.mem\[192\]\[2\] _01785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_147_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06300__A1 u2.mem\[147\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06300__B2 u2.mem\[169\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12153__CLK clknet_leaf_56_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08428__I0 _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13279__CLK clknet_leaf_380_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06851__A2 _02145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07667__I _02547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06571__I _02005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09970_ _04741_ _00690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06603__A2 _02080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08699__S _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08921_ _04017_ u2.mem\[19\]\[1\] _04074_ _04076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09928__I0 _04716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11735__I0 _05825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08852_ _03691_ _04032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08600__I0 _03825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_133_clock_I clknet_5_15_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07564__B1 _03034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06367__B2 u2.mem\[156\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07803_ u2.mem\[3\]\[12\] _03269_ _03215_ _03270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_61_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08783_ _03983_ _03984_ _03985_ _03986_ _03987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_05995_ _01503_ _01504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07734_ u2.mem\[8\]\[10\] _03093_ _03094_ u2.mem\[4\]\[10\] _03203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_72_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06119__A1 _01586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07867__A1 u2.mem\[32\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07665_ u2.mem\[60\]\[9\] _03059_ _03060_ u2.mem\[62\]\[9\] _03135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11652__I _05787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09404_ _04170_ _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06616_ _01992_ _02001_ _02101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_77_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07596_ u2.mem\[26\]\[8\] _02908_ _02909_ u2.mem\[10\]\[8\] _03067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_40_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09335_ _04342_ _00454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08667__I0 _03913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06547_ _01985_ _02025_ _02032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10474__I0 _04992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09266_ _04301_ _00426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06478_ u2.mem\[193\]\[11\] _01960_ _01948_ u2.mem\[192\]\[11\] _01964_ _01968_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_21_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_180_clock clknet_5_27_0_clock clknet_leaf_180_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08217_ _03566_ u2.mem\[3\]\[9\] _03618_ _03620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08419__I0 _03684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09197_ _04255_ _00403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_58_clock_I clknet_5_12_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09993__S _04750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08148_ _03577_ u2.mem\[1\]\[14\] _03573_ _03578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06481__I _01920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12646__CLK clknet_leaf_94_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10932__S _05326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08079_ _03492_ _03528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_195_clock clknet_5_31_0_clock clknet_leaf_195_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_161_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10110_ _04797_ u2.mem\[46\]\[6\] _04825_ _04828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09919__I0 _04709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11090_ _05420_ u2.mem\[143\]\[0\] _05435_ _05436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10041_ _04781_ _00721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10731__I _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06358__A1 u2.mem\[166\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06358__B2 u2.mem\[161\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06373__A4 _01875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12026__CLK clknet_leaf_304_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11992_ _00004_ clknet_leaf_331_clock u2.mem\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10943_ _05341_ _01063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07858__B2 u2.mem\[48\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_133_clock clknet_5_15_0_clock clknet_leaf_133_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_147_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10874_ _05294_ u2.mem\[130\]\[0\] _05297_ _05298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_335_clock_I clknet_5_18_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12613_ _00492_ clknet_leaf_92_clock u2.mem\[30\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12544_ _00423_ clknet_leaf_188_clock u2.mem\[26\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07086__A2 _02559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_148_clock clknet_5_13_0_clock clknet_leaf_148_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12475_ _00354_ clknet_leaf_177_clock u2.mem\[22\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06833__A2 _02042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11426_ _04094_ _05645_ _05646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07389__A3 _02862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11357_ _05593_ u2.mem\[159\]\[4\] _05597_ _05603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09408__S _04385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10308_ _04948_ _00821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11288_ _05548_ u2.mem\[155\]\[1\] _05559_ _05561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_45_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13027_ _00906_ clknet_leaf_30_clock u2.mem\[56\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10239_ _04906_ _00794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06349__A1 u2.mem\[184\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11193__I1 u2.mem\[149\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08111__I _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09143__S _04218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12519__CLK clknet_leaf_125_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11472__I _03505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07450_ u2.mem\[5\]\[5\] _02922_ _02923_ u2.mem\[38\]\[5\] _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08982__S _04107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06566__I _02050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07864__A4 _03330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06401_ u2.mem\[173\]\[5\] _01719_ _01721_ u2.mem\[185\]\[5\] _01903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07381_ u2.mem\[5\]\[4\] _02689_ _02690_ u2.mem\[38\]\[4\] _02856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09120_ _04202_ _04208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_52_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09310__I1 u2.mem\[27\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06332_ u2.mem\[170\]\[3\] _01687_ _01689_ u2.mem\[156\]\[3\] _01836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08781__I mem_address_trans\[6\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07077__A2 _02553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12669__CLK clknet_leaf_217_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09051_ _04163_ _04164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06285__B1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06285__C2 _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06263_ _01765_ _01766_ _01767_ _01768_ _01769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_117_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07397__I _02419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08002_ u2.active_mem\[11\] _03461_ _03462_ u2.active_mem\[10\] _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_102_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08026__A1 _03479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06194_ _01700_ _01701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06007__S _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10752__S _05223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06588__A1 u2.mem\[184\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09953_ _04731_ _00683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08904_ _04039_ u2.mem\[18\]\[11\] _04061_ _04065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_170_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12049__CLK clknet_2_1__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09884_ _04686_ _00659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_284_clock_I clknet_5_20_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_11_0_clock clknet_3_5_0_clock clknet_4_11_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_4119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08835_ _04020_ _00276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08766_ _03975_ _00252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07860__I _02611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_50_clock clknet_5_7_0_clock clknet_leaf_50_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_input11_I data_in_a[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06760__A1 u2.mem\[188\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07717_ u2.mem\[61\]\[10\] _03132_ _03133_ u2.mem\[63\]\[10\] _03186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12199__CLK clknet_leaf_42_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08697_ _03935_ _00223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13444__CLK clknet_leaf_364_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10695__I0 _05115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07648_ u2.mem\[54\]\[9\] _03116_ _03117_ u2.mem\[55\]\[9\] _03118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_41_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07579_ _02527_ _03050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_65_clock clknet_5_9_0_clock clknet_leaf_65_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_107_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09318_ _04331_ _00448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09301__I1 u2.mem\[27\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08691__I _03708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10590_ _05124_ u2.mem\[57\]\[13\] _05122_ _05125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_16_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06276__B1 _01663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09249_ _04254_ u2.mem\[26\]\[1\] _04290_ _04292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06276__C2 u2.mem\[176\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12260_ _00139_ clknet_leaf_72_clock u2.mem\[8\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09065__I0 _04174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11758__S _05848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11211_ _05511_ u2.mem\[150\]\[3\] _05502_ _05512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09765__A1 _04180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12191_ _00070_ clknet_leaf_252_clock u2.mem\[4\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07776__B1 _03156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11572__A1 _05411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09228__S _04270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput43 net43 driver_io[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_11142_ _05467_ _01136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07240__A2 _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08132__S _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11557__I _05605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10461__I _05029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11073_ _05339_ _05424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10024_ _04761_ _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_118_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11875__A2 _05926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07543__A3 _03013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08866__I _04014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_18_clock clknet_5_2_0_clock clknet_leaf_18_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06751__A1 u2.mem\[179\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06751__B2 u2.mem\[191\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11975_ _05970_ _05985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_3985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09540__I1 u2.mem\[33\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10686__I0 _05106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10926_ _05301_ u2.mem\[133\]\[2\] _05327_ _05330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12811__CLK clknet_leaf_184_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10857_ _05286_ _05287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_71_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13576_ _01455_ clknet_leaf_32_clock u2.mem\[194\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10788_ _05245_ _01004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_169_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12527_ _00406_ clknet_leaf_189_clock u2.mem\[25\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06806__A2 _02043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10636__I _05151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12961__CLK clknet_leaf_168_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12458_ _00337_ clknet_leaf_135_clock u2.mem\[20\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11668__S _05787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11409_ _05635_ u2.mem\[162\]\[5\] _05624_ _05636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12389_ _00268_ clknet_leaf_79_clock u2.mem\[16\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07767__B1 _03069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06950_ _02399_ _02429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_101_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07519__B1 _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input3_I col_select_a[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06881_ _02359_ _02360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08620_ _03878_ _03884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__12341__CLK clknet_leaf_94_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13467__CLK clknet_leaf_361_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08551_ _03814_ u2.mem\[10\]\[7\] _03840_ _03844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07502_ u2.mem\[45\]\[7\] _02866_ _02867_ u2.mem\[34\]\[7\] _02974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_39_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10677__I0 _05097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07298__A2 _02586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08482_ _03657_ _03544_ _03775_ _03798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_35_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07433_ _02901_ _02902_ _02903_ _02906_ _02907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_22_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07364_ _02576_ _02839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09295__I0 _04260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08217__S _03618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09103_ _04198_ _00366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09400__I _04166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06258__B1 _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06315_ _01815_ _01816_ _01817_ _01818_ _01819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_31_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07295_ u2.mem\[28\]\[3\] _02580_ _02582_ u2.mem\[31\]\[3\] _02771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09034_ _04150_ _04151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06246_ u2.mem\[171\]\[1\] _01610_ _01615_ u2.mem\[157\]\[1\] _01752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08016__I mem_address_trans\[4\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07470__A2 _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11578__S _05739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06177_ _01683_ _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07758__B1 _03054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09048__S _04155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07222__A2 _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08270__I1 u2.mem\[4\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10281__I _04922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06430__B1 _01929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09936_ _04687_ u2.mem\[42\]\[2\] _04719_ _04722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06981__A1 _02439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09867_ _04675_ _00653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08818_ _03936_ u2.mem\[16\]\[14\] _04005_ _04008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09798_ _04612_ u2.mem\[38\]\[14\] _04633_ _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06733__A1 u2.mem\[188\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06733__B2 u2.mem\[175\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07930__B1 _02555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08749_ _03911_ u2.mem\[15\]\[3\] _03962_ _03966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10668__I0 _05126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11760_ _05837_ u2.mem\[184\]\[5\] _05848_ _05855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07289__A2 _02537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10711_ _03903_ _05172_ _05195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11691_ _05792_ u2.mem\[180\]\[2\] _05810_ _05813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10657__S _05162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13430_ _01309_ clknet_leaf_351_clock u2.mem\[175\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10642_ _05155_ _00948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09286__I0 _04246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06934__I _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_23_0_clock_I clknet_4_11_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13361_ _01240_ clknet_leaf_369_clock u2.mem\[163\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10573_ _05094_ _05113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_158_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07997__B1 _03459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12312_ _00191_ clknet_leaf_117_clock u2.mem\[11\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12214__CLK clknet_leaf_72_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13292_ _01171_ clknet_leaf_382_clock u2.mem\[152\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06264__A3 _01769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11488__S _05683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12243_ _00122_ clknet_leaf_75_clock u2.mem\[7\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12174_ _00053_ clknet_leaf_232_clock u2.mem\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07213__A2 _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10191__I _04864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11125_ _05456_ _01130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11056_ _05380_ u2.mem\[141\]\[0\] _05413_ _05414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10007_ _04681_ u2.mem\[44\]\[0\] _04762_ _04763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06724__A1 u2.mem\[171\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06724__B2 u2.mem\[157\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10659__I0 _05117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11958_ _05909_ u2.mem\[194\]\[2\] _05975_ _05976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09421__S _04396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10909_ _05320_ _01050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10567__S _05104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11889_ u2.mem\[192\]\[5\] _03510_ _05932_ _05936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_232_clock_I clknet_5_28_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13559_ _01438_ clknet_leaf_33_clock u2.mem\[193\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_146_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07988__B1 _02629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06100_ _01596_ _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10831__I0 u2.mem\[63\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07080_ _02558_ _02559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06031_ _01531_ _01534_ _01539_ _01516_ _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_172_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12707__CLK clknet_leaf_65_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11387__I1 u2.mem\[161\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07982_ _03442_ _03443_ _03444_ _03445_ _03446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_101_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06963__A1 _02441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12857__CLK clknet_5_13_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06933_ _02386_ _02412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_45_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09721_ _04583_ u2.mem\[37\]\[5\] _04580_ _04584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08500__S _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09652_ _04494_ u2.mem\[35\]\[13\] _04537_ _04539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06864_ _01984_ _02007_ _02009_ row_select_trans\[1\].data_sync _02343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_41_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07912__B1 _02426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08603_ _03873_ _00191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09583_ _04499_ _00545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06795_ u2.mem\[149\]\[4\] _02176_ _02177_ u2.mem\[175\]\[4\] _02276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06191__A2 _01665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11861__S _05918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08534_ _03657_ _03725_ _03775_ _03834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_23_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09331__S _04336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08465_ _03788_ _00138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07416_ _02517_ _02890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12237__CLK clknet_leaf_226_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08396_ _03745_ _00112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07347_ u2.mem\[43\]\[4\] _02820_ _02821_ u2.mem\[20\]\[4\] _02822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_17_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07443__A2 _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07278_ u2.mem\[53\]\[3\] _02476_ _02483_ u2.mem\[56\]\[3\] _02754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09017_ _04137_ _00341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06229_ u2.mem\[145\]\[1\] _01640_ _01734_ u2.mem\[177\]\[1\] _01735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06403__B1 _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09919_ _04709_ u2.mem\[41\]\[12\] _04710_ _04711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_150_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08410__S _03753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_181_clock_I clknet_5_27_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12930_ _00809_ clknet_leaf_151_clock u2.mem\[50\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10889__I0 _05307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06929__I _02407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06706__A1 _02184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12861_ _00740_ clknet_leaf_203_clock u2.mem\[46\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11812_ _05887_ _05888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12792_ _00671_ clknet_leaf_339_clock u2.mem\[41\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11743_ _05835_ u2.mem\[183\]\[4\] _05839_ _05845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07682__A2 _03082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11674_ _05790_ u2.mem\[179\]\[1\] _05801_ _05803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13162__CLK clknet_leaf_279_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13413_ _01292_ clknet_5_5_0_clock u2.mem\[172\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11066__I0 _05392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10625_ _05145_ _00941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13344_ _01223_ clknet_leaf_6_clock u2.mem\[160\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10556_ _04997_ _05101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10487_ _05009_ u2.mem\[55\]\[7\] _05056_ _05060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13275_ _01154_ clknet_leaf_9_clock u2.mem\[149\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11369__I1 u2.mem\[160\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09187__A2 _03774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12226_ _00105_ clknet_leaf_241_clock u2.mem\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11946__S _05965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12157_ _00036_ clknet_leaf_213_clock u2.mem\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07737__A3 _03200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06945__A1 _02377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11108_ _05424_ u2.mem\[144\]\[1\] _05445_ _05447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12088_ row_col_select_trans.A clknet_leaf_303_clock row_col_select_trans.data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11039_ _04334_ _05402_ _05403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_83_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06580_ _02064_ _02028_ _02065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_75_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09498__I0 _04360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09151__S _04226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13505__CLK clknet_leaf_333_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10297__S _04938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_383_clock_I clknet_5_0_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08250_ _03557_ u2.mem\[4\]\[5\] _03639_ _03641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06574__I _02058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07673__A2 _03141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07201_ u2.mem\[9\]\[1\] _02572_ _02577_ u2.mem\[25\]\[1\] _02679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_21_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10096__I _04819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08181_ _03598_ _00044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07132_ _02587_ _02588_ _02488_ _02562_ _02611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__09670__I0 _04473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07063_ _02541_ _02542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11509__A1 _04248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06014_ u2.driver_mem\[7\] _01508_ _01523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_99_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06936__A1 _02414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08230__S _03623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07965_ u2.mem\[58\]\[15\] _03277_ _03278_ u2.mem\[36\]\[15\] _03429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_151_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11655__I _05667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13035__CLK clknet_leaf_264_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09704_ _04570_ u2.mem\[37\]\[1\] _04567_ _04571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06916_ _02394_ _02395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_112_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09725__I1 u2.mem\[37\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07896_ _03358_ _03359_ _03360_ _03361_ _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__11532__I1 u2.mem\[170\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09635_ _04529_ _00567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06847_ u2.mem\[148\]\[5\] _02128_ _02130_ u2.mem\[152\]\[5\] _02327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_3_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09489__I0 _04391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09566_ _04487_ u2.mem\[33\]\[10\] _04483_ _04488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06778_ _02256_ _02257_ _02258_ _02259_ _02260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__13185__CLK clknet_leaf_294_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09061__S _04168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08517_ _03822_ _00156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11296__I0 _05556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09497_ _04444_ _00514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09996__S _04755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10000__S _04755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08448_ _03663_ u2.mem\[8\]\[1\] _03777_ _03779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07664__A2 _03132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_128_clock_I clknet_5_15_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08379_ _03688_ u2.mem\[6\]\[7\] _03732_ _03736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11748__A1 _04223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10410_ _05013_ _00858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11390_ _05622_ _01229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09661__I0 _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10341_ _04889_ u2.mem\[52\]\[1\] _04966_ _04968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10734__I _03686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13060_ _00939_ clknet_leaf_29_clock u2.mem\[58\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10272_ _04922_ _04928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_152_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11766__S _05857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12011_ net27 clknet_2_1__leaf_clock_a mem_address_trans\[3\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_152_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06659__I _02143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12402__CLK clknet_leaf_171_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13528__CLK clknet_leaf_332_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12913_ _00792_ clknet_leaf_163_clock u2.mem\[49\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12844_ _00723_ clknet_leaf_215_clock u2.mem\[45\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12775_ _00654_ clknet_leaf_141_clock u2.mem\[40\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11726_ _05834_ _01353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06312__C1 _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11657_ _05791_ _01327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10845__S _05278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10608_ _05130_ _05136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_127_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09652__I0 _04494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11588_ _05747_ _05748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_156_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13327_ _01206_ clknet_leaf_0_clock u2.mem\[158\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10539_ _05023_ u2.mem\[56\]\[13\] _05088_ _05090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08080__A2 _03528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06091__A1 _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08114__I _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13258_ _01137_ clknet_leaf_285_clock u2.mem\[146\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11676__S _05801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13058__CLK clknet_leaf_250_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12209_ _00088_ clknet_leaf_252_clock u2.mem\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10580__S _05113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13189_ _01068_ clknet_leaf_296_clock u2.mem\[135\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11911__A1 _03534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07040__B1 _02518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07186__A4 _02663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06394__A2 _01889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07750_ u2.mem\[50\]\[11\] _03113_ _03114_ u2.mem\[51\]\[11\] _03218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_81_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06569__I _02053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12082__CLK clknet_leaf_380_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06701_ _02103_ _02185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07681_ u2.mem\[17\]\[9\] _03079_ _03080_ u2.mem\[24\]\[9\] _03151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_168_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06146__A2 _01630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08391__I0 _03709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09420_ _04398_ _00483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06632_ _02116_ _02117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08784__I _03987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09351_ _04335_ _04351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06563_ u2.mem\[180\]\[0\] _02043_ _02047_ u2.mem\[150\]\[0\] _02048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10819__I _05252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08302_ _03677_ _00086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09282_ _03747_ _04247_ _04310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_55_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06494_ u2.mem\[0\]\[15\] _01980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08233_ _03628_ _03629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10755__S _05223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08164_ _03552_ u2.mem\[2\]\[3\] _03585_ _03589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09643__I0 _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07115_ _02593_ _02594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_174_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_146_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07949__A3 _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11450__I0 _05633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08095_ _03483_ _03539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06082__A1 _01586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07046_ _02524_ _02525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10490__S _05061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input41_I row_select_a[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08997_ _04120_ _04121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07084__B _02417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08895__S _04056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07948_ u2.mem\[6\]\[14\] _02622_ _02624_ u2.mem\[47\]\[14\] _03413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_54_clock_I clknet_5_12_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09323__A2 _04334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07879_ u2.mem\[58\]\[13\] _03277_ _03278_ u2.mem\[36\]\[13\] _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_44_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12575__CLK clknet_leaf_184_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08382__I0 _03692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09618_ _04519_ _00560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10890_ _05308_ _01043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09549_ _04144_ _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12560_ _00439_ clknet_leaf_159_clock u2.mem\[27\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07637__A2 _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07103__I _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06845__B1 _02134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11511_ _05663_ u2.mem\[169\]\[0\] _05700_ _05701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_279_clock_I clknet_5_23_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12491_ _00370_ clknet_leaf_177_clock u2.mem\[23\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06942__I _02362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11442_ _05623_ u2.mem\[165\]\[0\] _05655_ _05656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09634__I0 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08135__S _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08437__I1 u2.mem\[7\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11373_ _05593_ u2.mem\[160\]\[4\] _05607_ _05613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10324_ _04957_ _00828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13112_ _00991_ clknet_leaf_45_clock u2.mem\[61\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07270__B1 _02452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_331_clock_I clknet_5_18_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10255_ _04917_ _00799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_363_clock clknet_5_4_0_clock clknet_leaf_363_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13043_ _00922_ clknet_leaf_31_clock u2.mem\[57\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08869__I _03713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13350__CLK clknet_leaf_7_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10186_ _04872_ _00775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12918__CLK clknet_leaf_87_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06781__C1 u2.mem\[181\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_378_clock clknet_5_0_0_clock clknet_leaf_378_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_75_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08373__I0 _03675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07876__A2 _02493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10180__I0 _04790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12827_ _00706_ clknet_leaf_184_clock u2.mem\[44\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_301_clock clknet_5_21_0_clock clknet_leaf_301_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08125__I0 _03561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12758_ _00637_ clknet_leaf_71_clock u2.mem\[39\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07628__A2 _03017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09873__I0 _04612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11709_ _05796_ u2.mem\[181\]\[4\] _05817_ _05823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11680__I0 _05796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06836__B1 _02105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12689_ _00568_ clknet_leaf_155_clock u2.mem\[35\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06300__A2 _01676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_316_clock clknet_5_17_0_clock clknet_leaf_316_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_163_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09625__I0 _04467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11432__I0 _05629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10374__I _04117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06064__A1 _01547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12448__CLK clknet_leaf_168_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07261__B1 _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08920_ _04075_ _00306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08779__I mem_address_trans\[4\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11735__I1 u2.mem\[183\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08851_ _04031_ _00281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06367__A2 _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07802_ _02469_ _03269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08782_ mem_address_trans\[7\].data_sync _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05994_ u2.select_mem_row\[1\] u2.select_mem_col\[1\] _01502_ _01503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09604__S _04511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07733_ u2.mem\[39\]\[10\] _03090_ _03091_ u2.mem\[48\]\[10\] _03202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11499__I0 _05668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07316__A1 u2.mem\[40\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06119__A2 _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07316__B2 u2.mem\[30\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08364__I0 _03656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07664_ u2.mem\[61\]\[9\] _03132_ _03133_ u2.mem\[63\]\[9\] _03134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09403_ _04386_ _00478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06615_ _02028_ _02060_ _02100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_164_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07595_ _03058_ _03061_ _03064_ _03065_ _03066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_111_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08116__I0 _03554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09334_ _04260_ u2.mem\[28\]\[4\] _04341_ _04342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06546_ _02005_ _02031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08019__I mem_address_trans\[1\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09864__I0 _04599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_280_clock_I clknet_5_23_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09265_ _04269_ u2.mem\[26\]\[8\] _04300_ _04301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10485__S _05056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06477_ u2.mem\[194\]\[11\] _01946_ _01967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13223__CLK clknet_leaf_301_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08216_ _03619_ _00058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09196_ _04254_ u2.mem\[25\]\[1\] _04252_ _04255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11423__I0 _05635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07079__B _02430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08147_ _03532_ _03577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08078_ data_in_trans\[12\].data_sync _03527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13373__CLK clknet_leaf_371_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07029_ _02507_ _02508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10040_ _04716_ u2.mem\[44\]\[15\] _04777_ _04781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06430__C _01914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09514__S _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07307__A1 _02767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11991_ _00003_ clknet_leaf_331_clock u2.mem\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10942_ _05340_ u2.mem\[134\]\[1\] _05337_ _05341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10873_ _05296_ _05297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_32_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12612_ _00491_ clknet_leaf_82_clock u2.mem\[30\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09855__I0 _04586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12543_ _00422_ clknet_leaf_189_clock u2.mem\[26\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11662__I0 _05794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10395__S _05002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06294__A1 u2.mem\[144\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06294__B2 u2.mem\[182\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12474_ _00353_ clknet_leaf_127_clock u2.mem\[21\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11425_ _05605_ _05645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06046__A1 _01547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07243__B1 _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11356_ _05602_ _01215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10307_ _04893_ u2.mem\[51\]\[3\] _04944_ _04948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08599__I _03855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12740__CLK clknet_leaf_24_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11287_ _05560_ _01188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13026_ _00905_ clknet_leaf_265_clock u2.mem\[56\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10238_ _04904_ u2.mem\[49\]\[8\] _04905_ _04906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06349__A2 _01778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10169_ _03477_ mem_address_trans\[5\].data_sync _04861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07008__I _02486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12890__CLK clknet_leaf_57_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_240_clock clknet_5_25_0_clock clknet_leaf_240_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_47_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12120__CLK clknet_leaf_348_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13246__CLK clknet_leaf_289_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06400_ u2.mem\[144\]\[5\] _01670_ _01672_ u2.mem\[182\]\[5\] _01902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07380_ _02845_ _02848_ _02851_ _02854_ _02855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_91_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09846__I0 _04573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06331_ u2.mem\[173\]\[3\] _01720_ _01722_ u2.mem\[185\]\[3\] _01835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11653__I0 _05786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07678__I _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09050_ data_in_trans\[11\].data_sync _04163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06285__A1 u2.mem\[145\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06285__B2 u2.mem\[163\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06262_ u2.mem\[189\]\[1\] _01649_ _01651_ u2.mem\[176\]\[1\] u2.mem\[172\]\[1\]
+ _01653_ _01768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_30_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13396__CLK clknet_leaf_327_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08001_ _03460_ _03463_ _03464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06193_ _01616_ _01607_ _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08026__A2 _03486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07234__B1 _02483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08503__S _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09952_ _04703_ u2.mem\[42\]\[9\] _04729_ _04731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08903_ _04064_ _00300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11988__CLK clknet_leaf_380_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09883_ _04685_ u2.mem\[41\]\[1\] _04683_ _04686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_227_clock_I clknet_5_22_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08834_ _04019_ u2.mem\[17\]\[2\] _04015_ _04020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08765_ _03927_ u2.mem\[15\]\[10\] _03972_ _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08337__I0 _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06760__A2 _02185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_208_clock clknet_5_30_0_clock clknet_leaf_208_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07716_ _03169_ _03174_ _03179_ _03184_ _03185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08696_ _03934_ u2.mem\[13\]\[13\] _03932_ _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07647_ _02500_ _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07578_ u2.mem\[14\]\[8\] _02892_ _02893_ u2.mem\[12\]\[8\] _03049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09837__I0 _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12613__CLK clknet_leaf_92_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09317_ _04283_ u2.mem\[27\]\[14\] _04328_ _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11644__I0 _05754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06529_ _01998_ _02014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06276__A1 u2.mem\[189\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07588__I _02541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09248_ _04291_ _00418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06276__B2 u2.mem\[180\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08017__A2 mem_address_trans\[5\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09179_ _04242_ _00398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12763__CLK clknet_leaf_219_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07225__B1 _02639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11210_ _05510_ _05511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09765__A2 _04542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12190_ _00069_ clknet_leaf_267_clock u2.mem\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11572__A2 _05729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11141_ _05466_ u2.mem\[146\]\[2\] _05462_ _05467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput44 net44 driver_io[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_89_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13119__CLK clknet_leaf_257_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11072_ _05423_ _01110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10023_ _04771_ _00713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12143__CLK clknet_leaf_239_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11573__I _05738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13269__CLK clknet_leaf_384_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06751__A2 _02150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11088__A1 _04417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11974_ _05984_ _01451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09043__I _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10925_ _05329_ _01057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11883__I0 u2.mem\[192\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09828__I0 _04602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10856_ _05285_ _05276_ _05286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13575_ _01454_ clknet_leaf_33_clock u2.mem\[194\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10787_ _05218_ u2.mem\[62\]\[10\] _05242_ _05245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08500__I0 _03810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12526_ _00405_ clknet_leaf_198_clock u2.mem\[25\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_176_clock_I clknet_5_27_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12457_ _00336_ clknet_leaf_128_clock u2.mem\[20\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09419__S _04396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11408_ _05516_ _05635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06019__B2 _01516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12388_ _00267_ clknet_leaf_79_clock u2.mem\[16\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11339_ _05591_ u2.mem\[158\]\[3\] _05585_ _05592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09218__I _04251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08567__I0 _03830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07519__B2 u2.mem\[12\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13009_ _00888_ clknet_leaf_253_clock u2.mem\[55\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06880_ _02358_ _02359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08550_ _03843_ _00168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06577__I _02061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10126__I0 _04813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12636__CLK clknet_leaf_215_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07501_ _01945_ _02784_ _02952_ _02973_ _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_35_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08481_ _03655_ _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07432_ u2.mem\[57\]\[5\] _02904_ _02905_ u2.mem\[41\]\[5\] _02906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_194_clock clknet_5_31_0_clock clknet_leaf_194_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09819__I0 _04589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11626__I0 _05750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07363_ _02571_ _02838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09295__I1 u2.mem\[27\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12786__CLK clknet_leaf_338_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09102_ _04167_ u2.mem\[22\]\[12\] _04197_ _04198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06258__A1 u2.mem\[180\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07455__B1 _02928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06258__B2 u2.mem\[150\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06314_ u2.mem\[172\]\[3\] _01654_ _01664_ u2.mem\[180\]\[3\] _01818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07294_ u2.mem\[9\]\[3\] _02572_ _02577_ u2.mem\[25\]\[3\] _02770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_149_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09033_ data_in_trans\[7\].data_sync _04150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06245_ u2.mem\[167\]\[1\] _01749_ _01750_ u2.mem\[183\]\[1\] _01751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12016__CLK clknet_leaf_315_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07207__B1 _02591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09329__S _04336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06176_ _01622_ _01641_ _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11658__I _05670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_132_clock clknet_5_15_0_clock clknet_leaf_132_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_131_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06430__A1 u2.mem\[193\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09935_ _04721_ _00675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06430__B2 u2.mem\[192\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08032__I _03492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_378_clock_I clknet_5_0_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08558__I0 _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12166__CLK clknet_leaf_79_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09866_ _04602_ u2.mem\[40\]\[11\] _04671_ _04675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06718__C1 _02019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08817_ _04007_ _00271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_147_clock clknet_5_13_0_clock clknet_leaf_147_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_86_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09797_ _04635_ _00623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11393__I _05624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06733__A2 _02185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07092__B _02546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08748_ _03965_ _00244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10117__I0 _04804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13561__CLK clknet_leaf_32_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11865__I0 _05909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10668__I1 u2.mem\[59\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08679_ _03904_ _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10938__S _05337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_9_0_clock clknet_3_4_0_clock clknet_4_9_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__08730__I0 _03929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10710_ _04986_ _05194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08408__S _03753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11690_ _05812_ _01339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10641_ _05099_ u2.mem\[59\]\[2\] _05152_ _05155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10737__I _03690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09286__I1 u2.mem\[27\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13360_ _01239_ clknet_leaf_371_clock u2.mem\[163\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10572_ _03690_ _05112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12311_ _00190_ clknet_leaf_115_clock u2.mem\[11\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_166_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13291_ _01170_ clknet_leaf_378_clock u2.mem\[152\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_5_27_0_clock_I clknet_4_13_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12242_ _00121_ clknet_leaf_239_clock u2.mem\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07749__A1 _03212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12173_ _00052_ clknet_leaf_231_clock u2.mem\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09038__I _04153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11124_ _05426_ u2.mem\[145\]\[2\] _05453_ _05456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_150_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08549__I0 _03812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13091__CLK clknet_leaf_26_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11055_ _05412_ _05413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_42_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10006_ _04761_ _04762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_49_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06724__A2 _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10108__I0 _04795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11957_ _05971_ _05975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_166_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08721__I0 _03920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06488__A1 _01973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10908_ _05294_ u2.mem\[132\]\[0\] _05319_ _05320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_75_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11888_ _05935_ _01414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11608__I0 _05746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10839_ _03477_ _03984_ _05274_ _05275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_60_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12039__CLK clknet_2_2__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13558_ _01437_ clknet_leaf_16_clock u2.mem\[193\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12509_ _00388_ clknet_leaf_196_clock u2.mem\[24\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10583__S _05113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10831__I1 _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13489_ _01368_ clknet_leaf_306_clock u2.mem\[185\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06030_ _01504_ _01536_ _01538_ _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06660__A1 _02005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12189__CLK clknet_leaf_267_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06412__A1 _01911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07981_ u2.mem\[28\]\[15\] _03307_ _03308_ u2.mem\[31\]\[15\] _03445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06963__A2 _02429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_64_clock clknet_5_9_0_clock clknet_leaf_64_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09720_ _04582_ _04583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06932_ u2.mem\[40\]\[0\] _02403_ _02410_ u2.mem\[30\]\[0\] _02411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07691__I _02623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09651_ _04538_ _00574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08704__A3 _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06863_ col_select_trans\[5\].data_sync _02024_ _02016_ col_select_trans\[4\].data_sync
+ _02342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_83_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07912__A1 u2.mem\[27\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08602_ _03828_ u2.mem\[11\]\[13\] _03871_ _03873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08960__I0 _04017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09582_ _04498_ u2.mem\[33\]\[15\] _04492_ _04499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06794_ u2.mem\[166\]\[4\] _02096_ _02098_ u2.mem\[161\]\[4\] u2.mem\[159\]\[4\]
+ _02174_ _02275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
Xclkbuf_leaf_79_clock clknet_5_8_0_clock clknet_leaf_79_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06191__A3 _01678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08533_ _03833_ _00161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06100__I _01596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10758__S _05223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08712__I0 _03911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11941__I _05949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06479__A1 _01966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07676__B1 _03075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08464_ _03692_ u2.mem\[8\]\[8\] _03787_ _03788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08228__S _03623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07415_ _02513_ _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08395_ _03718_ u2.mem\[6\]\[14\] _03742_ _03745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07346_ _02507_ _02821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08027__I _03487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10822__I1 _03520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07277_ u2.mem\[54\]\[3\] _02650_ _02651_ u2.mem\[55\]\[3\] _02753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_17_clock clknet_5_2_0_clock clknet_leaf_17_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09016_ _04136_ u2.mem\[21\]\[3\] _04124_ _04137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06228_ _01583_ _01734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07087__B _02485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06159_ _01612_ _01665_ _01591_ _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__08898__S _04061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06403__A1 u2.mem\[191\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09918_ _04682_ _04710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_77_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08156__A1 _03479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_124_clock_I clknet_5_15_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09849_ _04665_ _00645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06706__A2 _02188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12860_ _00739_ clknet_leaf_215_clock u2.mem\[46\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12951__CLK clknet_leaf_147_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11811_ _04333_ _05886_ _05887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__06010__I _01503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12791_ _00670_ clknet_leaf_339_clock u2.mem\[41\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11742_ _05844_ _01359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08138__S _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10510__I0 _04987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13307__CLK clknet_leaf_370_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11673_ _05802_ _01332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13412_ _01291_ clknet_leaf_358_clock u2.mem\[172\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10624_ _05119_ u2.mem\[58\]\[11\] _05141_ _05145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11499__S _05692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13343_ _01222_ clknet_leaf_2_clock u2.mem\[160\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12331__CLK clknet_leaf_234_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10813__I1 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10555_ _05100_ _00916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_49_clock_I clknet_5_7_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13457__CLK clknet_leaf_325_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13274_ _01153_ clknet_leaf_7_clock u2.mem\[149\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10486_ _05059_ _00888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11298__I _05442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12225_ _00104_ clknet_leaf_242_clock u2.mem\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10577__I0 _05115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12481__CLK clknet_leaf_172_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12156_ _00035_ clknet_leaf_219_clock u2.mem\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06945__A2 _02391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11107_ _05446_ _01122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12087_ net36 clknet_2_3__leaf_clock_a row_col_select_trans.A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11038_ _05275_ _05402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_42_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08400__I _03483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11962__S _05975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07370__A2 _02682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11829__I0 _05868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09498__I1 u2.mem\[32\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12989_ _00868_ clknet_leaf_274_clock u2.mem\[54\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_166_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07658__B1 _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10501__I0 _05023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09231__I _04251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_326_clock_I clknet_5_16_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10377__I _04988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06330__B1 _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07200_ u2.mem\[29\]\[1\] _02559_ _02564_ u2.mem\[11\]\[1\] _02678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_32_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08180_ _03568_ u2.mem\[2\]\[10\] _03595_ _03598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07131_ _02609_ _02610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10804__I1 _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09670__I1 u2.mem\[36\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07686__I _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07062_ _02477_ _02529_ _02530_ _02512_ _02541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__06633__A1 u2.mem\[144\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12824__CLK clknet_leaf_129_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11509__A2 _05690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06013_ _01511_ _01522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06397__B1 _01714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06936__A2 _02350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10840__I _05275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07964_ u2.mem\[53\]\[15\] _03274_ _03275_ u2.mem\[56\]\[15\] _03428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12974__CLK clknet_leaf_271_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09703_ _04569_ _04570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06915_ _02362_ _02394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08310__I _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07895_ u2.mem\[28\]\[13\] _03307_ _03308_ u2.mem\[31\]\[13\] _03361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09634_ _04476_ u2.mem\[35\]\[5\] _04527_ _04529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07897__B1 _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06846_ u2.mem\[153\]\[5\] _02136_ _02137_ u2.mem\[160\]\[5\] _02326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_55_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12204__CLK clknet_leaf_271_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09565_ _04160_ _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06777_ u2.mem\[145\]\[3\] _02081_ _02091_ u2.mem\[177\]\[3\] _02259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_55_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11671__I _05800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08516_ _03821_ u2.mem\[9\]\[10\] _03817_ _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07649__B1 _03042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11296__I1 u2.mem\[155\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09496_ _04356_ u2.mem\[32\]\[0\] _04443_ _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07113__A2 _02586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08447_ _03778_ _00130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12354__CLK clknet_leaf_162_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08378_ _03735_ _00104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11748__A2 _05847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07329_ u2.mem\[3\]\[4\] _02803_ _02749_ _02804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_109_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_50_clock_I clknet_5_7_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11112__S _05445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10340_ _04967_ _00834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10271_ _04927_ _00805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12010_ mem_address_trans\[2\].A clknet_leaf_315_clock mem_address_trans\[2\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06388__B1 _01732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06927__A2 _02400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10750__I _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_275_clock_I clknet_5_23_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11782__S _05866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12912_ _00791_ clknet_leaf_162_clock u2.mem\[49\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12843_ _00722_ clknet_leaf_214_clock u2.mem\[45\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12774_ _00653_ clknet_leaf_76_clock u2.mem\[40\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09051__I _04163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07104__A2 _02580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_3_6_0_clock clknet_0_clock clknet_3_6_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_37_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11987__A2 _05972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11725_ _05833_ u2.mem\[182\]\[3\] _05827_ _05834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06312__B1 _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06312__C2 u2.mem\[181\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09986__I _04739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06863__A1 col_select_trans\[5\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11656_ _05790_ u2.mem\[178\]\[1\] _05788_ _05791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10607_ _05135_ _00933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11587_ _04393_ _05729_ _05747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_122_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11022__S _05381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10798__I0 _05229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13326_ _01205_ clknet_leaf_324_clock u2.mem\[157\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06615__A1 _02028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10538_ _05089_ _00910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06091__A2 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13257_ _01136_ clknet_leaf_286_clock u2.mem\[146\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10469_ _05049_ _00881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12208_ _00087_ clknet_leaf_241_clock u2.mem\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11211__I1 u2.mem\[150\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06379__B1 _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13188_ _01067_ clknet_leaf_291_clock u2.mem\[134\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11911__A2 _05929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12139_ _00018_ clknet_leaf_230_clock u2.mem\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06700_ u2.mem\[171\]\[1\] _02065_ _02067_ u2.mem\[157\]\[1\] _02183_ _02184_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_42_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07680_ u2.mem\[23\]\[9\] _03148_ _03149_ u2.mem\[22\]\[9\] _03150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_93_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10722__I0 _05202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06631_ _02015_ _02046_ _02116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12377__CLK clknet_leaf_114_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09350_ _04350_ _00461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10101__S _04820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06562_ _02045_ _02046_ _02047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09340__I0 _04267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08301_ _03675_ u2.mem\[5\]\[4\] _03676_ _03677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09281_ _04309_ _00433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06493_ u2.mem\[194\]\[15\] _01979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_33_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08232_ mem_address_trans\[1\].data_sync mem_address_trans\[0\].data_sync _03628_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08506__S _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08163_ _03588_ _00036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10789__I0 _05220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07114_ _02447_ _02449_ _02458_ _02575_ _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_118_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06606__A1 _02080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08305__I _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11450__I1 u2.mem\[165\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08094_ _03491_ _03538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_8_0_clock clknet_4_4_0_clock clknet_5_8_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_109_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11867__S _05918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07045_ _02522_ _02523_ _02512_ _02450_ _02524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__10771__S _05232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08241__S _03634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08996_ _03900_ _03749_ _04120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_130_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input34_I mem_write_n_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13152__CLK clknet_leaf_260_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08040__I _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07084__C _02562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07947_ u2.mem\[8\]\[14\] _03326_ _03327_ u2.mem\[4\]\[14\] _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_25_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08975__I _04096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07878_ u2.mem\[53\]\[13\] _03274_ _03275_ u2.mem\[56\]\[13\] _03344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10713__I0 _05194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09617_ _04496_ u2.mem\[34\]\[14\] _04516_ _04519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06829_ _02305_ _02306_ _02307_ _02308_ _02309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_16_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10011__S _04762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09548_ _04475_ _00534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09331__I0 _04258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09800__S _04633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09479_ _04432_ _00508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10946__S _05337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11510_ _05699_ _05700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06845__A1 u2.mem\[194\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12490_ _00369_ clknet_leaf_127_clock u2.mem\[22\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11441_ _05654_ _05655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_7_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11372_ _05612_ _01221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13111_ _00990_ clknet_leaf_39_clock u2.mem\[61\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10323_ _04909_ u2.mem\[51\]\[10\] _04954_ _04957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10681__S _05174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09247__S _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09398__I0 _04382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13042_ _00921_ clknet_leaf_336_clock u2.mem\[57\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10254_ _04916_ u2.mem\[49\]\[13\] _04914_ _04917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08151__S _03573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10480__I _05050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10185_ _04795_ u2.mem\[48\]\[5\] _04870_ _04872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_65_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09046__I data_in_trans\[10\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06781__B1 _02034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06781__C2 _02038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10704__I0 _05124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12826_ _00705_ clknet_leaf_129_clock u2.mem\[43\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07089__A1 _02560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12757_ _00636_ clknet_leaf_71_clock u2.mem\[39\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09873__I1 u2.mem\[40\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11708_ _05822_ _01347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06836__A1 u2.mem\[188\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12688_ _00567_ clknet_leaf_157_clock u2.mem\[35\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11680__I1 u2.mem\[179\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11639_ _05780_ _01320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13025__CLK clknet_leaf_253_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11432__I1 u2.mem\[164\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11687__S _05810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13309_ _01188_ clknet_leaf_363_clock u2.mem\[155\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09389__I0 _04375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09157__S _04226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08850_ _04030_ u2.mem\[17\]\[7\] _04024_ _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07564__A2 _03033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07801_ u2.mem\[16\]\[12\] _03266_ _03267_ u2.mem\[33\]\[12\] _03268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08781_ mem_address_trans\[6\].data_sync _03985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_22_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05993_ row_col_select_trans.data_sync _01502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_78_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07732_ u2.mem\[5\]\[10\] _03155_ _03156_ u2.mem\[38\]\[10\] _03201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08795__I _03989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11499__I1 u2.mem\[168\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07663_ _02554_ _03133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_92_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09402_ _04384_ u2.mem\[29\]\[12\] _04385_ _04386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06614_ _02098_ _02099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07594_ u2.mem\[57\]\[8\] _02904_ _02905_ u2.mem\[41\]\[8\] _03065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_168_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07204__I _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09313__I0 _04278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09333_ _04335_ _04341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_146_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06545_ _02029_ _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11120__I0 _05420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09864__I1 u2.mem\[40\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_223_clock_I clknet_5_23_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06827__A1 u2.mem\[167\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09264_ _04289_ _04300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06827__B2 u2.mem\[183\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06476_ u2.mem\[0\]\[11\] _01966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08215_ _03563_ u2.mem\[3\]\[8\] _03618_ _03619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09195_ _04127_ _04254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08146_ _03576_ _00031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08035__I data_in_trans\[1\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11423__I1 u2.mem\[163\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07079__C _02506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13518__CLK clknet_leaf_354_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08077_ _03488_ _03526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07028_ _02447_ _02449_ _02488_ _02506_ _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_66_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11187__I0 _05466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11396__I _05504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12542__CLK clknet_leaf_198_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07555__A2 _03021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08979_ _04109_ _00331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11990_ _00002_ clknet_leaf_334_clock u2.mem\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_152_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07307__A2 _02772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10941_ _05339_ _05340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10872_ _05295_ _05276_ _05296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_71_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09304__I0 _04269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12611_ _00490_ clknet_leaf_85_clock u2.mem\[30\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09855__I1 u2.mem\[40\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12542_ _00421_ clknet_leaf_198_clock u2.mem\[26\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06953__I _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11811__A1 _04333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11662__I1 u2.mem\[178\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12473_ _00352_ clknet_leaf_169_clock u2.mem\[21\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12072__CLK clknet_leaf_379_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11424_ _05644_ _01241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13198__CLK clknet_leaf_293_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06046__A2 _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11355_ _05591_ u2.mem\[159\]\[3\] _05598_ _05602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07243__B2 u2.mem\[63\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10306_ _04947_ _00820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11286_ _05544_ u2.mem\[155\]\[0\] _05559_ _05560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_79_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13025_ _00904_ clknet_leaf_253_clock u2.mem\[56\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10237_ _04886_ _04905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_80_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09791__I0 _04602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10168_ _04860_ _00769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07010__A4 _02488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06754__B1 _02143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_172_clock_I clknet_5_26_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10099_ _04786_ u2.mem\[46\]\[1\] _04820_ _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09504__I _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09543__I0 _04471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06349__B _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12809_ _00688_ clknet_leaf_129_clock u2.mem\[42\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_163_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09846__I1 u2.mem\[40\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06330_ u2.mem\[154\]\[3\] _01698_ _01700_ u2.mem\[162\]\[3\] _01833_ _01834_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11653__I1 u2.mem\[178\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06285__A2 _01639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06261_ u2.mem\[190\]\[1\] _01703_ _01710_ u2.mem\[160\]\[1\] _01705_ u2.mem\[194\]\[1\]
+ _01767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__07482__A1 u2.mem\[37\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08000_ u2.active_mem\[7\] _03461_ _03462_ u2.active_mem\[6\] _03463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_102_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06192_ _01698_ _01699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_141_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_97_clock_I clknet_5_10_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12565__CLK clknet_leaf_105_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09951_ _04730_ _00682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11169__I0 _05460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08902_ _04037_ u2.mem\[18\]\[10\] _04061_ _04064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09882_ _04569_ _04685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10916__I0 _05305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09615__S _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08833_ _03666_ _04019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09782__I0 _04589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06745__B1 _02200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08764_ _03974_ _00251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09534__I0 _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09414__I _04393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07715_ _03180_ _03181_ _03182_ _03183_ _03184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08695_ _03713_ _03934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_2_3__f_clock_a clknet_0_clock_a clknet_2_3__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_54_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11880__S _05929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07646_ _02498_ _03116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11892__I1 _03512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07577_ u2.mem\[44\]\[8\] _02889_ _02890_ u2.mem\[42\]\[8\] _03048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_94_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10496__S _05061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_362_clock clknet_5_4_0_clock clknet_leaf_362_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_167_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09316_ _04330_ _00447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_374_clock_I clknet_5_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06528_ _02012_ _02013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12095__CLK clknet_leaf_338_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11644__I1 u2.mem\[177\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07068__A4 _02546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13340__CLK clknet_leaf_2_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09247_ _04246_ u2.mem\[26\]\[0\] _04290_ _04291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07473__A1 _02942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06459_ u2.mem\[193\]\[7\] _01942_ _01948_ u2.mem\[192\]\[7\] _01949_ _01953_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_31_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12908__CLK clknet_leaf_202_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09178_ _04167_ u2.mem\[24\]\[12\] _04241_ _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_377_clock clknet_5_0_0_clock clknet_leaf_377_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_147_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08017__A3 mem_address_trans\[6\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07225__A1 u2.mem\[27\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08129_ _03563_ u2.mem\[1\]\[8\] _03564_ _03565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06028__A2 _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13490__CLK clknet_leaf_307_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11120__S _05453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10080__I0 _04808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07776__A2 _03155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11140_ _05342_ _05466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_4_5_0_clock clknet_3_2_0_clock clknet_4_5_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_134_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_300_clock clknet_5_21_0_clock clknet_leaf_300_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_122_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11071_ _05420_ u2.mem\[142\]\[0\] _05422_ _05423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_1_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07109__I _02413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07528__A2 _02997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10022_ _04698_ u2.mem\[44\]\[7\] _04767_ _04771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09525__S _04458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09773__I0 _04576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06013__I _01511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06736__B1 _02099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11580__I0 _05715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_315_clock clknet_5_17_0_clock clknet_leaf_315_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09324__I _04335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09525__I0 _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11973_ _05216_ u2.mem\[194\]\[9\] _05980_ _05984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10924_ _05299_ u2.mem\[133\]\[1\] _05327_ _05329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12438__CLK clknet_leaf_102_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11883__I1 _03499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07700__A2 _03166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_2_3__f_clock_a_I clknet_0_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10855_ _04012_ _05285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_77_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13574_ _01453_ clknet_leaf_16_clock u2.mem\[194\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10786_ _05244_ _01003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07059__A4 _02417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12525_ _00404_ clknet_leaf_198_clock u2.mem\[25\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12588__CLK clknet_leaf_205_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_119_clock_I clknet_5_14_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12456_ _00335_ clknet_leaf_128_clock u2.mem\[20\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08604__S _03871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11407_ _05634_ _01234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12387_ _00266_ clknet_leaf_81_clock u2.mem\[16\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11030__S _05395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07767__A2 _03068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10071__I0 _04801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11338_ _05510_ _05591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12072__D data_in_trans\[11\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11269_ _05504_ _05548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07519__A2 _02892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09435__S _04406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13008_ _00887_ clknet_leaf_251_clock u2.mem\[55\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09234__I _04170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09516__I0 _04378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11323__I0 _05554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_1_0_clock_I clknet_4_0_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07500_ _02957_ _02962_ _02967_ _02972_ _02973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_63_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08480_ _03796_ _00145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13363__CLK clknet_leaf_374_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07431_ _02549_ _02905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07362_ u2.mem\[29\]\[4\] _02835_ _02836_ u2.mem\[11\]\[4\] _02837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_143_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11626__I1 u2.mem\[176\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09101_ _04181_ _04197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06313_ u2.mem\[189\]\[3\] _01650_ _01652_ u2.mem\[176\]\[3\] _01817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06258__A2 _01664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07293_ u2.mem\[29\]\[3\] _02559_ _02564_ u2.mem\[11\]\[3\] _02769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11004__I _05334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09032_ _04149_ _00344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06244_ _01624_ _01750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06175_ _01681_ _01682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07758__A2 _03053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08313__I data_in_trans\[7\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09934_ _04685_ u2.mem\[42\]\[1\] _04719_ _04721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09345__S _04346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09755__I0 _04609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09865_ _04674_ _00652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06718__B1 _02012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11562__I0 _05711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06718__C2 u2.mem\[189\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08816_ _03934_ u2.mem\[16\]\[13\] _04005_ _04007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09796_ _04609_ u2.mem\[38\]\[13\] _04633_ _04635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07391__B1 _02824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09507__I0 _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07930__A2 _02553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08747_ _03909_ u2.mem\[15\]\[2\] _03962_ _03965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07092__C _02443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08678_ _03691_ _03922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11865__I1 u2.mem\[191\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07629_ _02431_ _03099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07694__A1 _03140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12730__CLK clknet_leaf_47_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10640_ _05154_ _00947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06436__C _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06249__A2 _01751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_120_clock_I clknet_5_14_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10954__S _05336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10571_ _05111_ _00921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12310_ _00189_ clknet_leaf_97_clock u2.mem\[11\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07997__A2 _03458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13290_ _01169_ clknet_leaf_368_clock u2.mem\[151\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06008__I _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12880__CLK clknet_5_24_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12241_ _00120_ clknet_leaf_240_clock u2.mem\[7\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07749__A2 _03213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08223__I _03607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12172_ _00051_ clknet_leaf_231_clock u2.mem\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11785__S _05866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11123_ _05455_ _01129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12110__CLK clknet_leaf_381_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13236__CLK clknet_leaf_287_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09746__I0 _04602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11054_ _05411_ _05402_ _05412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_27_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11553__I0 _05717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06709__B1 _02192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_254_clock clknet_5_19_0_clock clknet_leaf_254_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_103_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10005_ _04334_ _04760_ _04761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09054__I data_in_trans\[12\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12260__CLK clknet_leaf_72_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13386__CLK clknet_leaf_323_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_45_clock_I clknet_5_6_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11305__I0 _05550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07134__B1 _02612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11956_ _05974_ _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_269_clock clknet_5_23_0_clock clknet_leaf_269_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10907_ _05318_ _05319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_11887_ u2.mem\[192\]\[4\] _03506_ _05932_ _05935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10838_ _05273_ mem_address_trans\[7\].data_sync _05274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__11608__I1 u2.mem\[175\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10864__S _05287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13557_ _01436_ clknet_leaf_16_clock u2.mem\[193\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10769_ _05200_ u2.mem\[62\]\[2\] _05232_ _05235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07988__A2 _02627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_173_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12508_ _00387_ clknet_leaf_195_clock u2.mem\[24\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13488_ _01367_ clknet_leaf_314_clock u2.mem\[184\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12439_ _00318_ clknet_leaf_119_clock u2.mem\[19\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10663__I _05151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06660__A2 _02125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_207_clock clknet_5_30_0_clock clknet_leaf_207_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_12_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06948__B1 _02426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11695__S _05809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_322_clock_I clknet_5_16_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06412__A2 _01912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07980_ u2.mem\[9\]\[15\] _03304_ _03305_ u2.mem\[25\]\[15\] _03444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_138_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12603__CLK clknet_leaf_214_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06931_ _02409_ _02410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06963__A3 _02416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11494__I _05605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09650_ _04491_ u2.mem\[35\]\[12\] _04537_ _04538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06862_ col_select_trans\[5\].data_sync _02025_ _02341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_94_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_0_clock clock clknet_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06176__A1 _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08601_ _03872_ _00190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08960__I1 u2.mem\[20\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07912__A2 _02420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09581_ _04176_ _04498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06793_ u2.mem\[177\]\[4\] _02091_ _02088_ u2.mem\[193\]\[4\] _02274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_97_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08532_ _03832_ u2.mem\[9\]\[15\] _03826_ _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12753__CLK clknet_leaf_247_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08712__I1 u2.mem\[14\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08463_ _03776_ _03787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06479__A2 _01955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07414_ _02882_ _02885_ _02886_ _02887_ _02888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_168_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08394_ _03744_ _00111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08308__I data_in_trans\[6\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13109__CLK clknet_leaf_21_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07212__I _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07345_ _02504_ _02820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10774__S _05237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07428__B2 u2.mem\[62\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07276_ u2.mem\[50\]\[3\] _02647_ _02648_ u2.mem\[51\]\[3\] _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_34_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09015_ _04135_ _04136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08228__I0 _03577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06227_ u2.mem\[193\]\[1\] _01731_ _01732_ u2.mem\[168\]\[1\] _01733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12133__CLK clknet_leaf_12_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10573__I _05094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13259__CLK clknet_leaf_311_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08043__I data_in_trans\[3\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06158_ _01564_ _01665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_137_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07087__C _02408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06403__A2 _01681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06089_ _01587_ _01596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09075__S _04182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12283__CLK clknet_leaf_188_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09917_ _04604_ _04709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11535__I0 _05715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08156__A2 _03583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09848_ _04576_ u2.mem\[40\]\[3\] _04661_ _04665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06167__A1 u2.mem\[144\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06706__A3 _02189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09779_ _04625_ _00615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11810_ _05768_ _05886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12790_ _00669_ clknet_leaf_33_clock u2.mem\[41\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11741_ _05833_ u2.mem\[183\]\[3\] _05840_ _05844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_2_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11672_ _05786_ u2.mem\[179\]\[0\] _05801_ _05802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07122__I _02600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13411_ _01290_ clknet_leaf_358_clock u2.mem\[172\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10623_ _05144_ _00940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_271_clock_I clknet_5_23_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10684__S _05179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13342_ _01221_ clknet_leaf_2_clock u2.mem\[160\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06961__I _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10554_ _05099_ u2.mem\[57\]\[2\] _05095_ _05100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08219__I0 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06642__A2 _02052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13273_ _01152_ clknet_leaf_7_clock u2.mem\[149\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10485_ _05007_ u2.mem\[55\]\[6\] _05056_ _05059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12224_ _00103_ clknet_leaf_241_clock u2.mem\[6\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11774__I0 _05837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12155_ _00034_ clknet_leaf_231_clock u2.mem\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08888__I _04050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_2_0_clock clknet_0_clock clknet_3_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_69_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_193_clock clknet_5_30_0_clock clknet_leaf_193_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_150_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11106_ _05420_ u2.mem\[144\]\[0\] _05445_ _05446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06945__A3 _02416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12086_ mem_write_n_trans.A clknet_leaf_317_clock mem_write_n_trans.data_sync vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11526__I0 _05707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11037_ _05401_ _01097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06201__I _01707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12006__CLK clknet_leaf_315_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11829__I1 u2.mem\[189\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12988_ _00867_ clknet_leaf_274_clock u2.mem\[54\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11939_ _05220_ u2.mem\[193\]\[11\] _05960_ _05964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_131_clock clknet_5_15_0_clock clknet_leaf_131_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08128__I _03545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06330__A1 u2.mem\[154\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07032__I _02373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06330__B2 u2.mem\[162\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12156__CLK clknet_leaf_219_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13401__CLK clknet_leaf_318_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07130_ _02573_ _02574_ _02401_ _02450_ _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_118_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08083__A1 _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_146_clock clknet_5_13_0_clock clknet_leaf_146_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10393__I _05000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07061_ u2.mem\[37\]\[0\] _02537_ _02539_ u2.mem\[59\]\[0\] _02540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_173_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07830__A1 u2.mem\[37\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06012_ _01516_ _01520_ _01521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08630__I0 _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06397__A1 u2.mem\[152\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07594__B1 _02905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07963_ u2.mem\[54\]\[15\] _02499_ _02501_ u2.mem\[55\]\[15\] _03427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_4_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11517__I0 _05674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06914_ _02390_ _02391_ _02392_ _02393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_09702_ _04126_ _04569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07894_ u2.mem\[9\]\[13\] _03304_ _03305_ u2.mem\[25\]\[13\] _03360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09623__S _04522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09633_ _04528_ _00566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06845_ u2.mem\[194\]\[5\] _02133_ _02134_ u2.mem\[190\]\[5\] _02325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10769__S _05232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11952__I _05971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09564_ _04486_ _00539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08239__S _03634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06776_ u2.mem\[165\]\[3\] _02075_ _02078_ u2.mem\[163\]\[3\] _02258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_5_4_0_clock clknet_4_2_0_clock clknet_5_4_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_110_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08515_ _03700_ _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09495_ _04442_ _04443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_19_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08446_ _03656_ u2.mem\[8\]\[0\] _03777_ _03778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_24_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06321__A1 u2.mem\[159\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06321__B2 u2.mem\[149\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06872__A2 _02350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08377_ _03684_ u2.mem\[6\]\[6\] _03732_ _03735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13081__CLK clknet_leaf_340_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07328_ _02469_ _02803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12649__CLK clknet_leaf_114_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11399__I _05507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07259_ u2.mem\[39\]\[2\] _02617_ _02619_ u2.mem\[48\]\[2\] _02736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06624__A2 _02037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10009__S _04762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10270_ _04893_ u2.mem\[50\]\[3\] _04923_ _04927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08702__S _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11756__I0 _05833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08621__I0 _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12799__CLK clknet_leaf_167_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06388__A1 u2.mem\[145\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06388__B2 u2.mem\[168\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06927__A3 _02392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_218_clock_I clknet_5_29_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12029__CLK clknet_2_2__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11133__A1 _05295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07117__I _02595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12911_ _00790_ clknet_leaf_162_clock u2.mem\[49\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10679__S _05174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12842_ _00721_ clknet_leaf_131_clock u2.mem\[44\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12773_ _00652_ clknet_leaf_76_clock u2.mem\[40\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13424__CLK clknet_leaf_361_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11724_ _03669_ _05833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06312__A1 u2.mem\[174\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06312__B2 u2.mem\[150\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11655_ _05667_ _05790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_63_clock clknet_5_9_0_clock clknet_leaf_63_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10247__I0 _04911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10606_ _05101_ u2.mem\[58\]\[3\] _05131_ _05135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11586_ _05662_ _05746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13574__CLK clknet_leaf_16_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07812__A1 u2.mem\[58\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10537_ _05020_ u2.mem\[56\]\[12\] _05088_ _05089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13325_ _01204_ clknet_leaf_323_clock u2.mem\[157\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06615__A2 _02060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08860__I0 _04037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07812__B2 u2.mem\[36\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_78_clock clknet_5_8_0_clock clknet_leaf_78_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_109_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09708__S _04567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08612__S _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10468_ _05027_ u2.mem\[54\]\[15\] _05045_ _05049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13256_ _01135_ clknet_leaf_287_clock u2.mem\[146\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12207_ _00086_ clknet_leaf_241_clock u2.mem\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10941__I _05339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08612__I0 _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13187_ _01066_ clknet_leaf_292_clock u2.mem\[134\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06379__A1 u2.mem\[180\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10399_ _05005_ u2.mem\[53\]\[5\] _05002_ _05006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06379__B2 u2.mem\[150\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12138_ _01464_ clknet_leaf_38_clock u2.driver_mem\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07040__A2 _02514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11973__S _05980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12080__D data_in_trans\[15\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12069_ net8 clknet_2_1__leaf_clock_a data_in_trans\[10\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07027__I _02347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07879__A1 u2.mem\[58\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07879__B2 u2.mem\[36\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06630_ _02114_ _02115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_16_clock clknet_5_2_0_clock clknet_leaf_16_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_20_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06561_ _02032_ _02036_ _02046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10388__I _04134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08300_ _03658_ _03676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_61_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09280_ _04285_ u2.mem\[26\]\[15\] _04305_ _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09340__I1 u2.mem\[28\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06303__A1 _01773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06492_ _01976_ _01970_ _01977_ _01978_ _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08231_ _03627_ _00065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10238__I0 _04904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08162_ _03550_ u2.mem\[2\]\[2\] _03585_ _03588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08056__A1 _01878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_167_clock_I clknet_5_26_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10789__I1 u2.mem\[62\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07113_ u2.mem\[17\]\[0\] _02586_ _02591_ u2.mem\[24\]\[0\] _02592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_146_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08093_ _03536_ _03537_ _00017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06606__A2 _01999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12941__CLK clknet_leaf_221_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11012__I _05342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07044_ _02448_ _02523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_118_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11363__A1 _03486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08321__I _03658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08995_ _04118_ _04119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11883__S _05932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07946_ u2.mem\[39\]\[14\] _03323_ _03324_ u2.mem\[48\]\[14\] _03411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_5_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06790__A1 _02245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input27_I mem_address_a[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10499__S _05066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07877_ u2.mem\[54\]\[13\] _02499_ _02501_ u2.mem\[55\]\[13\] _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_25_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_5_27_0_clock clknet_4_13_0_clock clknet_5_27_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_84_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12321__CLK clknet_leaf_167_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10713__I1 u2.mem\[61\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09616_ _04518_ _00559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06828_ u2.mem\[184\]\[5\] _02072_ _01994_ _02308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_44_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09547_ _04473_ u2.mem\[33\]\[4\] _04474_ _04475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06759_ u2.mem\[187\]\[3\] _02186_ _02187_ u2.mem\[192\]\[3\] _02241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_24_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12471__CLK clknet_leaf_127_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09478_ _04380_ u2.mem\[31\]\[10\] _04429_ _04432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08429_ _03766_ _00124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06845__A2 _02133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_156_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11440_ _04120_ _05645_ _05654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09095__I0 _04158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11371_ _05591_ u2.mem\[160\]\[3\] _05608_ _05612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10322_ _04956_ _00827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13110_ _00989_ clknet_leaf_20_clock u2.mem\[61\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07270__A2 _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13041_ _00920_ clknet_leaf_336_clock u2.mem\[57\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10253_ _04608_ _04916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07558__B1 _03028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10184_ _04871_ _00774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_369_clock_I clknet_5_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06781__A1 u2.mem\[150\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06781__B2 u2.mem\[174\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12814__CLK clknet_leaf_186_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12825_ _00704_ clknet_leaf_129_clock u2.mem\[43\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10468__I0 _05027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07089__A2 _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12756_ _00635_ clknet_leaf_71_clock u2.mem\[39\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11707_ _05794_ u2.mem\[181\]\[3\] _05818_ _05822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12687_ _00566_ clknet_leaf_157_clock u2.mem\[35\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08038__A1 _01727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09086__I0 _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11638_ _05746_ u2.mem\[177\]\[0\] _05779_ _05780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11569_ _05736_ _01294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13308_ _01187_ clknet_leaf_369_clock u2.mem\[154\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07261__A2 _02694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13239_ _01118_ clknet_leaf_303_clock u2.mem\[143\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09237__I _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08141__I _03545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07800_ _02466_ _03267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08780_ mem_address_trans\[5\].data_sync _03984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_111_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06772__A1 u2.mem\[184\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09173__S _04236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07731_ _03196_ _03197_ _03198_ _03199_ _03200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_37_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_93_clock_I clknet_5_10_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07662_ _02552_ _03132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12494__CLK clknet_leaf_197_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09401_ _04357_ _04385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_92_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06613_ _02006_ _02080_ _02098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_37_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07593_ u2.mem\[37\]\[8\] _03062_ _03063_ u2.mem\[59\]\[8\] _03064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_94_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09313__I1 u2.mem\[27\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09332_ _04340_ _00453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06544_ _02023_ _02028_ _02029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11120__I1 u2.mem\[145\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09263_ _04299_ _00425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06475_ _01962_ _01955_ _01963_ _01965_ _01459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_166_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08214_ _03607_ _03618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_21_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09077__I0 _04128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09194_ _04253_ _00402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11878__S _05929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08145_ _03575_ u2.mem\[1\]\[13\] _03573_ _03576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10631__I0 _05126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08076_ _01966_ _03516_ _03525_ _00012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_162_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07027_ _02347_ _02506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_122_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06460__B1 _01952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11187__I1 u2.mem\[149\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_370_clock_I clknet_5_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07555__A3 _03024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08978_ _04035_ u2.mem\[20\]\[9\] _04107_ _04109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_25_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06763__A1 u2.mem\[154\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06763__B2 u2.mem\[162\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12837__CLK clknet_leaf_88_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09001__I0 _04119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07929_ _03378_ _03383_ _03388_ _03393_ _03394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_60_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07307__A3 _02777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10022__S _04767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10940_ _04126_ _05339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07712__B1 _03126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06439__C _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10871_ _03582_ _05295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_45_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_1_0_clock clknet_3_0_0_clock clknet_4_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_38_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12987__CLK clknet_leaf_264_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09304__I1 u2.mem\[27\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12610_ _00489_ clknet_leaf_160_clock u2.mem\[30\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_61_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12541_ _00420_ clknet_leaf_198_clock u2.mem\[26\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12217__CLK clknet_leaf_44_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12472_ _00351_ clknet_leaf_123_clock u2.mem\[21\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11788__S _05866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11423_ _05635_ u2.mem\[163\]\[5\] _05637_ _05644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07779__B1 _03161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10622__I0 _05117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11354_ _05601_ _01214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08162__S _03585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07243__A2 _02666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10305_ _04891_ u2.mem\[51\]\[2\] _04944_ _04947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11285_ _05558_ _05559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_3_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10236_ _04591_ _04904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13024_ _00903_ clknet_leaf_265_clock u2.mem\[56\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10167_ _04817_ u2.mem\[47\]\[15\] _04856_ _04860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06754__A1 u2.mem\[169\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_115_clock_I clknet_5_14_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07951__B1 _03394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06754__B2 u2.mem\[147\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06410__S _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10098_ _04821_ _00738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11028__S _05395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_1_0_clock_I clknet_3_0_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09543__I1 u2.mem\[33\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07703__B1 _03034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12808_ _00687_ clknet_leaf_130_clock u2.mem\[42\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08337__S _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12739_ _00618_ clknet_leaf_29_clock u2.mem\[38\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06260_ u2.mem\[148\]\[1\] _01715_ _01698_ u2.mem\[154\]\[1\] u2.mem\[162\]\[1\]
+ _01700_ _01766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_54_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13142__CLK clknet_leaf_19_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06191_ _01567_ _01665_ _01678_ _01698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_156_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10613__I0 _05108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07234__A2 _02476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09950_ _04700_ u2.mem\[42\]\[8\] _04729_ _04730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13292__CLK clknet_leaf_382_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08901_ _04063_ _00299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09881_ _04684_ _00658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08832_ _04018_ _00275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06745__A1 u2.mem\[153\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06745__B2 u2.mem\[160\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08763_ _03925_ u2.mem\[15\]\[9\] _03972_ _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07714_ u2.mem\[43\]\[10\] _03053_ _03054_ u2.mem\[20\]\[10\] _03183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09534__I1 u2.mem\[33\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08694_ _03933_ _00222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07645_ u2.mem\[50\]\[9\] _03113_ _03114_ u2.mem\[51\]\[9\] _03115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07576_ _03039_ _03040_ _03043_ _03046_ _03047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_317_clock_I clknet_5_16_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09315_ _04281_ u2.mem\[27\]\[13\] _04328_ _04330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06527_ _02006_ _02011_ _02012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_167_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10576__I _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09246_ _04289_ _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_55_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06458_ u2.mem\[194\]\[7\] _01946_ _01952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07473__A2 _02943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09177_ _04225_ _04241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_147_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06389_ u2.mem\[187\]\[5\] _01633_ _01636_ u2.mem\[192\]\[5\] _01891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_147_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08017__A4 mem_address_trans\[7\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08128_ _03545_ _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10604__I0 _05099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07225__A2 _02638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08059_ _01945_ _03504_ _03513_ _00007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09806__S _04639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11070_ _05421_ _05422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09222__I0 _04272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08710__S _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10021_ _04770_ _00712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09773__I1 u2.mem\[38\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06736__B2 u2.mem\[161\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07933__B1 _02550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11580__I1 u2.mem\[173\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13015__CLK clknet_leaf_149_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09525__I1 u2.mem\[32\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11972_ _05983_ _01450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07125__I _02603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10923_ _05328_ _01056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06964__I _02394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10854_ _05284_ _01031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13165__CLK clknet_leaf_281_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13573_ _01452_ clknet_leaf_16_clock u2.mem\[194\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10785_ _05216_ u2.mem\[62\]\[9\] _05242_ _05244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11796__A1 _04310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12524_ _00403_ clknet_leaf_198_clock u2.mem\[25\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10843__I0 _05194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12455_ _00334_ clknet_leaf_135_clock u2.mem\[20\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_41_clock_I clknet_5_6_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11311__S _05567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11406_ _05633_ u2.mem\[162\]\[4\] _05624_ _05634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12386_ _00265_ clknet_leaf_158_clock u2.mem\[16\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11337_ _05590_ _01208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06975__A1 _02428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11268_ _05547_ _01182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13007_ _00886_ clknet_leaf_254_clock u2.mem\[55\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10219_ _04892_ _00788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11199_ _05500_ u2.mem\[150\]\[0\] _05502_ _05503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06727__A1 u2.mem\[150\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07924__B1 _02518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_266_clock_I clknet_5_22_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09516__I1 u2.mem\[32\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07035__I _02513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07430_ _02547_ _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_5_0_clock_I clknet_4_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07361_ _02563_ _02836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09100_ _04196_ _00365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06312_ u2.mem\[174\]\[3\] _01656_ _01666_ u2.mem\[150\]\[3\] _01660_ u2.mem\[181\]\[3\]
+ _01816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_52_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07292_ u2.mem\[26\]\[3\] _02675_ _02676_ u2.mem\[10\]\[3\] _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_149_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08652__A1 _03479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07455__A2 _02927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09031_ _04148_ u2.mem\[21\]\[6\] _04141_ _04149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06243_ _01621_ _01749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07207__A2 _02586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08404__A1 _03479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06174_ _01581_ _01600_ _01681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_171_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09933_ _04720_ _00674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09755__I1 u2.mem\[37\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09864_ _04599_ u2.mem\[40\]\[10\] _04671_ _04674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06718__A1 u2.mem\[176\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09425__I _04395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06718__B2 u2.mem\[172\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11562__I1 u2.mem\[172\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08815_ _04006_ _00270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09795_ _04634_ _00622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07391__A1 _01843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07391__B2 _02865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09507__I1 u2.mem\[32\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08746_ _03964_ _00243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12062__CLK clknet_leaf_374_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08677_ _03921_ _00217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08191__I0 _03579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07628_ _01954_ _03017_ _03057_ _03098_ _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_14_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07694__A2 _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06351__C1 u2.mem\[165\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07559_ _02456_ _03030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10570_ _05110_ u2.mem\[57\]\[7\] _05104_ _05111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09229_ _04277_ _00413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12240_ _00119_ clknet_leaf_240_clock u2.mem\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06406__B1 _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12171_ _00050_ clknet_leaf_233_clock u2.mem\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11122_ _05424_ u2.mem\[145\]\[1\] _05453_ _05455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_1_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11002__I0 _05352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11053_ _03902_ _05411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_67_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06709__A1 u2.mem\[180\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06709__B2 u2.mem\[150\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12405__CLK clknet_leaf_103_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10004_ _04440_ _04760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11553__I1 u2.mem\[171\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09271__S _04300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11305__I1 u2.mem\[156\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11955_ _05907_ u2.mem\[194\]\[1\] _05972_ _05974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12555__CLK clknet_leaf_206_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08182__I0 _03570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10906_ _04095_ _05317_ _05318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_44_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11886_ _05934_ _01413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10837_ mem_address_trans\[6\].data_sync _05273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11105__I _05444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13556_ _01435_ clknet_leaf_14_clock u2.mem\[193\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10768_ _05234_ _00995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12507_ _00386_ clknet_leaf_191_clock u2.mem\[24\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10944__I _04130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13487_ _01366_ clknet_leaf_314_clock u2.mem\[184\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11041__S _05404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10699_ _05119_ u2.mem\[60\]\[11\] _05184_ _05188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12438_ _00317_ clknet_leaf_102_clock u2.mem\[19\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08414__I _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11976__S _05985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10880__S _05297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12369_ _00248_ clknet_leaf_184_clock u2.mem\[15\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06948__A1 u2.mem\[27\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_361_clock clknet_5_4_0_clock clknet_leaf_361_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06930_ _02387_ _02389_ _02406_ _02408_ _02409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_113_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12085__CLK clknet_2_2__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input1_I col_select_a[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13330__CLK clknet_leaf_1_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06861_ row_select_trans\[0\].data_sync row_select_trans\[2\].data_sync _02340_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_45_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06176__A2 _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07373__B2 u2.mem\[24\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08600_ _03825_ u2.mem\[11\]\[12\] _03871_ _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09580_ _04497_ _00544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06792_ u2.mem\[151\]\[4\] _02084_ _02086_ u2.mem\[158\]\[4\] u2.mem\[168\]\[4\]
+ _02093_ _02273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_167_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_376_clock clknet_5_1_0_clock clknet_leaf_376_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08531_ _03721_ _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08173__I0 _03561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13480__CLK clknet_leaf_303_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08462_ _03786_ _00137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07676__A2 _03074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07413_ u2.mem\[58\]\[5\] _02811_ _02812_ u2.mem\[36\]\[5\] _02887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08393_ _03714_ u2.mem\[6\]\[13\] _03742_ _03744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11015__I _05345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07344_ u2.mem\[49\]\[4\] _02817_ _02818_ u2.mem\[46\]\[4\] _02819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07275_ _02746_ _02747_ _02748_ _02750_ _02751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_148_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09014_ _04134_ _04135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_314_clock clknet_5_17_0_clock clknet_leaf_314_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06226_ _01589_ _01732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08324__I data_in_trans\[9\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_0_0_clock clknet_4_0_0_clock clknet_5_0_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_163_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06157_ _01663_ _01664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12428__CLK clknet_leaf_192_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09356__S _04351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07061__B1 _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06088_ _01594_ _01595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_329_clock clknet_5_19_0_clock clknet_leaf_329_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_67_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09916_ _04708_ _00669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11535__I1 u2.mem\[170\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09847_ _04664_ _00644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12578__CLK clknet_leaf_185_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_9_clock_I clknet_5_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08994__I _04117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09778_ _04583_ u2.mem\[38\]\[5\] _04623_ _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08729_ _03954_ _00236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08164__I0 _03552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11126__S _05453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11740_ _05843_ _01358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10965__S _05356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11671_ _05800_ _05801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_53_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_214_clock_I clknet_5_29_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13410_ _01289_ clknet_leaf_323_clock u2.mem\[171\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10622_ _05117_ u2.mem\[58\]\[10\] _05141_ _05144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08435__S _03768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06627__B1 _02099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13341_ _01220_ clknet_leaf_1_clock u2.mem\[160\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10764__I _05231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10553_ _04994_ _05099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13203__CLK clknet_leaf_294_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13272_ _01151_ clknet_leaf_6_clock u2.mem\[148\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08234__I mem_address_trans\[2\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10484_ _05058_ _00887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12223_ _00102_ clknet_leaf_242_clock u2.mem\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11774__I1 u2.mem\[185\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12154_ _00033_ clknet_leaf_57_clock u2.mem\[1\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13353__CLK clknet_leaf_376_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11105_ _05444_ _05445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12085_ net34 clknet_2_2__leaf_clock_a mem_write_n_trans.A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11526__I1 u2.mem\[170\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11036_ _05392_ u2.mem\[139\]\[5\] _05394_ _05401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10004__I _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12987_ _00866_ clknet_leaf_264_clock u2.mem\[54\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11036__S _05394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07658__A2 _03050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11938_ _05963_ _01436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12078__D data_in_trans\[14\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11869_ _05913_ u2.mem\[191\]\[4\] _05917_ _05923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06330__A2 _01698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_158_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11462__I0 _05668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13539_ _01418_ clknet_leaf_11_clock u2.mem\[192\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10674__I _05173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08083__A2 _03528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07060_ _02538_ _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08144__I _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06011_ u2.driver_mem\[0\] _01512_ _01518_ _01519_ _01520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_173_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06397__A2 _01712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10115__S _04830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07962_ u2.mem\[50\]\[15\] _02493_ _02495_ u2.mem\[51\]\[15\] _03426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12720__CLK clknet_leaf_248_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_13_0_clock_I clknet_4_6_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11517__I1 u2.mem\[169\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09701_ _04568_ _00594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06913_ _02348_ _02350_ _02392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_101_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07893_ u2.mem\[29\]\[13\] _03301_ _03302_ u2.mem\[11\]\[13\] _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_25_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_163_clock_I clknet_5_26_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09632_ _04473_ u2.mem\[35\]\[4\] _04527_ _04528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06844_ u2.mem\[144\]\[5\] _02114_ _02116_ u2.mem\[182\]\[5\] _02324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07897__A2 _02594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09563_ _04485_ u2.mem\[33\]\[9\] _04483_ _04486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06775_ u2.mem\[151\]\[3\] _02084_ _02086_ u2.mem\[158\]\[3\] u2.mem\[193\]\[3\]
+ _02088_ _02257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_43_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08514_ _03820_ _00155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09494_ _03982_ _04441_ _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07649__A2 _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08319__I _03690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08445_ _03776_ _03777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_169_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12100__CLK clknet_leaf_246_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10785__S _05242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08376_ _03734_ _00103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07327_ u2.mem\[16\]\[4\] _02800_ _02801_ u2.mem\[33\]\[4\] _02802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_253_clock clknet_5_19_0_clock clknet_leaf_253_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_20_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07282__B1 _02660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12250__CLK clknet_leaf_56_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08054__I _03509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_23_0_clock clknet_4_11_0_clock clknet_5_23_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_07258_ u2.mem\[5\]\[2\] _02689_ _02690_ u2.mem\[38\]\[2\] _02735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__13376__CLK clknet_leaf_8_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_88_clock_I clknet_5_11_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06209_ u2.mem\[152\]\[0\] _01713_ _01715_ u2.mem\[148\]\[0\] _01716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07189_ _02554_ _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_156_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09086__S _04187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11756__I1 u2.mem\[184\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_268_clock clknet_5_22_0_clock clknet_leaf_268_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_155_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08621__I1 u2.mem\[12\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06388__A2 _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10025__S _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12910_ _00789_ clknet_leaf_202_clock u2.mem\[49\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10192__I0 _04801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12841_ _00720_ clknet_leaf_130_clock u2.mem\[44\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_206_clock clknet_5_31_0_clock clknet_leaf_206_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12772_ _00651_ clknet_leaf_64_clock u2.mem\[40\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07133__I _02611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11723_ _05832_ _01352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10695__S _05184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06312__A2 _01656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_365_clock_I clknet_5_4_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11654_ _05789_ _01326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11444__I0 _05627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10605_ _05134_ _00932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11585_ _05745_ _01301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06076__A1 _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13324_ _01203_ clknet_leaf_322_clock u2.mem\[157\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10536_ _05072_ _05088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_170_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13255_ _01134_ clknet_leaf_286_clock u2.mem\[146\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10467_ _05048_ _00880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12743__CLK clknet_leaf_43_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12206_ _00085_ clknet_leaf_227_clock u2.mem\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13186_ _01065_ clknet_leaf_293_clock u2.mem\[134\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06379__A2 _01664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10398_ _05004_ _05005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12137_ _01463_ clknet_leaf_38_clock u2.driver_mem\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12893__CLK clknet_leaf_224_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12068_ data_in_trans\[9\].A clknet_leaf_378_clock data_in_trans\[9\].data_sync vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11019_ _05390_ u2.mem\[138\]\[4\] _05381_ _05391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10183__I0 _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12123__CLK clknet_leaf_37_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13249__CLK clknet_leaf_302_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06551__A2 _01989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06560_ _02044_ _02045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07043__I _02446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06839__B1 _02099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10635__A1 _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06491_ u2.mem\[193\]\[14\] _01917_ _01919_ u2.mem\[192\]\[14\] _01920_ _01978_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_21_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07500__A1 _02957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08230_ _03579_ u2.mem\[3\]\[15\] _03623_ _03627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12273__CLK clknet_leaf_176_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06882__I _02360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13399__CLK clknet_leaf_314_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08161_ _03587_ _00035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07112_ _02590_ _02591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07264__B1 _02719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08092_ u2.driver_enable output_active_hold\[1\] output_active_hold\[0\] _03537_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_146_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07043_ _02446_ _02522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09800__I0 _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07567__A1 _03029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08994_ _04117_ _04118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06775__C1 u2.mem\[193\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07945_ u2.mem\[5\]\[14\] _02627_ _02629_ u2.mem\[38\]\[14\] _03410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_87_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06790__A2 _02249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07876_ u2.mem\[50\]\[13\] _02493_ _02495_ u2.mem\[51\]\[13\] _03342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10174__I0 _04782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09615_ _04494_ u2.mem\[34\]\[13\] _04516_ _04518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06827_ u2.mem\[167\]\[5\] _02059_ _02062_ u2.mem\[183\]\[5\] _02307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10579__I _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08119__I0 _03557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09546_ _04464_ _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08049__I _03505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06758_ u2.mem\[159\]\[3\] _02174_ _02176_ u2.mem\[149\]\[3\] _02240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12616__CLK clknet_leaf_136_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11674__I0 _05790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09477_ _04431_ _00507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06689_ u2.mem\[145\]\[1\] _02082_ _02094_ u2.mem\[168\]\[1\] _02173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08428_ _03701_ u2.mem\[7\]\[10\] _03763_ _03766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_192_clock clknet_5_30_0_clock clknet_leaf_192_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09619__I0 _04498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08359_ _03723_ _00097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12766__CLK clknet_leaf_219_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06058__A1 _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07255__B1 _02601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11370_ _05611_ _01220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10321_ _04907_ u2.mem\[51\]\[9\] _04954_ _04956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13040_ _00919_ clknet_leaf_336_clock u2.mem\[57\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08512__I _03696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10252_ _04915_ _00798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10183_ _04792_ u2.mem\[48\]\[4\] _04870_ _04871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_130_clock clknet_5_15_0_clock clknet_leaf_130_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_117_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08358__I0 _03722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06781__A2 _02047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_1_0_clock_I clknet_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06967__I _02386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10165__I0 _04815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11901__I1 _03522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10489__I _05050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12824_ _00703_ clknet_leaf_129_clock u2.mem\[43\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12296__CLK clknet_leaf_116_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13541__CLK clknet_leaf_18_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11665__I0 _05796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12755_ _00634_ clknet_leaf_68_clock u2.mem\[39\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06297__A1 u2.mem\[191\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11706_ _05821_ _01346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06297__B2 u2.mem\[179\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12686_ _00565_ clknet_leaf_216_clock u2.mem\[35\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11417__I0 _05629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11637_ _05778_ _05779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09086__I1 u2.mem\[22\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_111_clock_I clknet_5_11_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07246__B1 _02672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11568_ _05717_ u2.mem\[172\]\[4\] _05730_ _05736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_171_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13307_ _01186_ clknet_leaf_370_clock u2.mem\[154\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10952__I _04138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10519_ _05001_ u2.mem\[56\]\[4\] _05078_ _05079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11499_ _05668_ u2.mem\[168\]\[1\] _05692_ _05694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_48_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13238_ _01117_ clknet_leaf_302_clock u2.mem\[143\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08597__I0 _03823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11984__S _05971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12091__D net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13169_ _01048_ clknet_leaf_283_clock u2.mem\[131\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13071__CLK clknet_leaf_250_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07730_ u2.mem\[18\]\[10\] _03085_ _03086_ u2.mem\[19\]\[10\] _03199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_84_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10156__I0 _04806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12639__CLK clknet_leaf_159_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10856__A1 _05285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_36_clock_I clknet_5_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07661_ _03107_ _03112_ _03121_ _03130_ _03131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09400_ _04166_ _04384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06612_ _02096_ _02097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07592_ _02538_ _03063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09331_ _04258_ u2.mem\[28\]\[3\] _04336_ _04340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_146_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11656__I0 _05790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06543_ _02026_ _02027_ _02028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06288__A1 _01789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09262_ _04267_ u2.mem\[26\]\[7\] _04295_ _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07485__B1 _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06474_ u2.mem\[193\]\[10\] _01960_ _01948_ u2.mem\[192\]\[10\] _01964_ _01965_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_166_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08213_ _03617_ _00057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09193_ _04246_ u2.mem\[25\]\[0\] _04252_ _04253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09629__S _04522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12019__CLK clknet_2_3__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07237__B1 _02657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08144_ _03530_ _03575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08075_ _03524_ _03518_ _03525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10631__I1 u2.mem\[58\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07026_ _02504_ _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06460__A1 _01951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12169__CLK clknet_leaf_60_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08588__I0 _03814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11894__S _05937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_313_clock_I clknet_5_17_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10395__I0 _05001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06212__A1 _01613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08977_ _04108_ _00330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_62_clock clknet_5_9_0_clock clknet_leaf_62_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_102_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07928_ _03389_ _03390_ _03391_ _03392_ _03393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__10303__S _04944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10147__I0 _04797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13564__CLK clknet_leaf_10_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07859_ _02609_ _03326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07712__A1 u2.mem\[14\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10870_ _04986_ _05294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08708__S _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_77_clock clknet_5_8_0_clock clknet_leaf_77_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_25_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09529_ _04391_ u2.mem\[32\]\[15\] _04458_ _04462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12540_ _00419_ clknet_leaf_198_clock u2.mem\[26\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06455__C _01949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12471_ _00350_ clknet_leaf_127_clock u2.mem\[21\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10973__S _05355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07228__B1 _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11422_ _05643_ _01240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11024__A1 _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07779__A1 u2.mem\[6\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11353_ _05589_ u2.mem\[159\]\[2\] _05598_ _05601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10622__I1 u2.mem\[58\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_15_clock clknet_5_2_0_clock clknet_leaf_15_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_10_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10304_ _04946_ _00819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11284_ _04310_ _05527_ _05558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__08579__I0 _03805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13023_ _00902_ clknet_leaf_254_clock u2.mem\[56\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13094__CLK clknet_leaf_19_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10235_ _04903_ _00793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10386__I0 _04995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10166_ _04859_ _00768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07951__A1 _01976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06754__A2 _02141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11309__S _05567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10138__I0 _04788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10097_ _04782_ u2.mem\[46\]\[0\] _04820_ _04821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_59_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07703__A1 u2.mem\[16\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12931__CLK clknet_leaf_65_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08618__S _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_4_5_0_clock_I clknet_3_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12807_ _00686_ clknet_leaf_131_clock u2.mem\[42\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11638__I0 _05746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08503__I0 _03812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10999_ _05377_ _01083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12738_ _00617_ clknet_leaf_248_clock u2.mem\[38\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10310__I0 _04895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10883__S _05297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12669_ _00548_ clknet_leaf_217_clock u2.mem\[34\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_262_clock_I clknet_5_22_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06190_ u2.mem\[147\]\[0\] _01676_ _01680_ u2.mem\[169\]\[0\] _01696_ _01697_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_156_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11778__I _05865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12311__CLK clknet_leaf_115_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10613__I1 u2.mem\[58\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06442__A1 u2.mem\[194\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08900_ _04035_ u2.mem\[18\]\[9\] _04061_ _04063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09880_ _04681_ u2.mem\[41\]\[0\] _04683_ _04684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08195__A1 _03480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09184__S _04241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08831_ _04017_ u2.mem\[17\]\[1\] _04015_ _04018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12461__CLK clknet_leaf_194_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11219__S _05501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08762_ _03973_ _00250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07713_ u2.mem\[49\]\[10\] _03050_ _03051_ u2.mem\[46\]\[10\] _03182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09912__S _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08693_ _03931_ u2.mem\[13\]\[12\] _03932_ _03933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11018__I _05348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07644_ _02494_ _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10857__I _05286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07575_ u2.mem\[58\]\[8\] _03044_ _03045_ u2.mem\[36\]\[8\] _03046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_53_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09314_ _04329_ _00446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07458__B1 _02898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06526_ _02010_ _02000_ _02011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10301__I0 _04885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11889__S _05932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09245_ _04288_ _04250_ _04289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06457_ u2.mem\[0\]\[7\] _01951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_72_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07473__A3 _02944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06681__A1 u2.mem\[144\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09176_ _04240_ _00397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08263__S _03644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06681__B2 u2.mem\[182\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06388_ u2.mem\[145\]\[5\] _01640_ _01732_ u2.mem\[168\]\[5\] _01890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10592__I _03716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08127_ _03517_ _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10604__I1 u2.mem\[58\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06433__A1 u2.mem\[192\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08058_ _03512_ _03507_ _03513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07009_ _02441_ _02381_ _02382_ _02488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA__09222__I1 u2.mem\[25\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10368__I0 _04916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08997__I _04120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10020_ _04696_ u2.mem\[44\]\[6\] _04767_ _04770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07528__A4 _02999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06736__A2 _02097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07933__A1 u2.mem\[57\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12954__CLK clknet_leaf_146_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08011__B _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07406__I _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09822__S _04649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11971_ _05213_ u2.mem\[194\]\[8\] _05980_ _05983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10922_ _05294_ u2.mem\[133\]\[0\] _05327_ _05328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07697__B1 _03020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10853_ _05207_ u2.mem\[128\]\[5\] _05277_ _05284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13572_ _01451_ clknet_leaf_15_clock u2.mem\[194\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10784_ _05243_ _01002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12523_ _00402_ clknet_leaf_187_clock u2.mem\[25\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11796__A2 _05847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12334__CLK clknet_leaf_234_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09269__S _04300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06672__A1 _02125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12454_ _00333_ clknet_leaf_89_clock u2.mem\[20\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06980__I _02394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11405_ _05513_ _05633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12385_ _00264_ clknet_leaf_235_clock u2.mem\[16\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09068__I _04176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06424__A1 u2.mem\[194\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12484__CLK clknet_leaf_107_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07621__B1 _03091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11336_ _05589_ u2.mem\[158\]\[2\] _05585_ _05590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06975__A2 _02390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10359__I0 _04907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11267_ _05544_ u2.mem\[154\]\[0\] _05546_ _05547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13006_ _00885_ clknet_leaf_270_clock u2.mem\[55\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10218_ _04891_ u2.mem\[49\]\[2\] _04887_ _04892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11198_ _05501_ _05502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_67_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_209_clock_I clknet_5_28_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06727__A2 _02192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10149_ _04799_ u2.mem\[47\]\[7\] _04846_ _04850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08724__I0 _03922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07688__B1 _03091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09531__I _04118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07152__A2 _02620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11236__A1 _04223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07360_ _02558_ _02835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08147__I _03532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08101__A1 _03482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06311_ u2.mem\[155\]\[3\] _01659_ _01815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07291_ _02763_ _02764_ _02765_ _02766_ _02767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__08652__A2 _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09030_ _04147_ _04148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_5_9_0_clock_I clknet_4_4_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06890__I _02368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06242_ u2.mem\[178\]\[1\] _01746_ _01747_ u2.mem\[164\]\[1\] _01748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12827__CLK clknet_leaf_184_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06173_ _01679_ _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08404__A2 _03751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08811__S _04000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09932_ _04681_ u2.mem\[42\]\[0\] _04719_ _04720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12977__CLK clknet_leaf_253_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09706__I _04130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09863_ _04673_ _00651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08814_ _03931_ u2.mem\[16\]\[12\] _04005_ _04006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07915__B2 u2.mem\[7\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09794_ _04605_ u2.mem\[38\]\[12\] _04633_ _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12207__CLK clknet_leaf_241_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06130__I _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08745_ _03907_ u2.mem\[15\]\[1\] _03962_ _03964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08715__I0 _03913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08676_ _03920_ u2.mem\[13\]\[7\] _03914_ _03921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_26_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07627_ _03066_ _03077_ _03088_ _03097_ _03098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_42_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12357__CLK clknet_leaf_95_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06351__B1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07694__A3 _03154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07558_ u2.mem\[15\]\[8\] _03027_ _03028_ u2.mem\[13\]\[8\] _03029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08057__I data_in_trans\[6\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06509_ _01993_ _01994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07489_ _02958_ _02959_ _02960_ _02961_ _02962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__09840__A1 _04224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09228_ _04276_ u2.mem\[25\]\[11\] _04270_ _04277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_5_clock_I clknet_5_0_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_158_clock_I clknet_5_25_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09159_ _04225_ _04231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_159_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06406__A1 u2.mem\[147\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12170_ _00049_ clknet_leaf_59_clock u2.mem\[2\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06305__I _01808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11121_ _05454_ _01128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11950__A2 _05926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11052_ _05410_ _01103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_210_clock_I clknet_5_28_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06709__A2 _02043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10003_ _04759_ _00705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10761__I0 _05229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09659__A1 _04095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08706__I0 _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_18_0_clock clknet_4_9_0_clock clknet_5_18_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_3742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11954_ _05973_ _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09351__I _04335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07134__A2 _02610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10905_ _05275_ _05317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_166_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06342__B1 _01663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11885_ u2.mem\[192\]\[3\] _03502_ _05932_ _05934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13282__CLK clknet_leaf_383_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06342__C2 u2.mem\[176\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06893__A1 _02364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10836_ _05272_ _01025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13555_ _01434_ clknet_leaf_15_clock u2.mem\[193\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10767_ _05198_ u2.mem\[62\]\[1\] _05232_ _05234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12506_ _00385_ clknet_leaf_126_clock u2.mem\[23\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13486_ _01365_ clknet_leaf_306_clock u2.mem\[184\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10698_ _05187_ _00972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12437_ _00316_ clknet_leaf_102_clock u2.mem\[19\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06215__I _01721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12368_ _00247_ clknet_leaf_183_clock u2.mem\[15\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06948__A2 _02420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07070__A1 _02395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11319_ _05550_ u2.mem\[157\]\[2\] _05576_ _05579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12299_ _00178_ clknet_leaf_206_clock u2.mem\[11\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06860_ _02025_ _01989_ _02339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10752__I0 _05222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09462__S _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06791_ _01809_ _01995_ _02244_ _02272_ _01477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_48_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08530_ _03831_ _00160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08173__I1 u2.mem\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08461_ _03688_ u2.mem\[8\]\[7\] _03782_ _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07412_ u2.mem\[53\]\[5\] _02808_ _02809_ u2.mem\[56\]\[5\] _02886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_168_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10200__I _04864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08392_ _03743_ _00110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07343_ _02531_ _02818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07833__B1 _03142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07274_ u2.mem\[3\]\[3\] _02470_ _02749_ _02750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09013_ data_in_trans\[3\].data_sync _04134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06225_ _01577_ _01731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06156_ _01623_ _01618_ _01663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06125__I _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11966__I _05971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10870__I _04986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06087_ _01556_ _01569_ _01593_ _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_160_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13155__CLK clknet_leaf_281_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08340__I _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09915_ _04707_ u2.mem\[41\]\[11\] _04701_ _04708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09846_ _04573_ u2.mem\[40\]\[2\] _04661_ _04664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_63_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08010__B1 _03459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09372__S _04358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09777_ _04624_ _00614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06989_ u2.mem\[16\]\[0\] _02465_ _02467_ u2.mem\[33\]\[0\] _02468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08728_ _03927_ u2.mem\[14\]\[10\] _03951_ _03954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_84_clock_I clknet_5_9_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08659_ _03666_ _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11206__I _05507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06875__A1 row_select_trans\[1\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11670_ _04071_ _05769_ _05800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_53_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10621_ _05143_ _00939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13340_ _01219_ clknet_leaf_2_clock u2.mem\[160\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08515__I _03700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06627__B2 u2.mem\[161\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10552_ _05098_ _00915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07824__B1 _03133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08092__A3 output_active_hold\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13271_ _01150_ clknet_leaf_4_clock u2.mem\[148\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10483_ _05005_ u2.mem\[55\]\[5\] _05056_ _05058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09547__S _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12222_ _00101_ clknet_leaf_225_clock u2.mem\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11223__I1 u2.mem\[151\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06035__I _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11876__I _05927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07052__A1 _02395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12153_ _00032_ clknet_leaf_56_clock u2.mem\[1\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10982__I0 _05343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06260__C1 u2.mem\[162\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11104_ _03486_ _05443_ _05444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_12084_ net48 clknet_leaf_381_clock output_active_hold\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_361_clock_I clknet_5_4_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12522__CLK clknet_leaf_124_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11035_ _05400_ _01096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06563__B1 _02047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11317__S _05576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10221__S _04887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12986_ _00865_ clknet_leaf_50_clock u2.mem\[53\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09352__I0 _04278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11937_ _05218_ u2.mem\[193\]\[10\] _05960_ _05963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06866__A1 _02339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11868_ _05922_ _01407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09104__I0 _04171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10819_ _05252_ _05263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_105_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11799_ _05880_ _01380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06618__A1 _02014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07815__B1 _03126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11462__I1 u2.mem\[166\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13538_ _01417_ clknet_leaf_34_clock u2.mem\[192\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06094__A2 _01587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12094__D _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13469_ _01348_ clknet_leaf_360_clock u2.mem\[181\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_174_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06010_ _01503_ _01519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13178__CLK clknet_leaf_293_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10973__I0 _05352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07594__A2 _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07961_ _03421_ _03422_ _03423_ _03424_ _03425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_59_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09700_ _04565_ u2.mem\[37\]\[0\] _04567_ _04568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06912_ _02380_ _02391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_136_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07892_ u2.mem\[26\]\[13\] _02567_ _02569_ u2.mem\[10\]\[13\] _03358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_136_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06149__A3 _01596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_106_clock_I clknet_5_11_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09631_ _04521_ _04527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_28_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06843_ _02319_ _02320_ _02321_ _02322_ _02323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_55_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11227__S _05520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_17_0_clock_I clknet_4_8_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09562_ _04157_ _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06774_ u2.mem\[168\]\[3\] _02093_ _02256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09343__I0 _04269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08513_ _03819_ u2.mem\[9\]\[9\] _03817_ _03820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09493_ _04440_ _04441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11150__I0 _05472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06857__A1 _02309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08444_ _03629_ _03541_ _03775_ _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__08536__S _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08375_ _03680_ u2.mem\[6\]\[5\] _03732_ _03734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07326_ _02466_ _02801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07806__B1 _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08335__I _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07282__A1 u2.mem\[14\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06085__A2 _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07257_ _02730_ _02731_ _02732_ _02733_ _02734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_20_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07282__B2 u2.mem\[12\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06208_ _01714_ _01715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07188_ _02552_ _02666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_151_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07034__A1 _02455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12545__CLK clknet_leaf_178_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06139_ _01645_ _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06793__B1 _02088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08909__I0 _04044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10105__I _04819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10716__I0 _05198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12695__CLK clknet_leaf_140_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09582__I0 _04498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09829_ _04653_ _00637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10192__I1 u2.mem\[48\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12840_ _00719_ clknet_leaf_130_clock u2.mem\[44\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09334__I0 _04260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12771_ _00650_ clknet_leaf_83_clock u2.mem\[40\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11141__I0 _05466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11722_ _05831_ u2.mem\[182\]\[2\] _05827_ _05832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08446__S _03777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_308_clock_I clknet_5_20_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11653_ _05786_ u2.mem\[178\]\[0\] _05788_ _05789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_360_clock clknet_5_5_0_clock clknet_leaf_360_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_122_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12075__CLK clknet_2_0__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10604_ _05099_ u2.mem\[58\]\[2\] _05131_ _05134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_174_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11444__I1 u2.mem\[165\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11584_ _05719_ u2.mem\[173\]\[5\] _05738_ _05745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13320__CLK clknet_leaf_323_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13323_ _01202_ clknet_leaf_322_clock u2.mem\[157\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10535_ _05087_ _00909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06076__A2 _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13254_ _01133_ clknet_leaf_308_clock u2.mem\[145\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10466_ _05025_ u2.mem\[54\]\[14\] _05045_ _05048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_375_clock clknet_5_1_0_clock clknet_leaf_375_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_108_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07025__A1 _02421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12205_ _00084_ clknet_leaf_267_clock u2.mem\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13185_ _01064_ clknet_leaf_294_clock u2.mem\[134\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13470__CLK clknet_leaf_360_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10397_ _04143_ _05004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07576__A2 _03040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12136_ _01462_ clknet_leaf_38_clock u2.driver_mem\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06784__B1 _02148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10015__I _04761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12067_ net22 clknet_2_1__leaf_clock_a data_in_trans\[9\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09573__I0 _04491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11018_ _05348_ _05390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11047__S _05404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06536__C2 u2.mem\[189\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06000__A2 _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_313_clock clknet_5_17_0_clock clknet_leaf_313_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09325__I0 _04246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12089__D net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10886__S _05296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12969_ _00848_ clknet_leaf_127_clock u2.mem\[52\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06839__A1 u2.mem\[166\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06839__B2 u2.mem\[161\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06490_ u2.mem\[194\]\[14\] _01933_ _01977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12418__CLK clknet_leaf_171_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07500__A2 _02962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_328_clock clknet_5_17_0_clock clknet_leaf_328_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_159_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08160_ _03548_ u2.mem\[2\]\[1\] _03585_ _03587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07111_ _02587_ _02588_ _02401_ _02589_ _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_14_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07264__A1 _01772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12568__CLK clknet_leaf_135_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07264__B2 _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08091_ output_active_hold\[3\] output_active_hold\[2\] _03536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_32_clock_I clknet_5_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07042_ _02520_ _02521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10126__S _04835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10946__I0 _05343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09915__S _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08993_ data_in_trans\[0\].data_sync _04117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06775__B1 _02086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06775__C2 _02088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07944_ _03405_ _03406_ _03407_ _03408_ _03409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_116_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09714__I _04138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_257_clock_I clknet_5_19_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06790__A3 _02250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07875_ _03337_ _03338_ _03339_ _03340_ _03341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_21_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11371__I0 _05591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09614_ _04517_ _00558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06826_ u2.mem\[164\]\[5\] _02051_ _02054_ u2.mem\[178\]\[5\] _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09545_ _04139_ _04473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06757_ _01773_ _01996_ _02239_ _01476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10796__S _05247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12098__CLK clknet_leaf_246_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09476_ _04378_ u2.mem\[31\]\[9\] _04429_ _04431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11674__I1 u2.mem\[179\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06688_ u2.mem\[151\]\[1\] _02085_ _02087_ u2.mem\[158\]\[1\] u2.mem\[193\]\[1\]
+ _02089_ _02172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_145_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13343__CLK clknet_leaf_2_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08427_ _03765_ _00123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10595__I _03720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08358_ _03722_ u2.mem\[5\]\[15\] _03710_ _03723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08065__I _03492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07255__A1 u2.mem\[52\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07309_ _02360_ _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08289_ _03666_ _03667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13493__CLK clknet_leaf_309_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09097__S _04192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10320_ _04955_ _00826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10251_ _04913_ u2.mem\[49\]\[12\] _04914_ _04915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10036__S _04777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07558__A2 _03027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07409__I _02498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10182_ _04864_ _04870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_59_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07191__B1 _02544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09560__S _04483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12823_ _00702_ clknet_leaf_129_clock u2.mem\[43\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_3_5_0_clock_I clknet_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08176__S _03595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12754_ _00633_ clknet_leaf_247_clock u2.mem\[39\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11665__I1 u2.mem\[178\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11705_ _05792_ u2.mem\[181\]\[2\] _05818_ _05821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12685_ _00564_ clknet_leaf_217_clock u2.mem\[35\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12710__CLK clknet_leaf_65_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11636_ _05285_ _05769_ _05778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__11417__I1 u2.mem\[163\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08904__S _04061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11567_ _05735_ _01293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11330__S _05585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13306_ _01185_ clknet_leaf_376_clock u2.mem\[154\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10518_ _05072_ _05078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_156_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11498_ _05693_ _01266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12860__CLK clknet_leaf_215_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13237_ _01116_ clknet_leaf_302_clock u2.mem\[143\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10449_ _05038_ _00872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_152_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10928__I0 _05303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07319__I _02444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09794__I0 _04605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06223__I _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13168_ _01047_ clknet_leaf_279_clock u2.mem\[131\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07013__A4 _02393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13216__CLK clknet_leaf_297_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12119_ _01482_ clknet_leaf_343_clock u2.select_mem_col\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13099_ _00978_ clknet_leaf_260_clock u2.mem\[61\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_252_clock clknet_5_19_0_clock clknet_leaf_252_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11353__I0 _05589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07660_ _03124_ _03127_ _03128_ _03129_ _03130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_37_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06611_ _02006_ _02046_ _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_168_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07591_ _02536_ _03062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09330_ _04339_ _00452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11505__S _05691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06542_ _01988_ _02009_ _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_267_clock clknet_5_22_0_clock clknet_leaf_267_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11656__I1 u2.mem\[178\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09261_ _04298_ _00424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06473_ _01913_ _01964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08212_ _03561_ u2.mem\[3\]\[7\] _03613_ _03617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09192_ _04251_ _04252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_159_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08143_ _03574_ _00030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08285__I0 _03663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11240__S _05529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08074_ data_in_trans\[11\].data_sync _03524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07252__A4 _02728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07025_ _02421_ _02433_ _02434_ _02417_ _02504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__06460__A2 _01938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_205_clock clknet_5_31_0_clock clknet_leaf_205_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_162_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_161_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09645__S _04532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09785__I0 _04592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06133__I _01639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11592__I0 _05750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06212__A2 _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08976_ _04032_ u2.mem\[20\]\[8\] _04107_ _04108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_25_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input32_I mem_address_a[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09537__I0 _04467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07927_ u2.mem\[43\]\[14\] _03286_ _03287_ u2.mem\[20\]\[14\] _03392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_152_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07858_ u2.mem\[39\]\[12\] _03323_ _03324_ u2.mem\[48\]\[12\] _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_29_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07712__A2 _03125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06809_ _02286_ _02287_ _02288_ _02289_ _02290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_56_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07789_ _02409_ _03256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12733__CLK clknet_leaf_271_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11415__S _05638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09528_ _04461_ _00528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_149_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09459_ _04421_ _00499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06279__A2 _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11214__I _05513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12470_ _00349_ clknet_leaf_103_clock u2.mem\[21\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08724__S _03951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11421_ _05633_ u2.mem\[163\]\[4\] _05637_ _05643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07228__B2 u2.mem\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11150__S _05461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07779__A2 _03160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11352_ _05600_ _01213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10303_ _04889_ u2.mem\[51\]\[1\] _04944_ _04946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_12_0_clock_I clknet_3_6_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13239__CLK clknet_leaf_303_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11283_ _05557_ _01187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09776__I0 _04579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13022_ _00901_ clknet_leaf_272_clock u2.mem\[56\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10234_ _04902_ u2.mem\[49\]\[7\] _04896_ _04903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06043__I col_select_trans\[5\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06739__B1 _02089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07400__A1 _02868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06978__I _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10165_ _04815_ u2.mem\[47\]\[14\] _04856_ _04859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_171_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12263__CLK clknet_leaf_54_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13389__CLK clknet_leaf_372_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10096_ _04819_ _04820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_134_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10838__A2 mem_address_trans\[7\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07164__B1 _02452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09290__S _04313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07703__A2 _03033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11325__S _05575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12806_ _00685_ clknet_leaf_87_clock u2.mem\[42\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11638__I1 u2.mem\[177\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10998_ _05346_ u2.mem\[137\]\[3\] _05373_ _05377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_167_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09700__I0 _04565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12737_ _00616_ clknet_leaf_247_clock u2.mem\[38\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_205_clock_I clknet_5_31_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_9_0_clock_I clknet_3_4_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08634__S _03889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12668_ _00547_ clknet_leaf_217_clock u2.mem\[34\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11619_ _05767_ _01313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12599_ _00478_ clknet_leaf_115_clock u2.mem\[29\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11060__S _05413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10074__I0 _04804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06442__A2 _01924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07049__I _02527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09767__I0 _04565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12606__CLK clknet_leaf_202_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11574__I0 _05707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08830_ _03662_ _04017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06888__I _02353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_191_clock clknet_5_30_0_clock clknet_leaf_191_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09264__I _04289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08761_ _03922_ u2.mem\[15\]\[8\] _03972_ _03973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07712_ u2.mem\[14\]\[10\] _03125_ _03126_ u2.mem\[12\]\[10\] _03181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12756__CLK clknet_leaf_71_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08692_ _03904_ _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_122_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08809__S _04000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07643_ _02492_ _03113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07574_ _02489_ _03045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09313_ _04278_ u2.mem\[27\]\[12\] _04328_ _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07458__A1 _01877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06525_ _02008_ _02009_ _02010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_40_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07458__B2 _02931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10301__I1 u2.mem\[51\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09244_ _04287_ _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_167_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06456_ _01945_ _01938_ _01947_ _01950_ _01470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12136__CLK clknet_leaf_38_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09175_ _04164_ u2.mem\[24\]\[11\] _04236_ _04240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10873__I _05296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06387_ u2.mem\[158\]\[5\] _01728_ _01729_ u2.mem\[151\]\[5\] _01577_ u2.mem\[193\]\[5\]
+ _01889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_08126_ _03562_ _00025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_144_clock clknet_5_13_0_clock clknet_leaf_144_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06433__A2 _01931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08057_ data_in_trans\[6\].data_sync _03512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07008_ _02486_ _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13531__CLK clknet_leaf_348_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10314__S _04949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08430__I0 _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_159_clock clknet_5_27_0_clock clknet_leaf_159_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_27_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06197__A1 _01552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07394__B1 _02867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07933__A2 _02548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08959_ _04098_ _00322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11317__I0 _05548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_1_clock_I clknet_5_0_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11209__I _03501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_154_clock_I clknet_5_24_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11970_ _05982_ _01449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07146__B1 _02624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07697__A1 u2.mem\[32\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10921_ _05326_ _05327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_3968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10852_ _05283_ _01030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08518__I _03704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08497__I0 _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10984__S _05365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13571_ _01450_ clknet_leaf_15_clock u2.mem\[194\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10783_ _05213_ u2.mem\[62\]\[8\] _05242_ _05243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12522_ _00401_ clknet_leaf_124_clock u2.mem\[24\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06038__I _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12453_ _00332_ clknet_leaf_90_clock u2.mem\[20\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06672__A2 _02014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13061__CLK clknet_leaf_29_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_14_0_clock clknet_4_7_0_clock clknet_5_14_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_11404_ _05632_ _01233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12384_ _00263_ clknet_leaf_234_clock u2.mem\[16\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_79_clock_I clknet_5_8_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11335_ _05507_ _05589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06424__A2 _01924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07621__B2 u2.mem\[48\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06975__A3 _02381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11266_ _05545_ _05546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_10_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10508__A1 _04224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10217_ _04572_ _04891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12779__CLK clknet_leaf_265_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13005_ _00884_ clknet_leaf_273_clock u2.mem\[55\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08421__I0 _03688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11197_ _04179_ _05482_ _05501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__06188__A1 u2.mem\[146\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11181__A1 _04120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07924__A2 _02514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10148_ _04849_ _00760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06501__I row_select_trans\[1\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11119__I _05452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10079_ _04601_ _04808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12009__CLK clknet_2_1__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09812__I _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08724__I1 u2.mem\[14\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07688__B2 u2.mem\[48\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06360__B2 u2.mem\[194\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12159__CLK clknet_leaf_236_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12097__D _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10295__I0 _04918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06310_ _01810_ _01811_ _01812_ _01813_ _01814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08101__A2 _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08364__S _03727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07290_ u2.mem\[57\]\[3\] _02671_ _02672_ u2.mem\[41\]\[3\] _02766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06112__A1 _01618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06241_ _01619_ _01747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_61_clock clknet_5_9_0_clock clknet_leaf_61_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_129_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06172_ _01678_ _01644_ _01588_ _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__13554__CLK clknet_leaf_10_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08660__I0 _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09931_ _04718_ _04719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_132_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_76_clock clknet_5_8_0_clock clknet_leaf_76_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11547__I0 _05711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08412__I0 _03671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09862_ _04596_ u2.mem\[40\]\[9\] _04671_ _04673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10134__S _04841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06179__A1 _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08813_ _03989_ _04005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09793_ _04617_ _04633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08744_ _03963_ _00242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07128__B1 _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09912__I0 _04705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08675_ _03687_ _03920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07626_ _03089_ _03092_ _03095_ _03096_ _03097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_42_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_14_clock clknet_5_2_0_clock clknet_leaf_14_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06351__A1 u2.mem\[145\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06351__B2 u2.mem\[163\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07557_ _02451_ _03028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08479__I0 _03722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13084__CLK clknet_leaf_277_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10286__I0 _04909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06508_ _01987_ _01991_ _01992_ _01993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_139_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07488_ u2.mem\[28\]\[6\] _02841_ _02842_ u2.mem\[31\]\[6\] _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_21_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06103__A1 _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07300__B1 _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09840__A2 _04659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_29_clock clknet_5_3_0_clock clknet_leaf_29_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09227_ _04163_ _04276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06654__A2 _02135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06439_ u2.mem\[193\]\[3\] _01928_ _01933_ u2.mem\[194\]\[3\] _01934_ _01937_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_167_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10038__I0 _04714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09158_ _04230_ _00389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_80_clock_I clknet_5_8_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08109_ _03550_ u2.mem\[1\]\[2\] _03546_ _03551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06406__A2 _01675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09089_ _04190_ _00360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11120_ _05420_ u2.mem\[145\]\[0\] _05453_ _05454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_162_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11538__I0 _05717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11051_ _05392_ u2.mem\[140\]\[5\] _05403_ _05410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10002_ _04716_ u2.mem\[43\]\[15\] _04755_ _04759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09833__S _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09659__A2 _04542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06590__A1 _02031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11953_ _05903_ u2.mem\[194\]\[0\] _05972_ _05973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12301__CLK clknet_leaf_205_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13427__CLK clknet_leaf_365_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10904_ _05316_ _01049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06342__A1 u2.mem\[189\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11884_ _05933_ _01412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06342__B2 u2.mem\[180\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10835_ u2.mem\[63\]\[15\] _05229_ _05268_ _05272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10277__I0 _04900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06991__I _02469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13554_ _01433_ clknet_leaf_10_clock u2.mem\[193\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12451__CLK clknet_leaf_112_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10766_ _05233_ _00994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13577__CLK clknet_leaf_35_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12505_ _00384_ clknet_leaf_126_clock u2.mem\[23\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06645__A2 _02070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13485_ _01364_ clknet_leaf_305_clock u2.mem\[184\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10697_ _05117_ u2.mem\[60\]\[10\] _05184_ _05187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11402__I _05510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10029__I0 _04705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12436_ _00315_ clknet_leaf_102_clock u2.mem\[19\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_2_2__f_clock_a clknet_0_clock_a clknet_2_2__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_153_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12367_ _00246_ clknet_leaf_183_clock u2.mem\[15\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06940__B _02417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11318_ _05578_ _01201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12298_ _00177_ clknet_leaf_122_clock u2.mem\[10\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11529__I0 _05711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11249_ _05535_ _01175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10201__I0 _04810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10889__S _05296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06790_ _02245_ _02249_ _02250_ _02271_ _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_83_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09542__I _04135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11701__I0 _05786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08460_ _03785_ _00136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06333__A1 u2.mem\[191\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06333__B2 u2.mem\[179\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07411_ u2.mem\[54\]\[5\] _02883_ _02884_ u2.mem\[55\]\[5\] _02885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08391_ _03709_ u2.mem\[6\]\[12\] _03742_ _03743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10268__I0 _04891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11513__S _05700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07342_ _02527_ _02817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08086__A1 _03532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07833__A1 u2.mem\[26\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07273_ _02358_ _02749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_102_clock_I clknet_5_10_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09012_ _04133_ _00340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12944__CLK clknet_leaf_151_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06224_ u2.mem\[163\]\[1\] _01643_ _01646_ u2.mem\[165\]\[1\] _01730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_157_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11768__I0 _05831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06155_ u2.mem\[174\]\[0\] _01657_ _01659_ u2.mem\[155\]\[0\] _01661_ u2.mem\[181\]\[0\]
+ _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_89_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06086_ _01573_ _01575_ _01593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__07061__A2 _02537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09914_ _04601_ _04707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09845_ _04663_ _00643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12324__CLK clknet_leaf_95_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09776_ _04579_ u2.mem\[38\]\[4\] _04623_ _04624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06988_ _02466_ _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08727_ _03953_ _00235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08068__I data_in_trans\[9\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08658_ _03908_ _00211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12474__CLK clknet_leaf_127_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07609_ _02590_ _03080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08589_ _03865_ _00185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11423__S _05637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10620_ _05115_ u2.mem\[58\]\[9\] _05141_ _05143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06627__A2 _02097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10551_ _05097_ u2.mem\[57\]\[1\] _05095_ _05098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11222__I _05519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09828__S _04649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13270_ _01149_ clknet_leaf_5_clock u2.mem\[148\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10482_ _05057_ _00886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12221_ _00100_ clknet_leaf_226_clock u2.mem\[6\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12152_ _00031_ clknet_leaf_65_clock u2.mem\[1\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10431__I0 _05027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08531__I _03721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11103_ _05442_ _05443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06260__B1 _01698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12083_ net47 clknet_leaf_381_clock output_active_hold\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_304_clock_I clknet_5_20_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06260__C2 _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09563__S _04483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11034_ _05390_ u2.mem\[139\]\[4\] _05394_ _05400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06051__I col_select_trans\[2\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06986__I _02464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06563__A1 u2.mem\[180\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09362__I _04357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06563__B2 u2.mem\[150\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12817__CLK clknet_leaf_167_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12985_ _00864_ clknet_leaf_50_clock u2.mem\[53\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11936_ _05962_ _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08907__S _04066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06866__A2 _02344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11867_ _05911_ u2.mem\[191\]\[3\] _05918_ _05922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12967__CLK clknet_leaf_128_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11333__S _05585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10818_ _05262_ _01017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11798_ _05864_ u2.mem\[187\]\[0\] _05879_ _05880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06618__A2 _02011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13537_ _01416_ clknet_leaf_34_clock u2.mem\[192\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08863__I0 _04039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10749_ _05221_ _00989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11132__I _05334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09738__S _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10670__I0 _05128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06226__I _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13468_ _01347_ clknet_leaf_360_clock u2.mem\[181\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07291__A2 _02764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12419_ _00298_ clknet_leaf_104_clock u2.mem\[18\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13399_ _01278_ clknet_leaf_314_clock u2.mem\[170\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10422__I0 _05020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08441__I mem_address_trans\[3\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12347__CLK clknet_leaf_209_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07960_ u2.mem\[3\]\[15\] _03269_ _02358_ _03424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_87_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06911_ _02376_ _02390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__09040__I0 _04154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07891_ _03353_ _03354_ _03355_ _03356_ _03357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_110_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09630_ _04526_ _00565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10412__S _05012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06842_ u2.mem\[145\]\[5\] _02082_ _02094_ u2.mem\[168\]\[5\] _02322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_28_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12497__CLK clknet_leaf_175_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07751__B1 _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09561_ _04484_ _00538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06773_ _02251_ _02252_ _02253_ _02254_ _02255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_55_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08512_ _03696_ _03819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10211__I _04886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06306__A1 u2.mem\[178\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09492_ _03985_ _03986_ _04439_ _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_93_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06306__B2 u2.mem\[164\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11150__I1 u2.mem\[146\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08443_ _03774_ _03775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_51_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08374_ _03733_ _00102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08059__A1 _01945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07325_ _02464_ _02800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08854__I0 _04032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_253_clock_I clknet_5_19_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07256_ u2.mem\[18\]\[2\] _02604_ _02606_ u2.mem\[19\]\[2\] _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_137_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06136__I _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10661__I0 _05119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07282__A2 _02659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13122__CLK clknet_leaf_257_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06207_ _01557_ _01618_ _01714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08606__I0 _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07187_ _02641_ _02646_ _02655_ _02664_ _02665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_151_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10169__A2 mem_address_trans\[5\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08351__I _03716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06138_ _01570_ _01644_ _01588_ _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_133_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13272__CLK clknet_leaf_6_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06069_ _01573_ _01575_ _01549_ _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__11118__A1 _05285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06793__A1 u2.mem\[177\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06793__B2 u2.mem\[193\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09031__I0 _04148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09828_ _04602_ u2.mem\[39\]\[11\] _04649_ _04653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07742__B1 _03105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09759_ _04612_ u2.mem\[37\]\[14\] _04606_ _04613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11217__I _03509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12770_ _00649_ clknet_leaf_152_clock u2.mem\[40\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11141__I1 u2.mem\[146\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11721_ _03665_ _05831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11652_ _05787_ _05788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_39_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07430__I _02547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06474__C _01964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10603_ _05133_ _00931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10992__S _05373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11583_ _05744_ _01300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13322_ _01201_ clknet_leaf_322_clock u2.mem\[157\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10652__I0 _05110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10534_ _05018_ u2.mem\[56\]\[11\] _05083_ _05087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10791__I _05231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10465_ _05047_ _00879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13253_ _01132_ clknet_leaf_307_clock u2.mem\[145\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12204_ _00083_ clknet_leaf_271_clock u2.mem\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07025__A2 _02433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13184_ _01063_ clknet_leaf_294_clock u2.mem\[134\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10396_ _05003_ _00854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07576__A3 _03043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12135_ _01461_ clknet_leaf_38_clock u2.driver_mem\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06784__A1 u2.mem\[170\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06784__B2 u2.mem\[156\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09022__I0 _04140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12066_ data_in_trans\[8\].A clknet_leaf_374_clock data_in_trans\[8\].data_sync vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11017_ _05389_ _01089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06536__A1 u2.mem\[176\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09092__I _04181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07733__B1 _03091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06536__B2 u2.mem\[172\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12968_ _00847_ clknet_leaf_128_clock u2.mem\[52\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06839__A2 _02097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11919_ _05909_ u2.mem\[193\]\[2\] _05950_ _05953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12899_ _00778_ clknet_leaf_70_clock u2.mem\[48\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07500__A3 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13145__CLK clknet_leaf_40_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07110_ _02347_ _02589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_119_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10643__I0 _05101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08090_ _01980_ _03526_ _03535_ _00016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11797__I _05878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07041_ _02387_ _02389_ _02406_ _02459_ _02520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_31_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13295__CLK clknet_leaf_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11199__I1 u2.mem\[150\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08992_ _04116_ _00337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06775__A1 u2.mem\[151\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06775__B2 u2.mem\[158\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07943_ u2.mem\[18\]\[14\] _03318_ _03319_ u2.mem\[19\]\[14\] _03408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_25_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11238__S _05529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06790__A4 _02271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07874_ u2.mem\[3\]\[13\] _03269_ _03215_ _03340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06527__A1 _02006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07724__B1 _03072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11371__I1 u2.mem\[160\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09613_ _04491_ u2.mem\[34\]\[12\] _04516_ _04517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06825_ u2.mem\[171\]\[5\] _02066_ _02068_ u2.mem\[157\]\[5\] _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_84_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09544_ _04472_ _00533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08547__S _03840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06756_ _02209_ _02214_ _02223_ _02238_ _02239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09475_ _04430_ _00506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06687_ _02164_ _02165_ _02166_ _02170_ _02171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_149_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08426_ _03697_ u2.mem\[7\]\[9\] _03763_ _03765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08346__I _03712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08357_ _03721_ _03722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12512__CLK clknet_leaf_176_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11587__A1 _04393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11701__S _05818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07308_ _01808_ _02361_ _02762_ _02783_ _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07255__A2 _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08288_ _03665_ _03666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07239_ u2.mem\[49\]\[2\] _02528_ _02532_ u2.mem\[46\]\[2\] _02716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_4_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09177__I _04225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10250_ _04886_ _04914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__12662__CLK clknet_leaf_83_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07007__A2 _02422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10181_ _04869_ _00773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07963__B1 _02501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09905__I _04682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13018__CLK clknet_leaf_149_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07425__I _02552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06469__C _01949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12822_ _00701_ clknet_leaf_89_clock u2.mem\[43\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08457__S _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12042__CLK clknet_leaf_315_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13168__CLK clknet_leaf_279_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09640__I _04521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11114__I1 u2.mem\[144\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12753_ _00632_ clknet_leaf_247_clock u2.mem\[39\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11704_ _05820_ _01345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08256__I _03633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12684_ _00563_ clknet_leaf_216_clock u2.mem\[35\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07160__I _02419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08818__I0 _03936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12192__CLK clknet_leaf_253_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11635_ _05777_ _01319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09288__S _04313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07246__A2 _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11566_ _05715_ u2.mem\[172\]\[3\] _05731_ _05735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_149_clock_I clknet_5_13_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13305_ _01184_ clknet_leaf_376_clock u2.mem\[154\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10517_ _05077_ _00901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11497_ _05663_ u2.mem\[168\]\[0\] _05692_ _05693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13236_ _01115_ clknet_leaf_287_clock u2.mem\[142\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06504__I row_select_trans\[3\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10448_ _05007_ u2.mem\[54\]\[6\] _05035_ _05038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_171_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_170_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13167_ _01046_ clknet_leaf_277_clock u2.mem\[131\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10379_ _04990_ _00850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06757__A1 _01773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12118_ _01481_ clknet_leaf_349_clock u2.select_mem_col\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_201_clock_I clknet_5_31_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13098_ _00977_ clknet_leaf_340_clock u2.mem\[60\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11058__S _05413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12049_ net7 clknet_2_1__leaf_clock_a data_in_trans\[0\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07706__B1 _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11353__I1 u2.mem\[159\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09751__S _04606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10897__S _05310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06610_ u2.mem\[177\]\[0\] _02092_ _02094_ u2.mem\[168\]\[0\] _02095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07590_ u2.mem\[60\]\[8\] _03059_ _03060_ u2.mem\[62\]\[8\] _03061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_92_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06541_ _02016_ _02025_ _02026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_146_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12535__CLK clknet_leaf_110_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09260_ _04265_ u2.mem\[26\]\[6\] _04295_ _04298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08166__I _03584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10864__I0 _05202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06472_ u2.mem\[194\]\[10\] _01946_ _01963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07485__A2 _02908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08211_ _03616_ _00056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09191_ _04249_ _04250_ _04251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08809__I0 _03927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08142_ _03572_ u2.mem\[1\]\[12\] _03573_ _03574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07237__A2 _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12685__CLK clknet_leaf_217_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08073_ _01962_ _03516_ _03523_ _00011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_140_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07024_ _02484_ _02491_ _02496_ _02502_ _02503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_162_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06414__I _01914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11041__I0 _05380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06748__A1 u2.mem\[154\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07945__B1 _02629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06748__B2 u2.mem\[162\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06212__A3 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08975_ _04096_ _04107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_9_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09537__I1 u2.mem\[33\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07926_ u2.mem\[49\]\[14\] _03283_ _03284_ u2.mem\[46\]\[14\] _03391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12065__CLK clknet_2_1__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09661__S _04544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input25_I mem_address_a[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13310__CLK clknet_leaf_363_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07857_ _02618_ _03324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06808_ u2.mem\[155\]\[4\] _02030_ _02192_ u2.mem\[150\]\[4\] _02289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10600__S _05131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07788_ _02402_ _03255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_374_clock clknet_5_1_0_clock clknet_leaf_374_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_37_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09527_ _04389_ u2.mem\[32\]\[14\] _04458_ _04461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_45_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06739_ u2.mem\[177\]\[2\] _02092_ _02089_ u2.mem\[193\]\[2\] _02222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13460__CLK clknet_leaf_360_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09458_ _04360_ u2.mem\[31\]\[1\] _04419_ _04421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08409_ _03755_ _00115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09389_ _04375_ u2.mem\[29\]\[8\] _04376_ _04377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11420_ _05642_ _01239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08804__I _03989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07228__A2 _02457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_150_clock_I clknet_5_24_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06436__B1 _01933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11351_ _05587_ u2.mem\[159\]\[1\] _05598_ _05600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06987__A1 _02421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_312_clock clknet_5_17_0_clock clknet_leaf_312_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_125_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10302_ _04945_ _00818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09225__I0 _04274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11282_ _05556_ u2.mem\[154\]\[5\] _05545_ _05557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13021_ _00900_ clknet_leaf_272_clock u2.mem\[56\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11032__I0 _05388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10233_ _04588_ _04902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06739__A1 u2.mem\[177\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06739__B2 u2.mem\[193\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12408__CLK clknet_leaf_124_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10164_ _04858_ _00767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_327_clock clknet_5_17_0_clock clknet_leaf_327_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_82_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10095_ _04394_ _04760_ _04819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07155__I _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10299__A1 _04072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_10_0_clock clknet_4_5_0_clock clknet_5_10_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__12558__CLK clknet_leaf_203_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06994__I _02346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_75_clock_I clknet_5_8_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10510__S _05073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08187__S _03600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12805_ _00684_ clknet_leaf_88_clock u2.mem\[42\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11405__I _05513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10997_ _05376_ _01082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12736_ _00615_ clknet_leaf_248_clock u2.mem\[38\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12667_ _00546_ clknet_leaf_211_clock u2.mem\[34\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11618_ _05758_ u2.mem\[175\]\[5\] _05760_ _05767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_54_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08714__I _03940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12598_ _00477_ clknet_leaf_97_clock u2.mem\[29\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11549_ _05713_ u2.mem\[171\]\[2\] _05722_ _05725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11140__I _05342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09746__S _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13219_ _01098_ clknet_leaf_301_clock u2.mem\[140\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12088__CLK clknet_leaf_303_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09545__I _04139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11574__I1 u2.mem\[173\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08195__A3 _03482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13333__CLK clknet_leaf_3_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_352_clock_I clknet_5_4_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08760_ _03961_ _03972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07065__I _02543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07711_ u2.mem\[44\]\[10\] _03122_ _03123_ u2.mem\[42\]\[10\] _03180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08691_ _03708_ _03931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13483__CLK clknet_leaf_306_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07642_ _03108_ _03109_ _03110_ _03111_ _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_96_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07573_ _02486_ _03044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09312_ _04312_ _04328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06524_ row_select_trans\[3\].data_sync _02009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09243_ _03581_ _04247_ _04287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06455_ u2.mem\[193\]\[6\] _01942_ _01948_ u2.mem\[192\]\[6\] _01949_ _01950_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_72_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09174_ _04239_ _00396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06386_ u2.mem\[177\]\[5\] _01583_ _01645_ u2.mem\[165\]\[5\] u2.mem\[163\]\[5\]
+ _01643_ _01888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_31_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08125_ _03561_ u2.mem\[1\]\[7\] _03555_ _03562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11262__I0 _05517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07091__B1 _02569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08560__S _03845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08056_ _01878_ _03504_ _03511_ _00006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_122_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07007_ _02473_ _02422_ _02423_ _02485_ _02486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_1_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11714__A1 _04179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09455__I _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06197__A2 _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08958_ _04010_ u2.mem\[20\]\[0\] _04097_ _04098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12700__CLK clknet_leaf_222_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11317__I1 u2.mem\[157\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07909_ u2.mem\[45\]\[14\] _02432_ _02436_ u2.mem\[34\]\[14\] _03374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08889_ _04023_ u2.mem\[18\]\[4\] _04056_ _04057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10330__S _04959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10920_ _04121_ _05317_ _05326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_3958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07697__A2 _03019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09190__I _03987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12850__CLK clknet_leaf_154_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10851_ _05204_ u2.mem\[128\]\[4\] _05277_ _05283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13570_ _01449_ clknet_leaf_13_clock u2.mem\[194\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09694__I0 _04498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10782_ _05231_ _05242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12521_ _00400_ clknet_leaf_125_clock u2.mem\[24\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13206__CLK clknet_leaf_287_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12452_ _00331_ clknet_leaf_90_clock u2.mem\[20\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09446__I0 _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11403_ _05631_ u2.mem\[162\]\[3\] _05625_ _05632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_251_clock clknet_5_19_0_clock clknet_leaf_251_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_165_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12383_ _00262_ clknet_leaf_158_clock u2.mem\[16\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09566__S _04483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12230__CLK clknet_leaf_73_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11334_ _05588_ _01207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07621__A2 _03090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13356__CLK clknet_leaf_377_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10505__S _05066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11265_ _04287_ _05527_ _05545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_4_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09365__I _04127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07909__B1 _02436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_266_clock clknet_5_22_0_clock clknet_leaf_266_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13004_ _00883_ clknet_leaf_273_clock u2.mem\[55\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10216_ _04890_ _00787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11196_ _05499_ _05500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10147_ _04797_ u2.mem\[47\]\[6\] _04846_ _04849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10078_ _04807_ _00732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07137__A1 _02459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08185__I0 _03572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11336__S _05585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07688__A2 _03090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_204_clock clknet_5_31_0_clock clknet_leaf_204_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08645__S _03894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09685__I0 _04489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11492__I0 _05680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08101__A3 _03544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12719_ _00598_ clknet_leaf_250_clock u2.mem\[37\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06112__A2 _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11071__S _05422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06240_ _01617_ _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09437__I0 _04378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_219_clock clknet_5_29_0_clock clknet_leaf_219_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_30_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06171_ _01677_ _01678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_157_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09476__S _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09930_ _04288_ _04659_ _04718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10415__S _05012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12723__CLK clknet_leaf_25_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11547__I1 u2.mem\[171\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09861_ _04672_ _00650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07376__B2 u2.mem\[21\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08812_ _04004_ _00269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09792_ _04632_ _00621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08743_ _03899_ u2.mem\[15\]\[0\] _03962_ _03963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08176__I0 _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11246__S _05528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08674_ _03919_ _00216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07625_ u2.mem\[6\]\[8\] _02927_ _02928_ u2.mem\[47\]\[8\] _03096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12103__CLK clknet_leaf_29_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13229__CLK clknet_leaf_301_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06351__A2 _01639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07556_ _02444_ _03027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06139__I _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09676__I0 _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06507_ row_select_trans\[5\].data_sync row_select_trans\[4\].data_sync _01992_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07487_ u2.mem\[9\]\[6\] _02838_ _02839_ u2.mem\[25\]\[6\] _02960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06103__A2 _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09226_ _04275_ _00412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09428__I0 _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06438_ u2.mem\[192\]\[3\] _01931_ _01936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13379__CLK clknet_leaf_367_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09157_ _04136_ u2.mem\[24\]\[3\] _04226_ _04230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06369_ u2.mem\[146\]\[4\] _01691_ _01693_ u2.mem\[186\]\[4\] _01872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_159_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_23_clock_I clknet_5_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08108_ _03499_ _03550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08290__S _03659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09088_ _04148_ u2.mem\[22\]\[6\] _04187_ _04190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_162_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08039_ data_in_trans\[2\].data_sync _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06811__B1 _02148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10325__S _04954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11050_ _05409_ _01102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06602__I _02086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10001_ _04758_ _00704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07906__A3 _03370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_248_clock_I clknet_5_18_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07119__A1 _02463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08167__I0 _03554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06590__A2 _02037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11156__S _05475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11952_ _05971_ _05972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10903_ _05307_ u2.mem\[131\]\[5\] _05309_ _05316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11883_ u2.mem\[192\]\[2\] _03499_ _05932_ _05933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10834_ _05271_ _01024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09667__I0 _04471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_300_clock_I clknet_5_21_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11474__I0 _05677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13553_ _01432_ clknet_leaf_10_clock u2.mem\[193\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10765_ _05194_ u2.mem\[62\]\[0\] _05232_ _05233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12504_ _00383_ clknet_leaf_126_clock u2.mem\[23\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_190_clock clknet_5_30_0_clock clknet_leaf_190_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09419__I0 _04360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13484_ _01363_ clknet_leaf_306_clock u2.mem\[184\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10696_ _05186_ _00971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12435_ _00314_ clknet_leaf_102_clock u2.mem\[19\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12746__CLK clknet_leaf_44_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12366_ _00245_ clknet_leaf_209_clock u2.mem\[15\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06940__C _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11317_ _05548_ u2.mem\[157\]\[1\] _05576_ _05578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_173_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06802__C2 u2.mem\[192\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12297_ _00176_ clknet_leaf_122_clock u2.mem\[10\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07608__I _02585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11529__I1 u2.mem\[170\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06512__I row_select_trans\[4\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11248_ _05517_ u2.mem\[152\]\[5\] _05528_ _05535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10201__I1 u2.mem\[48\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11179_ _05472_ u2.mem\[148\]\[5\] _05483_ _05490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08158__I0 _03538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12126__CLK clknet_leaf_349_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11066__S _05412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07343__I _02531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11701__I1 u2.mem\[181\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_143_clock clknet_5_13_0_clock clknet_leaf_143_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_91_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07410_ _02500_ _02884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12276__CLK clknet_leaf_100_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08390_ _03726_ _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_95_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13521__CLK clknet_leaf_4_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07341_ u2.mem\[14\]\[4\] _02659_ _02660_ u2.mem\[12\]\[4\] _02816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08086__A2 _03528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_158_clock clknet_5_25_0_clock clknet_leaf_158_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07294__B1 _02577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07272_ u2.mem\[16\]\[3\] _02465_ _02467_ u2.mem\[33\]\[3\] _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07833__A2 _03141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09011_ _04132_ u2.mem\[21\]\[2\] _04124_ _04133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06223_ _01572_ _01729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11768__I1 u2.mem\[185\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06154_ _01660_ _01661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_197_clock_I clknet_5_31_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10145__S _04846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06085_ _01564_ _01591_ _01588_ _01592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_160_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09934__S _04719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09913_ _04706_ _00668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08397__I0 _03722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09844_ _04570_ u2.mem\[40\]\[1\] _04661_ _04663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08010__A2 _03458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09733__I _04566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06021__A1 u2.driver_mem\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09775_ _04617_ _04623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06987_ _02421_ _02433_ _02434_ _02454_ _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_85_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13051__CLK clknet_leaf_264_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08726_ _03925_ u2.mem\[14\]\[9\] _03951_ _03953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12619__CLK clknet_leaf_206_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08657_ _03907_ u2.mem\[13\]\[1\] _03905_ _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_26_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07521__B2 u2.mem\[20\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07608_ _02585_ _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08285__S _03659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08588_ _03814_ u2.mem\[11\]\[7\] _03861_ _03865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07539_ u2.mem\[5\]\[7\] _02922_ _02923_ u2.mem\[38\]\[7\] _03011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_35_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10550_ _04991_ _05097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07824__A2 _03132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09209_ _04263_ u2.mem\[25\]\[5\] _04261_ _04264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10481_ _05001_ u2.mem\[55\]\[4\] _05056_ _05057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12220_ _00099_ clknet_leaf_226_clock u2.mem\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12151_ _00030_ clknet_leaf_56_clock u2.mem\[1\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09844__S _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11102_ _03983_ _03984_ _05274_ _05442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__06260__B2 u2.mem\[154\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12082_ net45 clknet_leaf_380_clock output_active_hold\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12149__CLK clknet_leaf_74_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08388__I0 _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11033_ _05399_ _01095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06012__A1 _01516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06563__A2 _02043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_60_clock clknet_5_12_0_clock clknet_leaf_60_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_91_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12299__CLK clknet_leaf_206_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12984_ _00863_ clknet_leaf_49_clock u2.mem\[53\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13544__CLK clknet_leaf_31_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11695__I0 _05796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11935_ _05216_ u2.mem\[193\]\[9\] _05960_ _05962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07512__A1 _02979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08560__I0 _03823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11614__S _05761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11866_ _05921_ _01406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_75_clock clknet_5_8_0_clock clknet_leaf_75_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_33_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10817_ u2.mem\[63\]\[7\] _03514_ _05258_ _05262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11797_ _05878_ _05879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_13_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07276__B1 _02648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13536_ _01415_ clknet_leaf_345_clock u2.mem\[192\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08923__S _04074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07815__A2 _03125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10748_ _05220_ u2.mem\[61\]\[11\] _05214_ _05221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_173_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13467_ _01346_ clknet_leaf_361_clock u2.mem\[181\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10679_ _05099_ u2.mem\[60\]\[2\] _05174_ _05177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12418_ _00297_ clknet_leaf_171_clock u2.mem\[18\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13398_ _01277_ clknet_leaf_325_clock u2.mem\[169\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12349_ _00228_ clknet_leaf_208_clock u2.mem\[14\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_13_clock clknet_5_2_0_clock clknet_leaf_13_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_138_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08379__I0 _03688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06910_ _02388_ _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_68_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07890_ u2.mem\[57\]\[13\] _02548_ _02550_ u2.mem\[41\]\[13\] _03356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_67_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07200__B1 _02564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06841_ u2.mem\[151\]\[5\] _02085_ _02087_ u2.mem\[158\]\[5\] u2.mem\[193\]\[5\]
+ _02089_ _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_28_clock clknet_5_3_0_clock clknet_leaf_28_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09560_ _04482_ u2.mem\[33\]\[8\] _04483_ _04484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06772_ u2.mem\[184\]\[3\] _02072_ _01994_ _02254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_23_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08511_ _03818_ _00154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09491_ _03983_ mem_address_trans\[5\].data_sync _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07503__A1 u2.mem\[32\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08551__I0 _03814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07503__B2 u2.mem\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12911__CLK clknet_leaf_162_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08442_ mem_address_trans\[2\].data_sync _03773_ _03774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06857__A3 _02323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06711__C1 _02127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11438__I0 _05635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08373_ _03675_ u2.mem\[6\]\[4\] _03732_ _03733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_17_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07267__B1 _02410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07324_ u2.mem\[1\]\[4\] _02797_ _02798_ u2.mem\[7\]\[4\] _02799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_165_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10110__I0 _04797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07806__A2 _03116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07255_ u2.mem\[52\]\[2\] _02599_ _02601_ u2.mem\[21\]\[2\] _02732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_149_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06206_ _01712_ _01713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07186_ _02658_ _02661_ _02662_ _02663_ _02664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_173_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06137_ _01593_ _01644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__11610__I0 _05750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13417__CLK clknet_leaf_314_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06242__A1 u2.mem\[178\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06242__B2 u2.mem\[164\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06152__I _01658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06068_ _01574_ _01575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_87_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06793__A2 _02091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07990__B2 u2.mem\[4\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12441__CLK clknet_leaf_119_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09827_ _04652_ _00636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13567__CLK clknet_leaf_14_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07742__A1 u2.mem\[27\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09758_ _04611_ _04612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08079__I _03492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08709_ _03943_ _00227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09689_ _04560_ _00590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08542__I0 _03805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11434__S _05647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11720_ _05830_ _01351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11651_ _05295_ _05769_ _05787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_14_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07258__B1 _02690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11054__A1 _05411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10602_ _05097_ u2.mem\[58\]\[1\] _05131_ _05133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_74_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10101__I0 _04788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08743__S _03962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11582_ _05717_ u2.mem\[173\]\[4\] _05738_ _05744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13321_ _01200_ clknet_leaf_321_clock u2.mem\[157\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_161_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10533_ _05086_ _00908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13252_ _01131_ clknet_leaf_295_clock u2.mem\[145\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10464_ _05023_ u2.mem\[54\]\[13\] _05045_ _05047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12203_ _00082_ clknet_leaf_229_clock u2.mem\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13097__CLK clknet_leaf_343_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11601__I0 _05756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13183_ _01062_ clknet_leaf_294_clock u2.mem\[134\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10395_ _05001_ u2.mem\[53\]\[4\] _05002_ _05003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06233__B2 u2.mem\[185\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12134_ _01460_ clknet_leaf_12_clock u2.driver_mem\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06784__A2 _02146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06997__I _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12065_ net21 clknet_2_1__leaf_clock_a data_in_trans\[8\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09022__I1 u2.mem\[21\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11016_ _05388_ u2.mem\[138\]\[3\] _05382_ _05389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12934__CLK clknet_leaf_63_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11668__I0 _05798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12967_ _00846_ clknet_leaf_128_clock u2.mem\[52\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11918_ _05952_ _01427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12898_ _00777_ clknet_leaf_245_clock u2.mem\[48\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11849_ _05910_ _01400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11143__I _05345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07249__B1 _02564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12314__CLK clknet_leaf_116_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13519_ _01398_ clknet_leaf_13_clock u2.mem\[190\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_146_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07040_ u2.mem\[44\]\[0\] _02514_ _02518_ u2.mem\[42\]\[0\] _02519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06472__A1 u2.mem\[194\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06224__A1 u2.mem\[163\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12464__CLK clknet_leaf_174_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06224__B2 u2.mem\[165\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08991_ _04048_ u2.mem\[20\]\[15\] _04112_ _04116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_170_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06775__A2 _02084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07942_ u2.mem\[52\]\[14\] _03315_ _03316_ u2.mem\[21\]\[14\] _03407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_151_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09283__I _04310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07873_ u2.mem\[16\]\[13\] _03266_ _03267_ u2.mem\[33\]\[13\] _03339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06527__A2 _02011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08772__I0 _03934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09612_ _04500_ _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_83_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06824_ _01844_ _01996_ _02304_ _01478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08828__S _04015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09543_ _04471_ u2.mem\[33\]\[3\] _04465_ _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11659__I0 _05792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06755_ _02224_ _02231_ _02232_ _02237_ _02238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_110_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11254__S _05537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11284__A1 _04310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09474_ _04375_ u2.mem\[31\]\[8\] _04429_ _04430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_64_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06686_ u2.mem\[146\]\[1\] _02156_ _02158_ u2.mem\[186\]\[1\] _02169_ _02170_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_93_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08425_ _03764_ _00122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08356_ _03720_ _03721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_347_clock_I clknet_5_5_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08563__S _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07307_ _02767_ _02772_ _02777_ _02782_ _02783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__11587__A2 _05729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11831__I0 _05870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10892__I _05309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08287_ _03498_ _03665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07238_ u2.mem\[14\]\[2\] _02659_ _02660_ u2.mem\[12\]\[2\] _02715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07169_ _02492_ _02647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07412__B1 _02809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10180_ _04790_ u2.mem\[48\]\[3\] _04865_ _04869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_65_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12957__CLK clknet_leaf_197_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08763__I0 _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10570__I0 _05110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09921__I _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07191__A2 _02542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12821_ _00700_ clknet_leaf_89_clock u2.mem\[43\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12752_ _00631_ clknet_leaf_247_clock u2.mem\[39\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07441__I _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11703_ _05790_ u2.mem\[181\]\[1\] _05818_ _05820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12337__CLK clknet_leaf_209_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12683_ _00562_ clknet_leaf_211_clock u2.mem\[35\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09569__S _04483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11634_ _05758_ u2.mem\[176\]\[5\] _05770_ _05777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06057__I _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08818__I1 u2.mem\[16\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11565_ _05734_ _01292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09368__I _04131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13304_ _01183_ clknet_leaf_378_clock u2.mem\[154\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12487__CLK clknet_leaf_125_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10516_ _04998_ u2.mem\[56\]\[3\] _05073_ _05077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11496_ _05691_ _05692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_137_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_71_clock_I clknet_5_8_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13235_ _01114_ clknet_leaf_288_clock u2.mem\[142\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10447_ _05037_ _00871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13166_ _01045_ clknet_leaf_277_clock u2.mem\[131\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10378_ _04987_ u2.mem\[53\]\[0\] _04989_ _04990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11339__S _05585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07954__B2 u2.mem\[30\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12117_ _01480_ clknet_leaf_348_clock u2.select_mem_col\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13097_ _00976_ clknet_leaf_343_clock u2.mem\[60\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12048_ col_select_trans\[5\].A clknet_leaf_304_clock col_select_trans\[5\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__11889__I0 u2.mem\[192\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08754__I0 _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_296_clock_I clknet_5_21_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10561__I0 _05103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13112__CLK clknet_leaf_45_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10977__I _05364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07721__A4 _03189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06390__B1 _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08506__I0 _03814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11074__S _05422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06540_ _02024_ _02025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07351__I _02541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06471_ u2.mem\[0\]\[10\] _01962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08210_ _03559_ u2.mem\[3\]\[6\] _03613_ _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09190_ _03987_ _04250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07890__B1 _02550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08809__I1 u2.mem\[16\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08141_ _03545_ _03573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_53_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11813__I0 _05864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10418__S _05012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06445__A1 u2.mem\[192\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08072_ _03522_ _03518_ _03523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06996__A2 _02422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07023_ u2.mem\[54\]\[0\] _02499_ _02501_ u2.mem\[55\]\[0\] _02502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_66_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08974_ _04106_ _00329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07925_ u2.mem\[14\]\[14\] _02521_ _02525_ u2.mem\[12\]\[14\] _03390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_5_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09698__A1 _04121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08745__I0 _03907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07856_ _02616_ _03323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08558__S _03845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09741__I _04598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06807_ u2.mem\[174\]\[4\] _02035_ _02039_ u2.mem\[181\]\[4\] _02288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input18_I data_in_a[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07787_ u2.mem\[32\]\[12\] _03252_ _03253_ u2.mem\[2\]\[12\] _03254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_71_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06920__A2 _02379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09526_ _04460_ _00527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08357__I _03721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06738_ u2.mem\[151\]\[2\] _02085_ _02087_ u2.mem\[158\]\[2\] u2.mem\[168\]\[2\]
+ _02094_ _02221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_43_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09457_ _04420_ _00498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06669_ u2.mem\[179\]\[0\] _02151_ _02153_ u2.mem\[191\]\[0\] _02154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09389__S _04376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08408_ _03663_ u2.mem\[7\]\[1\] _03753_ _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06684__A1 u2.mem\[179\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09388_ _04357_ _04376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07881__B1 _02518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08339_ data_in_trans\[12\].data_sync _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11804__I0 _05872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10328__S _04959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06436__A1 u2.mem\[193\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11350_ _05599_ _01212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06436__B2 u2.mem\[194\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06987__A2 _02433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10301_ _04885_ u2.mem\[51\]\[0\] _04944_ _04945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11281_ _05516_ _05556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13020_ _00899_ clknet_leaf_272_clock u2.mem\[56\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10232_ _04901_ _00792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06739__A2 _02092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10163_ _04813_ u2.mem\[47\]\[13\] _04856_ _04858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_43_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13135__CLK clknet_leaf_330_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10094_ _04818_ _00737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10998__S _05373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10299__A2 _04863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10543__I0 _05027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07164__A2 _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_18_clock_I clknet_5_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13285__CLK clknet_leaf_381_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12804_ _00683_ clknet_leaf_91_clock u2.mem\[42\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10996_ _05343_ u2.mem\[137\]\[2\] _05373_ _05376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12735_ _00614_ clknet_leaf_252_clock u2.mem\[38\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09299__S _04318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12666_ _00545_ clknet_leaf_60_clock u2.mem\[33\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11617_ _05766_ _01312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10238__S _04905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12597_ _00476_ clknet_leaf_97_clock u2.mem\[29\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11548_ _05724_ _01285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11479_ _05681_ _01259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13218_ _01097_ clknet_leaf_290_clock u2.mem\[139\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13149_ _01028_ clknet_leaf_277_clock u2.mem\[128\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07346__I _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12502__CLK clknet_leaf_107_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07710_ _03175_ _03176_ _03177_ _03178_ _03179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_152_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08690_ _03930_ _00221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07641_ u2.mem\[3\]\[9\] _03036_ _02982_ _03111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07572_ u2.mem\[53\]\[8\] _03041_ _03042_ u2.mem\[56\]\[8\] _03043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_53_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07081__I _02446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09311_ _04327_ _00445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06523_ _02007_ _02008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11532__S _05709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09242_ _04286_ _00417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06454_ _01913_ _01949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09173_ _04161_ u2.mem\[24\]\[10\] _04236_ _04239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06385_ _01883_ _01884_ _01885_ _01886_ _01887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_21_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08124_ _03514_ _03561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_147_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11411__A1 _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08055_ _03510_ _03507_ _03511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07006_ _02377_ _02400_ _02392_ _02485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA__09736__I data_in_trans\[9\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12032__CLK clknet_leaf_303_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13158__CLK clknet_leaf_260_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07918__A1 _03379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11714__A2 _05808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07394__A2 _02866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06160__I _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08957_ _04096_ _04097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_88_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12182__CLK clknet_leaf_76_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11707__S _05818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07908_ _01973_ _03250_ _03352_ _03373_ _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10611__S _05136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08888_ _04050_ _04056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_3904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10525__I0 _05009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07146__A2 _02622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07839_ u2.mem\[9\]\[12\] _03304_ _03305_ u2.mem\[25\]\[12\] _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10850_ _05282_ _01029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09143__I0 _04174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09509_ _04371_ u2.mem\[32\]\[6\] _04448_ _04451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10781_ _05241_ _01001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09694__I1 u2.mem\[36\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11442__S _05655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12520_ _00399_ clknet_leaf_124_clock u2.mem\[24\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12451_ _00330_ clknet_leaf_112_clock u2.mem\[20\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09446__I1 u2.mem\[30\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11402_ _05510_ _05631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06409__A1 _01878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12382_ _00261_ clknet_leaf_232_clock u2.mem\[16\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11333_ _05587_ u2.mem\[158\]\[1\] _05585_ _05588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11264_ _05499_ _05544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_4_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13003_ _00882_ clknet_leaf_266_clock u2.mem\[55\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12525__CLK clknet_leaf_198_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10215_ _04889_ u2.mem\[49\]\[1\] _04887_ _04890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11195_ _03490_ _05499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10146_ _04848_ _00759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10521__S _05078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10077_ _04806_ u2.mem\[45\]\[10\] _04802_ _04807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09381__I _04147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07137__A2 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09382__I0 _04371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12675__CLK clknet_leaf_62_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09134__I0 _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10979_ _05366_ _01074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06648__A1 _01992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12718_ _00597_ clknet_leaf_269_clock u2.mem\[37\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11492__I1 u2.mem\[167\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12649_ _00528_ clknet_leaf_114_clock u2.mem\[32\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12055__CLK clknet_2_0__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11244__I1 u2.mem\[152\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06170_ _01608_ _01677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_157_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13300__CLK clknet_leaf_383_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07073__A1 _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06820__A1 u2.mem\[144\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_373_clock clknet_5_1_0_clock clknet_leaf_373_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_154_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08948__I0 _04044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09860_ _04592_ u2.mem\[40\]\[8\] _04671_ _04672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10755__I0 _05225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07076__I _02554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06179__A3 _01587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08811_ _03929_ u2.mem\[16\]\[11\] _04000_ _04004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09791_ _04602_ u2.mem\[38\]\[11\] _04628_ _04632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06584__B1 _02068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08742_ _03961_ _03962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_100_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10431__S _05021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07128__A2 _02604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08673_ _03918_ u2.mem\[13\]\[6\] _03914_ _03919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10132__A1 _04417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_193_clock_I clknet_5_30_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06887__A1 _02339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07624_ u2.mem\[8\]\[8\] _03093_ _03094_ u2.mem\[4\]\[8\] _03095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_53_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_311_clock clknet_5_17_0_clock clknet_leaf_311_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09125__I0 _04148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07555_ _03018_ _03021_ _03024_ _03025_ _03026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_74_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11262__S _05536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06639__A1 u2.mem\[185\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06506_ _01990_ _01991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06639__B2 u2.mem\[173\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07486_ u2.mem\[29\]\[6\] _02835_ _02836_ u2.mem\[11\]\[6\] _02959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_139_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07300__A2 _02604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09225_ _04274_ u2.mem\[25\]\[10\] _04270_ _04275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_326_clock clknet_5_16_0_clock clknet_leaf_326_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06437_ _01773_ _01915_ _01932_ _01935_ _01466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09428__I1 u2.mem\[30\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09667__S _04544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09156_ _04229_ _00388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06368_ u2.mem\[191\]\[4\] _01681_ _01683_ u2.mem\[179\]\[4\] _01871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_148_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08107_ _03549_ _00019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12548__CLK clknet_leaf_100_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07064__A1 _02408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09087_ _04189_ _00359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10606__S _05131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06299_ _01801_ _01802_ _01803_ _01804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_135_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10994__I0 _05340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08038_ _01727_ _03489_ _03497_ _00002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_163_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06811__B2 u2.mem\[156\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08939__I0 _04035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11699__A1 _04120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10000_ _04714_ u2.mem\[43\]\[14\] _04755_ _04758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12698__CLK clknet_leaf_140_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09989_ _04703_ u2.mem\[43\]\[9\] _04750_ _04752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10341__S _04966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06327__B1 _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11951_ _05970_ _05971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11171__I0 _05464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06878__A1 _02347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10902_ _05315_ _01048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11882_ _05928_ _05932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_3789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09116__I0 _04132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10833_ u2.mem\[63\]\[14\] _03532_ _05268_ _05271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12078__CLK clknet_leaf_349_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11474__I1 u2.mem\[166\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13552_ _01431_ clknet_leaf_10_clock u2.mem\[193\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10764_ _05231_ _05232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_164_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13323__CLK clknet_leaf_322_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12503_ _00382_ clknet_leaf_125_clock u2.mem\[23\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13483_ _01362_ clknet_leaf_306_clock u2.mem\[184\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09419__I1 u2.mem\[30\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10695_ _05115_ u2.mem\[60\]\[9\] _05184_ _05186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_16_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12434_ _00313_ clknet_leaf_171_clock u2.mem\[19\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12365_ _00244_ clknet_leaf_210_clock u2.mem\[15\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10516__S _05073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13473__CLK clknet_leaf_308_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11316_ _05577_ _01200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06802__A1 u2.mem\[188\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06802__B2 u2.mem\[187\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12296_ _00175_ clknet_leaf_116_clock u2.mem\[10\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07070__A4 _02546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11247_ _05534_ _01174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07358__A2 _02828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11178_ _05489_ _01150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10251__S _04914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10129_ _04838_ _00752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06318__B1 _01732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11162__I0 _05470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11146__I _05348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_147_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07340_ u2.mem\[44\]\[4\] _02656_ _02657_ u2.mem\[42\]\[4\] _02815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07271_ u2.mem\[1\]\[3\] _02457_ _02461_ u2.mem\[7\]\[3\] _02747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_31_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09010_ _04131_ _04132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06222_ _01565_ _01728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08391__S _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06153_ _01570_ _01622_ _01644_ _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_145_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06084_ _01570_ _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__12840__CLK clknet_leaf_130_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09912_ _04705_ u2.mem\[41\]\[10\] _04701_ _04706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_171_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07349__A2 _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09843_ _04662_ _00642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06021__A2 _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06986_ _02464_ _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09774_ _04622_ _00613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09950__S _04729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08725_ _03952_ _00234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_250_clock clknet_5_19_0_clock clknet_leaf_250_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_113_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08656_ _03662_ _03907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12220__CLK clknet_leaf_226_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13346__CLK clknet_leaf_3_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07607_ u2.mem\[23\]\[8\] _02915_ _02916_ u2.mem\[22\]\[8\] _03078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_42_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08587_ _03864_ _00184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07538_ _03006_ _03007_ _03008_ _03009_ _03010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_168_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_265_clock clknet_5_22_0_clock clknet_leaf_265_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_74_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07469_ u2.mem\[50\]\[6\] _02880_ _02881_ u2.mem\[51\]\[6\] _02942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09208_ _04144_ _04263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10480_ _05050_ _05056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_148_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09139_ _04167_ u2.mem\[23\]\[12\] _04218_ _04219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10967__I0 _05343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08785__A1 _03982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12150_ _00029_ clknet_leaf_74_clock u2.mem\[1\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07052__A4 _02406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11101_ _05441_ _01121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12081_ net46 clknet_leaf_304_clock output_active_hold\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06260__A2 _01715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_203_clock clknet_5_31_0_clock clknet_leaf_203_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10719__I0 _05200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09924__I _04611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08388__I1 u2.mem\[6\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11032_ _05388_ u2.mem\[139\]\[3\] _05395_ _05399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_77_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_150_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10071__S _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_9_clock clknet_5_3_0_clock clknet_leaf_9_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_76_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09860__S _04671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_218_clock clknet_5_29_0_clock clknet_leaf_218_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_64_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12983_ _00862_ clknet_leaf_149_clock u2.mem\[53\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11144__I0 _05468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11934_ _05961_ _01434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11695__I1 u2.mem\[180\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11865_ _05909_ u2.mem\[191\]\[2\] _05918_ _05921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12713__CLK clknet_leaf_146_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08275__I _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10816_ _05261_ _01016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11796_ _04310_ _05847_ _05878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_60_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13535_ _01414_ clknet_leaf_334_clock u2.mem\[192\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10747_ _03703_ _05220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11630__S _05771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13466_ _01345_ clknet_leaf_361_clock u2.mem\[181\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10678_ _05176_ _00963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12863__CLK clknet_leaf_154_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_141_clock_I clknet_5_12_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12417_ _00296_ clknet_leaf_171_clock u2.mem\[18\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13397_ _01276_ clknet_leaf_327_clock u2.mem\[169\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10958__I0 _05352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07619__I _02616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12348_ _00227_ clknet_leaf_207_clock u2.mem\[14\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06787__B1 _02122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13219__CLK clknet_leaf_301_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12279_ _00158_ clknet_leaf_117_clock u2.mem\[9\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09576__I0 _04494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08379__I1 u2.mem\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11383__I0 _05589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11077__S _05422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06679__B _02163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06840_ u2.mem\[165\]\[5\] _02075_ _02078_ u2.mem\[163\]\[5\] _02092_ u2.mem\[177\]\[5\]
+ _02320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_151_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07354__I _02536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07751__A2 _03116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13369__CLK clknet_leaf_371_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06771_ u2.mem\[171\]\[3\] _02065_ _02067_ u2.mem\[157\]\[3\] _02253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11135__I0 _05460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08510_ _03816_ u2.mem\[9\]\[8\] _03817_ _03818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09490_ _04438_ _00513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08386__S _03737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_66_clock_I clknet_5_9_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08441_ mem_address_trans\[3\].data_sync _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_23_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12393__CLK clknet_leaf_140_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06711__B1 _02129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06711__C2 u2.mem\[162\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06857__A4 _02336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08372_ _03726_ _03732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_149_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11438__I1 u2.mem\[164\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09500__I0 _04362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07323_ _02460_ _02798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07267__A1 u2.mem\[40\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07267__B2 u2.mem\[30\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07254_ u2.mem\[17\]\[2\] _02586_ _02591_ u2.mem\[24\]\[2\] _02731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06205_ _01566_ _01586_ _01712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07185_ u2.mem\[43\]\[1\] _02505_ _02508_ u2.mem\[20\]\[1\] _02663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10156__S _04851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06490__A2 _01933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09945__S _04724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06136_ _01642_ _01643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07034__A4 _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06067_ col_select_trans\[1\].data_sync _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_160_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09744__I data_in_trans\[11\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_343_clock_I clknet_5_7_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09826_ _04599_ u2.mem\[39\]\[10\] _04649_ _04652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09319__I0 _04285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07742__A2 _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09757_ data_in_trans\[14\].data_sync _04611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06969_ _02388_ _02448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12736__CLK clknet_leaf_248_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08708_ _03907_ u2.mem\[14\]\[1\] _03941_ _03943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09688_ _04491_ u2.mem\[36\]\[12\] _04559_ _04560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08639_ _03825_ u2.mem\[12\]\[12\] _03894_ _03895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11650_ _05662_ _05786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08095__I _03483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12886__CLK clknet_leaf_71_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10601_ _05132_ _00930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11581_ _05743_ _01299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10532_ _05016_ u2.mem\[56\]\[10\] _05083_ _05086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13320_ _01199_ clknet_leaf_323_clock u2.mem\[156\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08823__I _03987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12116__CLK clknet_leaf_343_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10463_ _05046_ _00878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13251_ _01130_ clknet_leaf_307_clock u2.mem\[145\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12202_ _00081_ clknet_leaf_43_clock u2.mem\[4\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_174_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13182_ _01061_ clknet_leaf_284_clock u2.mem\[133\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10394_ _04988_ _05002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07025__A4 _02417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_142_clock clknet_5_13_0_clock clknet_leaf_142_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12133_ _01459_ clknet_leaf_12_clock u2.driver_mem\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12266__CLK clknet_leaf_54_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12064_ data_in_trans\[7\].A clknet_leaf_374_clock data_in_trans\[7\].data_sync vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13511__CLK clknet_leaf_332_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11365__I0 _05583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11015_ _05345_ _05388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08230__I0 _03579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_157_clock clknet_5_25_0_clock clknet_leaf_157_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_38_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09590__S _04501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07733__A2 _03090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12966_ _00845_ clknet_leaf_105_clock u2.mem\[52\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_161_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11917_ _05907_ u2.mem\[193\]\[1\] _05950_ _05952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12897_ _00776_ clknet_leaf_150_clock u2.mem\[48\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08934__S _04079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11848_ _05909_ u2.mem\[190\]\[2\] _05905_ _05910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_159_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11779_ _05864_ u2.mem\[186\]\[0\] _05866_ _05867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_174_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13518_ _01397_ clknet_leaf_354_clock u2.mem\[189\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_292_clock_I clknet_5_21_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06472__A2 _01946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13449_ _01328_ clknet_leaf_359_clock u2.mem\[178\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13041__CLK clknet_leaf_336_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06224__A2 _01643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08990_ _04115_ _00336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07972__A2 _03425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07941_ u2.mem\[17\]\[14\] _03312_ _03313_ u2.mem\[24\]\[14\] _03406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_142_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08221__I0 _03570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07872_ u2.mem\[1\]\[13\] _03263_ _03264_ u2.mem\[7\]\[13\] _03338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_25_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07185__B1 _02508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07724__A2 _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09611_ _04515_ _00557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06823_ _02285_ _02290_ _02303_ _02304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_7_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11108__I0 _05424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06932__B1 _02410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11535__S _05709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09542_ _04135_ _04471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06754_ u2.mem\[169\]\[2\] _02141_ _02143_ u2.mem\[147\]\[2\] _02236_ _02237_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_71_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09721__I0 _04583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09473_ _04418_ _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_93_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06685_ _02167_ _02168_ _02169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08424_ _03692_ u2.mem\[7\]\[8\] _03763_ _03764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06428__I _01927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12139__CLK clknet_leaf_230_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08355_ data_in_trans\[15\].data_sync _03720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11270__S _05546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07306_ _02778_ _02779_ _02780_ _02781_ _02782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_149_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08286_ _03664_ _00083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11831__I1 u2.mem\[189\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07237_ u2.mem\[44\]\[2\] _02656_ _02657_ u2.mem\[42\]\[2\] _02714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_153_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06463__A2 _01931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12289__CLK clknet_leaf_179_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07168_ _02642_ _02643_ _02644_ _02645_ _02646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_133_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13534__CLK clknet_leaf_333_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07007__A4 _02485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11595__I0 _05752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06119_ _01586_ _01623_ _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_160_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07099_ u2.mem\[9\]\[0\] _02572_ _02577_ u2.mem\[25\]\[0\] _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_156_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_74_clock clknet_5_8_0_clock clknet_leaf_74_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07963__A2 _02499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08212__I0 _03561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07176__B1 _02490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11898__I1 _03520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07715__A2 _03181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09809_ _04642_ _00628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_89_clock clknet_5_11_0_clock clknet_leaf_89_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12820_ _00699_ clknet_leaf_90_clock u2.mem\[43\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09712__I0 _04576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12751_ _00630_ clknet_leaf_247_clock u2.mem\[39\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11702_ _05819_ _01344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_12_clock clknet_5_2_0_clock clknet_leaf_12_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08754__S _03967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12682_ _00561_ clknet_leaf_144_clock u2.mem\[34\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06151__A1 _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07494__A4 _02966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11633_ _05776_ _01318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09649__I _04521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08553__I _03834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11564_ _05713_ u2.mem\[172\]\[2\] _05731_ _05734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13303_ _01182_ clknet_leaf_376_clock u2.mem\[154\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10515_ _05076_ _00900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11495_ _04223_ _05690_ _05691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_clkbuf_leaf_14_clock_I clknet_5_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07169__I _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13234_ _01113_ clknet_leaf_289_clock u2.mem\[142\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10446_ _05005_ u2.mem\[54\]\[5\] _05035_ _05037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10377_ _04988_ _04989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_13165_ _01044_ clknet_leaf_281_clock u2.mem\[131\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_152_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09384__I _04150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12116_ _01479_ clknet_leaf_343_clock u2.select_mem_row\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13096_ _00975_ clknet_leaf_342_clock u2.mem\[60\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08203__I0 _03552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12047_ net6 clknet_2_2__leaf_clock_a col_select_trans\[5\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11889__I1 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07706__A2 _03113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_239_clock_I clknet_5_25_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06390__B2 u2.mem\[188\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12949_ _00828_ clknet_leaf_63_clock u2.mem\[51\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13407__CLK clknet_leaf_320_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06470_ _01958_ _01955_ _01959_ _01961_ _01473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06142__A1 _01613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11090__S _05435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10077__I0 _04806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09559__I _04464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08140_ _03527_ _03572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08463__I _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11813__I1 u2.mem\[188\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12431__CLK clknet_leaf_169_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13557__CLK clknet_leaf_16_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06445__A2 _01931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08071_ data_in_trans\[10\].data_sync _03522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07022_ _02500_ _02501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_146_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12581__CLK clknet_leaf_100_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09294__I _04312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07807__I _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07945__A2 _02627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08973_ _04030_ u2.mem\[20\]\[7\] _04102_ _04106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11329__I _05584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07924_ u2.mem\[44\]\[14\] _02514_ _02518_ u2.mem\[42\]\[14\] _03389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07028__B _02488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07158__B1 _02397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09698__A2 _04542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07855_ u2.mem\[5\]\[12\] _03155_ _03156_ u2.mem\[38\]\[12\] _03322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_83_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06806_ u2.mem\[180\]\[4\] _02043_ _02013_ u2.mem\[172\]\[4\] _02287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_42_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08638__I _03878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07786_ _02396_ _03253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06381__B2 u2.mem\[164\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09525_ _04387_ u2.mem\[32\]\[13\] _04458_ _04460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06737_ u2.mem\[165\]\[2\] _02076_ _02079_ u2.mem\[163\]\[2\] u2.mem\[145\]\[2\]
+ _02081_ _02220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__11501__I0 _05671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13087__CLK clknet_5_19_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_149_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09456_ _04356_ u2.mem\[31\]\[0\] _04419_ _04420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06668_ _02152_ _02153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08407_ _03754_ _00114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09387_ _04153_ _04375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06599_ _02044_ _02057_ _02084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_61_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10609__S _05136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08338_ _03706_ _00093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11804__I1 u2.mem\[187\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07633__A1 u2.mem\[40\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08269_ _03651_ _00079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10408__I _04988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12924__CLK clknet_leaf_221_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10300_ _04943_ _04944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_140_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_188_clock_I clknet_5_30_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11280_ _05555_ _01186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06841__C1 u2.mem\[193\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11568__I0 _05717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10231_ _04900_ u2.mem\[49\]\[6\] _04896_ _04901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08433__I0 _03709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10162_ _04857_ _00766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10093_ _04817_ u2.mem\[45\]\[15\] _04811_ _04818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_120_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08749__S _03962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_240_clock_I clknet_5_25_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12304__CLK clknet_leaf_174_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11175__S _05484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06372__A1 _01867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12803_ _00682_ clknet_leaf_113_clock u2.mem\[42\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10995_ _05375_ _01081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11903__S _05942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12010__D mem_address_trans\[2\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12734_ _00613_ clknet_leaf_270_clock u2.mem\[38\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08484__S _03799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06124__A1 _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06675__A2 _02154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12665_ _00544_ clknet_leaf_141_clock u2.mem\[33\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10519__S _05078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11616_ _05756_ u2.mem\[175\]\[4\] _05760_ _05766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08283__I _03661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12596_ _00475_ clknet_leaf_95_clock u2.mem\[29\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_168_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10318__I _04943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11547_ _05711_ u2.mem\[171\]\[1\] _05722_ _05724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11478_ _05680_ u2.mem\[166\]\[5\] _05664_ _05681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13217_ _01096_ clknet_leaf_295_clock u2.mem\[139\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10254__S _04914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08424__I0 _03692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10429_ _05026_ _00864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07388__B1 _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10231__I0 _04900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13148_ _01027_ clknet_leaf_278_clock u2.mem\[128\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11149__I _05351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13079_ _00958_ clknet_leaf_47_clock u2.mem\[59\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_152_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11731__I0 _05837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07640_ u2.mem\[16\]\[9\] _03033_ _03034_ u2.mem\[33\]\[9\] _03110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_26_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07571_ _02482_ _03042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09310_ _04276_ u2.mem\[27\]\[11\] _04323_ _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06522_ _01988_ _02007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11813__S _05888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09241_ _04285_ u2.mem\[25\]\[15\] _04279_ _04286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06453_ _01918_ _01948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12947__CLK clknet_leaf_65_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09172_ _04238_ _00395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06384_ u2.mem\[184\]\[5\] _01778_ _01753_ _01886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11798__I0 _05864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08123_ _03560_ _00024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08663__I0 _03911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08054_ _03509_ _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07091__A2 _02567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07005_ u2.mem\[53\]\[0\] _02476_ _02483_ u2.mem\[56\]\[0\] _02484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_31_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08415__I0 _03675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06441__I _01914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08956_ _04095_ _03988_ _04096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08569__S _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input30_I mem_address_a[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09915__I0 _04707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07907_ _03357_ _03362_ _03367_ _03372_ _03373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_08887_ _04055_ _00293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11722__I0 _05831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07838_ _02576_ _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06354__A1 u2.mem\[187\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06354__B2 u2.mem\[192\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07769_ u2.mem\[28\]\[11\] _03074_ _03075_ u2.mem\[31\]\[11\] _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_44_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09508_ _04450_ _00519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10780_ _05211_ u2.mem\[62\]\[7\] _05237_ _05241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07854__A1 _03311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09439_ _04380_ u2.mem\[30\]\[10\] _04406_ _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10339__S _04966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12450_ _00329_ clknet_leaf_169_clock u2.mem\[20\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11401_ _05630_ _01232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07606__A1 _03067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06409__A2 _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08654__I0 _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12381_ _00260_ clknet_leaf_232_clock u2.mem\[16\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_166_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09927__I _04614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11332_ _05504_ _05587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13102__CLK clknet_leaf_282_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06290__B1 _01710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10074__S _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08406__I0 _03656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11263_ _05543_ _01181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07909__A2 _02432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13002_ _00881_ clknet_leaf_150_clock u2.mem\[54\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10214_ _04569_ _04889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11194_ _05498_ _01157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10145_ _04795_ u2.mem\[47\]\[5\] _04846_ _04848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13252__CLK clknet_leaf_295_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10802__S _05253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06593__A1 _02006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09906__I0 _04700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10076_ _04598_ _04806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07137__A3 _02615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07542__B1 _02928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_108_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10978_ _05335_ u2.mem\[136\]\[0\] _05365_ _05366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06648__A2 _02052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12717_ _00596_ clknet_leaf_269_clock u2.mem\[37\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08893__I0 _04028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12648_ _00527_ clknet_leaf_114_clock u2.mem\[32\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11994__CLK clknet_leaf_334_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08645__I0 _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12579_ _00458_ clknet_leaf_111_clock u2.mem\[28\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06281__B1 _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09773__S _04618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08948__I1 u2.mem\[19\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08810_ _04003_ _00268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11808__S _05878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09790_ _04631_ _00620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06584__A1 u2.mem\[171\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09572__I _04464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06584__B2 u2.mem\[157\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08741_ _03480_ _03605_ _03606_ _03877_ _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11607__I _05760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_136_clock_I clknet_5_14_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08672_ _03683_ _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06336__A1 u2.mem\[147\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10132__A2 _04760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06336__B2 u2.mem\[169\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07623_ _02611_ _03094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06887__A2 _02338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08089__A1 _03534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07554_ u2.mem\[27\]\[8\] _02871_ _02872_ u2.mem\[35\]\[8\] _03025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_41_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08916__I _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07820__I _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06505_ _01988_ _01989_ _01990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07485_ u2.mem\[26\]\[6\] _02908_ _02909_ u2.mem\[10\]\[6\] _02958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08884__I0 _04019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09224_ _04160_ _04274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07041__B _02406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06436_ u2.mem\[193\]\[2\] _01928_ _01933_ u2.mem\[194\]\[2\] _01934_ _01935_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_22_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13125__CLK clknet_leaf_21_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09155_ _04132_ u2.mem\[24\]\[2\] _04226_ _04229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08636__I0 _03823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06367_ u2.mem\[170\]\[4\] _01686_ _01688_ u2.mem\[156\]\[4\] _01870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_124_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08106_ _03548_ u2.mem\[1\]\[1\] _03546_ _03549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_120_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09086_ _04145_ u2.mem\[22\]\[5\] _04187_ _04189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_162_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06298_ u2.mem\[146\]\[2\] _01692_ _01694_ u2.mem\[186\]\[2\] _01803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06272__B1 _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08037_ _03496_ _03493_ _03497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_162_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06811__A2 _02146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09683__S _04554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09061__I0 _04171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11699__A2 _05808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10622__S _05141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09988_ _04751_ _00698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07772__B1 _03080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09482__I _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08939_ _04035_ u2.mem\[19\]\[9\] _04084_ _04086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10421__I _04988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08098__I mem_address_trans\[1\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11950_ _03582_ _05926_ _05970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06327__A1 u2.mem\[153\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06120__B _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06327__B2 u2.mem\[160\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07524__B1 _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10901_ _05305_ u2.mem\[131\]\[4\] _05309_ _05315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11881_ _05931_ _01411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10832_ _05270_ _01023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13551_ _01430_ clknet_leaf_9_clock u2.mem\[193\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10763_ _04394_ _05172_ _05231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12502_ _00381_ clknet_leaf_107_clock u2.mem\[23\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_338_clock_I clknet_5_18_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13482_ _01361_ clknet_leaf_306_clock u2.mem\[183\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10694_ _05185_ _00970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12433_ _00312_ clknet_leaf_171_clock u2.mem\[19\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08627__I0 _03814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12364_ _00243_ clknet_leaf_210_clock u2.mem\[15\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11315_ _05544_ u2.mem\[157\]\[0\] _05576_ _05577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_5_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06802__A2 _02185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12295_ _00174_ clknet_leaf_117_clock u2.mem\[10\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06081__I _01587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09052__I0 _04164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12642__CLK clknet_leaf_159_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11246_ _05514_ u2.mem\[152\]\[4\] _05528_ _05534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11628__S _05771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10532__S _05083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11177_ _05470_ u2.mem\[148\]\[4\] _05483_ _05489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07763__B1 _03063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10128_ _04815_ u2.mem\[46\]\[14\] _04835_ _04838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_48_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12792__CLK clknet_leaf_339_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07126__B _02424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10059_ _04794_ _00726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06318__A1 u2.mem\[145\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08937__S _04084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06318__B2 u2.mem\[168\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07515__B1 _02809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11162__I1 u2.mem\[147\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06965__B _02442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12022__CLK clknet_leaf_321_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13148__CLK clknet_leaf_278_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07270_ u2.mem\[15\]\[3\] _02445_ _02452_ u2.mem\[13\]\[3\] _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07294__A2 _02572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06221_ _01726_ _01727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12172__CLK clknet_leaf_231_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08618__I0 _03805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13298__CLK clknet_leaf_382_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10425__I0 _05023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06152_ _01658_ _01659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_62_clock_I clknet_5_9_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06083_ u2.mem\[177\]\[0\] _01583_ _01589_ u2.mem\[168\]\[0\] _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_132_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09911_ _04598_ _04705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07349__A3 _02814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11538__S _05708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09842_ _04565_ u2.mem\[40\]\[0\] _04661_ _04662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06557__A1 _02041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09773_ _04576_ u2.mem\[38\]\[3\] _04618_ _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06985_ _02412_ _02413_ _02383_ _02463_ _02464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_80_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08724_ _03922_ u2.mem\[14\]\[8\] _03951_ _03952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_85_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06309__A1 u2.mem\[184\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_287_clock_I clknet_5_20_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_14_0_clock clknet_3_7_0_clock clknet_4_14_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_27_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08655_ _03906_ _00210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11273__S _05546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07606_ _03067_ _03070_ _03073_ _03076_ _03077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_148_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06324__A4 _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08586_ _03812_ u2.mem\[11\]\[6\] _03861_ _03864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_74_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07537_ u2.mem\[18\]\[7\] _02852_ _02853_ u2.mem\[19\]\[7\] _03009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08857__I0 _04035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12515__CLK clknet_leaf_109_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10664__I0 _05121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06166__I _01672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07468_ _02937_ _02938_ _02939_ _02940_ _02941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_09207_ _04262_ _00406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06419_ _01913_ _01920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07399_ u2.mem\[27\]\[5\] _02871_ _02872_ u2.mem\[35\]\[5\] _02873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_10_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09138_ _04202_ _04218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_147_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08381__I _03726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12665__CLK clknet_leaf_141_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09069_ _04177_ u2.mem\[21\]\[15\] _04168_ _04178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11100_ _05432_ u2.mem\[143\]\[5\] _05434_ _05441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12080_ data_in_trans\[15\].A clknet_leaf_348_clock data_in_trans\[15\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11448__S _05655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11031_ _05398_ _01094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07745__B1 _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10151__I _04840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07760__A3 _03222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12982_ _00861_ clknet_leaf_55_clock u2.mem\[53\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12045__CLK clknet_2_2__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09940__I _04718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11144__I1 u2.mem\[146\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11933_ _05213_ u2.mem\[193\]\[8\] _05960_ _05961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11183__S _05492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11864_ _05920_ _01405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06720__A1 _02179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_372_clock clknet_5_1_0_clock clknet_leaf_372_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12195__CLK clknet_leaf_22_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10815_ u2.mem\[63\]\[6\] _03512_ _05258_ _05261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11795_ _05877_ _01379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09588__S _04501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13440__CLK clknet_leaf_354_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10655__I0 _05112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13534_ _01413_ clknet_leaf_333_clock u2.mem\[192\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07276__A2 _02647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10746_ _05219_ _00988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13465_ _01344_ clknet_leaf_362_clock u2.mem\[181\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10677_ _05097_ u2.mem\[60\]\[1\] _05174_ _05176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09387__I _04153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12416_ _00295_ clknet_leaf_170_clock u2.mem\[18\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13396_ _01275_ clknet_leaf_327_clock u2.mem\[169\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12347_ _00226_ clknet_leaf_209_clock u2.mem\[14\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06787__A1 u2.mem\[146\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06787__B2 u2.mem\[173\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_310_clock clknet_5_20_0_clock clknet_leaf_310_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_138_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12278_ _00157_ clknet_leaf_99_clock u2.mem\[9\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11229_ _05511_ u2.mem\[151\]\[3\] _05520_ _05524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07635__I _02425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11383__I1 u2.mem\[161\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07200__A2 _02559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_325_clock clknet_5_16_0_clock clknet_leaf_325_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_27_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06770_ u2.mem\[167\]\[3\] _02059_ _02062_ u2.mem\[183\]\[3\] _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_7_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09850__I _04660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11135__I1 u2.mem\[146\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12538__CLK clknet_leaf_117_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08440_ _03772_ _00129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06711__A1 u2.mem\[154\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08371_ _03731_ _00101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11821__S _05887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09498__S _04443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07322_ _02456_ _02797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10646__I0 _05103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07267__A2 _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12688__CLK clknet_leaf_157_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07253_ u2.mem\[23\]\[2\] _02682_ _02683_ u2.mem\[22\]\[2\] _02730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_165_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10437__S _05030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06204_ u2.mem\[153\]\[0\] _01708_ _01710_ u2.mem\[160\]\[0\] _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07184_ u2.mem\[49\]\[1\] _02528_ _02532_ u2.mem\[46\]\[1\] _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07019__A2 _02422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06714__I _02133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11071__I0 _05420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06135_ _01641_ _01597_ _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06227__B1 _01732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10236__I _04591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09016__I0 _04136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06066_ col_select_trans\[0\].data_sync _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07727__B1 _03149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09961__S _04734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09825_ _04651_ _00635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13313__CLK clknet_leaf_365_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09319__I1 u2.mem\[27\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09756_ _04610_ _00607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08577__S _03856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06968_ _02446_ _02447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__11126__I1 u2.mem\[145\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08707_ _03942_ _00226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09687_ _04543_ _04559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_104_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_2_1__f_clock_a clknet_0_clock_a clknet_2_1__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06899_ _01984_ _02008_ _02378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13463__CLK clknet_leaf_360_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08638_ _03878_ _03894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08569_ _03832_ u2.mem\[10\]\[15\] _03850_ _03854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10600_ _05093_ u2.mem\[58\]\[0\] _05131_ _05132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07258__A2 _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11580_ _05715_ u2.mem\[173\]\[3\] _05739_ _05743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10262__A1 _03583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10531_ _05085_ _00907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13250_ _01129_ clknet_leaf_295_clock u2.mem\[145\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10462_ _05020_ u2.mem\[54\]\[12\] _05045_ _05046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09000__I _04123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12201_ _00080_ clknet_leaf_42_clock u2.mem\[4\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11062__I0 _05388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13181_ _01060_ clknet_leaf_284_clock u2.mem\[133\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_163_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06769__A1 u2.mem\[164\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10393_ _05000_ _05001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11762__A1 _04248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06769__B2 u2.mem\[178\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12132_ _01473_ clknet_leaf_11_clock u2.driver_mem\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12063_ net20 clknet_2_1__leaf_clock_a data_in_trans\[7\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07718__B1 _03060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11365__I1 u2.mem\[160\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11014_ _05387_ _01088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08487__S _03799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_10_clock_I clknet_5_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12965_ _00844_ clknet_leaf_105_clock u2.mem\[52\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07404__B _02749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11916_ _05951_ _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12896_ _00775_ clknet_leaf_245_clock u2.mem\[48\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12830__CLK clknet_leaf_208_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11847_ _03665_ _05909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_92_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07249__A2 _02559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11778_ _05865_ _05866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_60_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13517_ _01396_ clknet_leaf_325_clock u2.mem\[189\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10257__S _04914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10729_ _05207_ u2.mem\[61\]\[5\] _05205_ _05208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_235_clock_I clknet_5_25_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13448_ _01327_ clknet_leaf_359_clock u2.mem\[178\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10005__A1 _04334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06209__B1 _01715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_173_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13379_ _01258_ clknet_leaf_367_clock u2.mem\[166\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13336__CLK clknet_leaf_14_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_173_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07940_ u2.mem\[23\]\[14\] _02594_ _02596_ u2.mem\[22\]\[14\] _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07972__A3 _03430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07709__B1 _03045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_264_clock clknet_5_22_0_clock clknet_leaf_264_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_116_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07871_ u2.mem\[15\]\[13\] _03260_ _03261_ u2.mem\[13\]\[13\] _03337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07185__B2 u2.mem\[20\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12360__CLK clknet_leaf_137_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09610_ _04489_ u2.mem\[34\]\[11\] _04511_ _04515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13486__CLK clknet_leaf_306_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06822_ _02295_ _02300_ _02301_ _02302_ _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_56_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08397__S _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06932__A1 u2.mem\[40\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11108__I1 u2.mem\[144\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06932__B2 u2.mem\[30\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09541_ _04470_ _00532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06753_ _02233_ _02234_ _02235_ _02236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xclkbuf_leaf_279_clock clknet_5_23_0_clock clknet_leaf_279_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_37_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09472_ _04428_ _00505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08196__I _03607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06684_ u2.mem\[179\]\[1\] _02151_ _02153_ u2.mem\[191\]\[1\] _02168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08423_ _03752_ _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06696__B1 _02053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_202_clock clknet_5_29_0_clock clknet_leaf_202_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08354_ _03719_ _00096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09485__I0 _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07305_ u2.mem\[6\]\[3\] _02694_ _02695_ u2.mem\[47\]\[3\] _02781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06448__B1 _01943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11292__I0 _05552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08285_ _03663_ u2.mem\[5\]\[1\] _03659_ _03664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09956__S _04729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_8_clock clknet_5_1_0_clock clknet_leaf_8_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07236_ _02709_ _02710_ _02711_ _02712_ _02713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__08860__S _04033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07660__A2 _03127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_217_clock clknet_5_29_0_clock clknet_leaf_217_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07167_ u2.mem\[3\]\[1\] _02470_ _02359_ _02645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_173_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07948__B1 _02624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11595__I1 u2.mem\[174\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06118_ u2.mem\[167\]\[0\] _01621_ _01624_ u2.mem\[183\]\[0\] _01625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07098_ _02576_ _02577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06049_ _01550_ _01551_ _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_82_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07176__A1 u2.mem\[58\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09808_ _04573_ u2.mem\[39\]\[2\] _04639_ _04642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06923__A1 _02363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09739_ _04597_ _00603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_184_clock_I clknet_5_30_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11525__I _05708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10858__I0 _05194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12750_ _00629_ clknet_leaf_271_clock u2.mem\[39\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07479__A2 _02941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11701_ _05786_ u2.mem\[181\]\[0\] _05818_ _05819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12681_ _00560_ clknet_leaf_144_clock u2.mem\[34\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13209__CLK clknet_leaf_300_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06151__A2 _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11632_ _05756_ u2.mem\[176\]\[4\] _05770_ _05776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09476__I0 _04378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06439__B1 _01933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10077__S _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11563_ _05733_ _01291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07100__A1 _02439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09866__S _04671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13302_ _01181_ clknet_leaf_5_clock u2.mem\[153\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10514_ _04995_ u2.mem\[56\]\[2\] _05073_ _05076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09228__I0 _04276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08770__S _03977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12233__CLK clknet_leaf_54_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11494_ _05605_ _05690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13233_ _01112_ clknet_leaf_303_clock u2.mem\[142\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12008__D mem_address_trans\[1\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10445_ _05036_ _00870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13164_ _01043_ clknet_leaf_285_clock u2.mem\[130\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10376_ _04121_ _04964_ _04988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12115_ _01478_ clknet_leaf_342_clock u2.select_mem_row\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13095_ _00974_ clknet_leaf_342_clock u2.mem\[60\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06303__B _01807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12046_ col_select_trans\[4\].A clknet_leaf_315_clock col_select_trans\[4\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06914__A1 _02390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09106__S _04197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06390__A2 _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10849__I0 _05202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12948_ _00827_ clknet_leaf_64_clock u2.mem\[51\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12879_ _00758_ clknet_leaf_243_clock u2.mem\[47\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06142__A2 _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11371__S _05608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09467__I0 _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07890__A2 _02548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09776__S _04623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09219__I0 _04269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08680__S _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08070_ _01958_ _03516_ _03521_ _00010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07021_ _02477_ _02479_ _02481_ _02458_ _02500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__11026__I0 _05380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06850__B1 _02122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06996__A4 _02474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12726__CLK clknet_leaf_24_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09575__I _04170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08972_ _04105_ _00328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07095__I _02448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12876__CLK clknet_leaf_220_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07923_ _03384_ _03385_ _03386_ _03387_ _03388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_116_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07028__C _02506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07158__A1 u2.mem\[32\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07158__B2 u2.mem\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07854_ _03311_ _03314_ _03317_ _03320_ _03321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_116_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10450__S _05035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06905__A1 _02363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09016__S _04124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06805_ u2.mem\[176\]\[4\] _02003_ _02020_ u2.mem\[189\]\[4\] _02286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07785_ _02384_ _03252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12106__CLK clknet_leaf_47_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09524_ _04459_ _00526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06736_ u2.mem\[166\]\[2\] _02097_ _02099_ u2.mem\[161\]\[2\] _02218_ _02219_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11501__I1 u2.mem\[168\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_141_clock clknet_5_12_0_clock clknet_leaf_141_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09455_ _04418_ _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_101_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06667_ _02104_ _02060_ _02152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_149_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07330__A1 _02796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08406_ _03656_ u2.mem\[7\]\[0\] _03753_ _03754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_40_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09386_ _04374_ _00473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09458__I0 _04360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12256__CLK clknet_leaf_229_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07881__A2 _02514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06598_ u2.mem\[165\]\[0\] _02076_ _02079_ u2.mem\[163\]\[0\] u2.mem\[145\]\[0\]
+ _02082_ _02083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_24_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13501__CLK clknet_leaf_354_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08337_ _03705_ u2.mem\[5\]\[11\] _03693_ _03706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_156_clock clknet_5_24_0_clock clknet_leaf_156_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08268_ _03575_ u2.mem\[4\]\[13\] _03649_ _03651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07219_ _02691_ _02692_ _02693_ _02696_ _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06841__B1 _02087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06987__A4 _02454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06841__C2 _02089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08199_ _03548_ u2.mem\[3\]\[1\] _03608_ _03610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11568__I1 u2.mem\[172\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10230_ _04585_ _04900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_156_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10161_ _04810_ u2.mem\[47\]\[12\] _04856_ _04857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10424__I _03712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10092_ _04614_ _04817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07149__A1 _02443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08197__I0 _03538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13031__CLK clknet_leaf_51_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06372__A2 _01868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12802_ _00681_ clknet_leaf_166_clock u2.mem\[42\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08765__S _03972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10994_ _05340_ u2.mem\[137\]\[1\] _05373_ _05375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_109_clock clknet_5_11_0_clock clknet_leaf_109_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_76_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12733_ _00612_ clknet_leaf_271_clock u2.mem\[38\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06124__A2 _01630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12664_ _00543_ clknet_leaf_141_clock u2.mem\[33\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11256__I0 _05508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11615_ _05765_ _01311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12595_ _00474_ clknet_leaf_112_clock u2.mem\[29\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12749__CLK clknet_leaf_223_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11546_ _05723_ _01284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11477_ _05679_ _05680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_5_22_0_clock_I clknet_4_11_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13216_ _01095_ clknet_leaf_297_clock u2.mem\[139\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10428_ _05025_ u2.mem\[53\]\[14\] _05021_ _05026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_48_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13147_ _01026_ clknet_leaf_262_clock u2.mem\[128\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10359_ _04907_ u2.mem\[52\]\[9\] _04976_ _04978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13078_ _00957_ clknet_leaf_22_clock u2.mem\[59\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12129__CLK clknet_leaf_36_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10270__S _04923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12029_ net39 clknet_2_2__leaf_clock_a row_select_trans\[2\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07643__I _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11731__I1 u2.mem\[182\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07570_ _02475_ _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12279__CLK clknet_leaf_117_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09688__I0 _04491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06521_ _02005_ _02006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13524__CLK clknet_leaf_7_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09240_ _04176_ _04285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06452_ u2.mem\[194\]\[6\] _01946_ _01947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07863__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_73_clock clknet_5_8_0_clock clknet_leaf_73_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_72_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09171_ _04158_ u2.mem\[24\]\[9\] _04236_ _04238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10509__I _05072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06383_ u2.mem\[171\]\[5\] _01611_ _01774_ u2.mem\[157\]\[5\] _01885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08112__I0 _03552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08122_ _03559_ u2.mem\[1\]\[6\] _03555_ _03560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11798__I1 u2.mem\[187\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09860__I0 _04592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_132_clock_I clknet_5_15_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08053_ data_in_trans\[5\].data_sync _03509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_88_clock clknet_5_11_0_clock clknet_leaf_88_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_31_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07004_ _02482_ _02483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_11_clock clknet_5_3_0_clock clknet_leaf_11_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08955_ _04094_ _04095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11276__S _05546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13054__CLK clknet_leaf_274_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07906_ _03368_ _03369_ _03370_ _03371_ _03372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08886_ _04021_ u2.mem\[18\]\[3\] _04051_ _04055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input23_I inverter_select_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11722__I1 u2.mem\[182\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07837_ _02571_ _03304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_26_clock clknet_5_2_0_clock clknet_leaf_26_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06169__I _01675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07768_ u2.mem\[9\]\[11\] _03071_ _03072_ u2.mem\[25\]\[11\] _03236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09679__I0 _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_57_clock_I clknet_5_12_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09507_ _04369_ u2.mem\[32\]\[5\] _04448_ _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11486__I0 _05671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06719_ _02195_ _02197_ _02201_ _02202_ _02203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_38_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07699_ u2.mem\[27\]\[10\] _03104_ _03105_ u2.mem\[35\]\[10\] _03168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09438_ _04408_ _00491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09369_ _04362_ u2.mem\[29\]\[2\] _04358_ _04363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08103__I0 _03538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11400_ _05629_ u2.mem\[162\]\[2\] _05625_ _05630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12380_ _00259_ clknet_leaf_213_clock u2.mem\[16\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09851__I0 _04579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11331_ _05586_ _01206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06290__A1 u2.mem\[153\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06290__B2 u2.mem\[160\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06632__I _02116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11262_ _05517_ u2.mem\[153\]\[5\] _05536_ _05543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13001_ _00880_ clknet_leaf_50_clock u2.mem\[54\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10213_ _04888_ _00786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11193_ _05472_ u2.mem\[149\]\[5\] _05491_ _05498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10144_ _04847_ _00758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06593__A2 _02077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_334_clock_I clknet_5_18_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07790__B2 u2.mem\[30\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10090__S _04811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10075_ _04805_ _00731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12421__CLK clknet_leaf_102_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07137__A4 _02458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13547__CLK clknet_leaf_36_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07542__A1 u2.mem\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06345__A2 _01846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10977_ _05364_ _05365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__12571__CLK clknet_leaf_186_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11713__I _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08294__I _03670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12716_ _00595_ clknet_leaf_269_clock u2.mem\[37\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12647_ _00526_ clknet_leaf_138_clock u2.mem\[32\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12578_ _00457_ clknet_leaf_185_clock u2.mem\[28\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09842__I0 _04565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11529_ _05711_ u2.mem\[170\]\[1\] _05709_ _05712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06281__A1 u2.mem\[175\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06281__B2 u2.mem\[188\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13077__CLK clknet_leaf_22_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07781__A1 _03233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06698__B _01993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06584__A2 _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11096__S _05435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08740_ _03960_ _00241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08671_ _03917_ _00215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06336__A2 _01676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07622_ _02609_ _03093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06887__A3 _02344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07553_ u2.mem\[40\]\[8\] _03022_ _03023_ u2.mem\[30\]\[8\] _03024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_81_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08089__A2 _03528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11623__I _05770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06504_ row_select_trans\[3\].data_sync _01989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07297__B1 _02683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10140__I0 _04790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07484_ _02953_ _02954_ _02955_ _02956_ _02957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_22_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09223_ _04273_ _00411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06435_ _01920_ _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07041__C _02459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09154_ _04228_ _00387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06366_ u2.mem\[173\]\[4\] _01719_ _01721_ u2.mem\[185\]\[4\] _01869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09833__I0 _04609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_10_0_clock clknet_3_5_0_clock clknet_4_10_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA_clkbuf_leaf_283_clock_I clknet_5_22_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08105_ _03496_ _03548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11640__I0 _05750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09085_ _04188_ _00358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06297_ u2.mem\[191\]\[2\] _01682_ _01684_ u2.mem\[179\]\[2\] _01802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07548__I _02384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06272__A1 u2.mem\[167\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08036_ _03495_ _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06272__B2 u2.mem\[183\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10903__S _05309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06024__A1 u2.driver_mem\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12444__CLK clknet_leaf_187_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07221__B1 _02665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09987_ _04700_ u2.mem\[43\]\[8\] _04750_ _04751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08938_ _04085_ _00314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07119__A4 _02488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08869_ _03713_ _04044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_18_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06327__A2 _01707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07524__A1 u2.mem\[61\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10900_ _05314_ _01047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11880_ u2.mem\[192\]\[1\] _03496_ _05929_ _05931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10831_ u2.mem\[63\]\[13\] _03530_ _05268_ _05270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13550_ _01429_ clknet_leaf_8_clock u2.mem\[193\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07288__B1 _02544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10762_ _05230_ _00993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09003__I data_in_trans\[1\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12501_ _00380_ clknet_leaf_119_clock u2.mem\[23\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13481_ _01360_ clknet_leaf_306_clock u2.mem\[183\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10693_ _05112_ u2.mem\[60\]\[8\] _05184_ _05185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12432_ _00311_ clknet_leaf_169_clock u2.mem\[19\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08627__I1 u2.mem\[12\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09824__I0 _04596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_165_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12363_ _00242_ clknet_leaf_234_clock u2.mem\[15\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11314_ _05575_ _05576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12294_ _00173_ clknet_leaf_99_clock u2.mem\[10\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11909__S _05928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12016__D mem_address_trans\[5\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11245_ _05533_ _01173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10198__I0 _04808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06015__A1 u2.driver_mem\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07358__A4 _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11176_ _05488_ _01149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10127_ _04837_ _00751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12937__CLK clknet_leaf_148_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08289__I _03666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07193__I _02547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10058_ _04792_ u2.mem\[45\]\[4\] _04793_ _04794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06318__A2 _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08563__I0 _03825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11644__S _05779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10370__I0 _04918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09114__S _04203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06965__C _02443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07279__B1 _02490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07142__B _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12317__CLK clknet_leaf_186_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06981__B _02458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06220_ u2.mem\[0\]\[1\] _01726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_129_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08618__I1 u2.mem\[12\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09815__I0 _04583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06151_ _01567_ _01609_ _01658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_172_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06254__A1 u2.mem\[187\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06254__B2 u2.mem\[192\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06082_ _01586_ _01588_ _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_160_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11819__S _05888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09910_ _04704_ _00667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10189__I0 _04799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09841_ _04660_ _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07349__A4 _02823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09772_ _04621_ _00612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06984_ _02407_ _02463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_112_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08723_ _03940_ _03951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_113_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11689__I0 _05790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07506__A1 _02974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06309__A2 _01778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08554__I0 _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08654_ _03899_ u2.mem\[13\]\[0\] _03905_ _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08927__I _04073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10361__I0 _04909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07605_ u2.mem\[28\]\[8\] _03074_ _03075_ u2.mem\[31\]\[8\] _03076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08585_ _03863_ _00183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08306__I0 _03680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07536_ u2.mem\[52\]\[7\] _02849_ _02850_ u2.mem\[21\]\[7\] _03008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09959__S _04734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08863__S _04033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06447__I _01923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08857__I1 u2.mem\[17\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07467_ u2.mem\[3\]\[6\] _02803_ _02749_ _02940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11861__I0 _05903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07285__A3 _02759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13242__CLK clknet_leaf_287_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08482__A2 _03544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09206_ _04260_ u2.mem\[25\]\[4\] _04261_ _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09758__I _04611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06418_ _01918_ _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08662__I _03670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07398_ _02425_ _02872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09806__I0 _04570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09137_ _04217_ _00381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06349_ u2.mem\[184\]\[4\] _01778_ _01554_ _01852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_159_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06245__A1 u2.mem\[167\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06182__I _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09068_ _04176_ _04177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06245__B2 u2.mem\[183\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13392__CLK clknet_leaf_369_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07993__A1 _03441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08019_ mem_address_trans\[1\].data_sync _03480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_11_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10633__S _05146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09493__I _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11030_ _05386_ u2.mem\[139\]\[2\] _05395_ _05398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06910__I _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_150_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08103__S _03546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold1_I output_active_hold\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11528__I _05667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08793__I0 _03911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07760__A4 _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12981_ _00860_ clknet_leaf_30_clock u2.mem\[53\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08545__I0 _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11932_ _05949_ _05960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10352__I0 _04900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06705__C1 _02092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11863_ _05907_ u2.mem\[191\]\[1\] _05918_ _05920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10814_ _05260_ _01015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11794_ _05876_ u2.mem\[186\]\[5\] _05865_ _05877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13533_ _01412_ clknet_leaf_333_clock u2.mem\[192\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10745_ _05218_ u2.mem\[61\]\[10\] _05214_ _05219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_159_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10808__S _05253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06484__A1 _01969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07681__B1 _03080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08572__I _03855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13464_ _01343_ clknet_leaf_360_clock u2.mem\[180\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06484__B2 _01972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10676_ _05175_ _00962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12415_ _00294_ clknet_leaf_170_clock u2.mem\[18\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11604__I0 _05758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13395_ _01274_ clknet_leaf_327_clock u2.mem\[169\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07188__I _02552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06236__A1 u2.mem\[146\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12346_ _00225_ clknet_leaf_139_clock u2.mem\[13\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06236__B2 u2.mem\[186\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_179_clock_I clknet_5_27_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06787__A2 _02156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12277_ _00156_ clknet_leaf_104_clock u2.mem\[9\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11907__I1 _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11228_ _05523_ _01166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11159_ _05478_ _01142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_231_clock_I clknet_5_28_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08536__I0 _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10343__I0 _04891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13265__CLK clknet_leaf_311_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06711__A2 _02126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08370_ _03671_ u2.mem\[6\]\[3\] _03727_ _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08683__S _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07321_ u2.mem\[15\]\[4\] _02794_ _02795_ u2.mem\[13\]\[4\] _02796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_149_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09578__I _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06475__A1 _01962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07252_ _02725_ _02726_ _02727_ _02728_ _02729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_143_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06203_ _01709_ _01710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_160_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07183_ u2.mem\[14\]\[1\] _02659_ _02660_ u2.mem\[12\]\[1\] _02661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_157_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07098__I _02576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06227__A1 u2.mem\[193\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06227__B2 u2.mem\[168\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06134_ _01573_ _01574_ _01549_ _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06778__A2 _02257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10453__S _05040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06065_ _01567_ _01571_ _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07826__I _02543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11348__I _05597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09824_ _04596_ u2.mem\[39\]\[9\] _04649_ _04651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06967_ _02386_ _02446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09755_ _04609_ u2.mem\[37\]\[13\] _04606_ _04610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08706_ _03899_ u2.mem\[14\]\[0\] _03941_ _03942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10334__I0 _04920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09686_ _04558_ _00589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06898_ _02376_ _02377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08637_ _03893_ _00205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11039__A1 _04334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06177__I _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08568_ _03853_ _00176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08593__S _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12632__CLK clknet_leaf_112_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07519_ u2.mem\[14\]\[7\] _02892_ _02893_ u2.mem\[12\]\[7\] _02991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_126_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08499_ _03679_ _03810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10530_ _05014_ u2.mem\[56\]\[9\] _05083_ _05085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10262__A2 _04863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10427__I _03716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10461_ _05029_ _05045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_136_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12782__CLK clknet_leaf_268_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12200_ _00079_ clknet_leaf_42_clock u2.mem\[4\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_180_clock_I clknet_5_27_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13180_ _01059_ clknet_leaf_279_clock u2.mem\[133\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10392_ _04138_ _05000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11762__A2 _05847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12131_ _01472_ clknet_leaf_11_clock u2.driver_mem\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10363__S _04976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12012__CLK clknet_leaf_315_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13138__CLK clknet_leaf_330_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12062_ data_in_trans\[6\].A clknet_leaf_374_clock data_in_trans\[6\].data_sync vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11013_ _05386_ u2.mem\[138\]\[2\] _05382_ _05387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07718__B2 u2.mem\[62\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12162__CLK clknet_leaf_236_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13288__CLK clknet_leaf_383_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12964_ _00843_ clknet_leaf_106_clock u2.mem\[52\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10325__I0 _04911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11915_ _05903_ u2.mem\[193\]\[0\] _05950_ _05951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12895_ _00774_ clknet_leaf_245_clock u2.mem\[48\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11846_ _05908_ _01399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11777_ _04287_ _05847_ _05865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11721__I _03665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07654__B1 _03123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13516_ _01395_ clknet_leaf_347_clock u2.mem\[189\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10728_ _05004_ _05207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13447_ _01326_ clknet_leaf_359_clock u2.mem\[178\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10659_ _05117_ u2.mem\[59\]\[10\] _05162_ _05165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06209__A1 u2.mem\[152\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10005__A2 _04760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13378_ _01257_ clknet_leaf_351_clock u2.mem\[166\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11369__S _05608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12329_ _00208_ clknet_leaf_135_clock u2.mem\[12\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10273__S _04928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07646__I _02498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06550__I _02034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07972__A4 _03435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07709__A1 u2.mem\[58\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11168__I _05483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07870_ _03332_ _03333_ _03334_ _03335_ _03336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_9_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10564__I0 _05106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07185__A2 _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_382_clock_I clknet_5_0_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06821_ u2.mem\[185\]\[4\] _02121_ _02123_ u2.mem\[173\]\[4\] _02302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06393__B1 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06932__A2 _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09540_ _04469_ u2.mem\[33\]\[2\] _04465_ _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06752_ u2.mem\[146\]\[2\] _02155_ _02157_ u2.mem\[186\]\[2\] _02235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10316__I0 _04902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09182__I0 _04174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12655__CLK clknet_leaf_236_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09471_ _04373_ u2.mem\[31\]\[7\] _04424_ _04428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06683_ u2.mem\[170\]\[1\] _02146_ _02148_ u2.mem\[156\]\[1\] _02167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_64_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08422_ _03762_ _00121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06696__A1 u2.mem\[164\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06696__B2 u2.mem\[178\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08353_ _03718_ u2.mem\[5\]\[14\] _03710_ _03719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10448__S _05035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07304_ u2.mem\[8\]\[3\] _02610_ _02612_ u2.mem\[4\]\[3\] _02780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_36_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06448__A1 u2.mem\[193\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07645__B1 _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08284_ _03662_ _03663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11292__I1 u2.mem\[155\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06448__B2 u2.mem\[194\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09101__I _04181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07235_ u2.mem\[58\]\[2\] _02487_ _02490_ u2.mem\[36\]\[2\] _02712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_34_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07660__A3 _03128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12035__CLK clknet_2_3__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07166_ u2.mem\[16\]\[1\] _02465_ _02467_ u2.mem\[33\]\[1\] _02644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11279__S _05545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06117_ _01571_ _01623_ _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_145_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07097_ _02573_ _02574_ _02546_ _02575_ _02576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_69_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07556__I _02444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06620__A1 _02056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_371_clock clknet_5_1_0_clock clknet_leaf_371_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06048_ _01554_ _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12185__CLK clknet_leaf_59_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07176__A2 _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09807_ _04641_ _00627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07999_ _01665_ _03462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10710__I _04986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10307__I0 _04893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09738_ _04596_ u2.mem\[37\]\[9\] _04593_ _04597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_127_clock_I clknet_5_15_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09173__I0 _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07479__A3 _02946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09669_ _04543_ _04549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11700_ _05817_ _05818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_27_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12680_ _00559_ clknet_leaf_142_clock u2.mem\[34\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11631_ _05775_ _01317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06439__A1 u2.mem\[193\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07636__B1 _03105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11562_ _05711_ u2.mem\[172\]\[1\] _05731_ _05733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_24_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06439__B2 u2.mem\[194\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10513_ _05075_ _00899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13301_ _01180_ clknet_leaf_0_clock u2.mem\[153\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_324_clock clknet_5_16_0_clock clknet_leaf_324_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11493_ _05689_ _01265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13232_ _01111_ clknet_leaf_302_clock u2.mem\[142\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10444_ _05001_ u2.mem\[54\]\[4\] _05035_ _05036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08987__I0 _04044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11189__S _05492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12528__CLK clknet_leaf_189_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10093__S _04811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13163_ _01042_ clknet_leaf_280_clock u2.mem\[130\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10375_ _04986_ _04987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10794__I0 _05225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12114_ _01477_ clknet_leaf_349_clock u2.select_mem_row\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_339_clock clknet_5_7_0_clock clknet_leaf_339_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_139_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06611__A1 _02006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13094_ _00973_ clknet_leaf_19_clock u2.mem\[60\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08739__I0 _03938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11917__S _05950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12045_ net5 clknet_2_2__leaf_clock_a col_select_trans\[4\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07167__A2 _02470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12678__CLK clknet_leaf_63_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06914__A2 _02391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08297__I _03505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09164__I0 _04148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12947_ _00826_ clknet_leaf_65_clock u2.mem\[51\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08911__I0 _04046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12878_ _00757_ clknet_leaf_225_clock u2.mem\[47\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10268__S _04923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11829_ _05868_ u2.mem\[189\]\[1\] _05896_ _05898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_159_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12058__CLK clknet_leaf_375_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06545__I _02029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_329_clock_I clknet_5_19_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13303__CLK clknet_leaf_376_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07020_ _02498_ _02499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06850__A1 u2.mem\[185\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08760__I _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08978__I0 _04035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13453__CLK clknet_leaf_320_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10785__I0 _05216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08971_ _04028_ u2.mem\[20\]\[6\] _04102_ _04105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11827__S _05896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07922_ u2.mem\[58\]\[14\] _03277_ _03278_ u2.mem\[36\]\[14\] _03387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09147__A3 _03774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10537__I0 _05020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07158__A2 _02385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07853_ u2.mem\[18\]\[12\] _03318_ _03319_ u2.mem\[19\]\[12\] _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_25_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08201__S _03608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06366__B1 _01721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06804_ _02277_ _02282_ _02283_ _02284_ _02285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_151_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07784_ u2.mem\[45\]\[12\] _03099_ _03100_ u2.mem\[34\]\[12\] _03251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09155__I0 _04132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09523_ _04384_ u2.mem\[32\]\[12\] _04458_ _04459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06735_ _02215_ _02216_ _02217_ _02218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06118__B1 _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11562__S _05731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08902__I0 _04037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09454_ _04417_ _04011_ _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06669__A1 u2.mem\[179\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07866__B1 _02436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06666_ _02150_ _02151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06669__B2 u2.mem\[191\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07330__A2 _02799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08405_ _03752_ _03753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_36_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09385_ _04373_ u2.mem\[29\]\[7\] _04367_ _04374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06597_ _02081_ _02082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08336_ _03704_ _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07618__B1 _02923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08267_ _03650_ _00078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09766__I _04617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07218_ u2.mem\[6\]\[1\] _02694_ _02695_ u2.mem\[47\]\[1\] _02696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06841__A1 u2.mem\[151\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08198_ _03609_ _00050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06841__B2 u2.mem\[158\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08969__I0 _04026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_53_clock_I clknet_5_12_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07149_ _02443_ _02614_ _02615_ _02497_ _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_106_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10776__I0 _05207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10160_ _04840_ _04856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_160_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12820__CLK clknet_leaf_90_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11737__S _05840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10091_ _04816_ _00736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10641__S _05152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10528__I0 _05011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07149__A2 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12970__CLK clknet_leaf_127_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_278_clock_I clknet_5_23_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12801_ _00680_ clknet_leaf_166_clock u2.mem\[42\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10993_ _05374_ _01080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12732_ _00611_ clknet_leaf_271_clock u2.mem\[38\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12200__CLK clknet_leaf_42_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12663_ _00542_ clknet_leaf_58_clock u2.mem\[33\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11614_ _05754_ u2.mem\[175\]\[3\] _05761_ _05765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_330_clock_I clknet_5_18_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_263_clock clknet_5_22_0_clock clknet_leaf_263_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_15_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11256__I1 u2.mem\[153\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12594_ _00473_ clknet_leaf_180_clock u2.mem\[29\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12350__CLK clknet_leaf_208_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11545_ _05707_ u2.mem\[171\]\[0\] _05722_ _05723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13476__CLK clknet_leaf_309_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06832__A1 u2.mem\[176\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06832__B2 u2.mem\[189\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11476_ _03509_ _05679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10427_ _03716_ _05025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13215_ _01094_ clknet_leaf_296_clock u2.mem\[139\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_278_clock clknet_5_23_0_clock clknet_leaf_278_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_136_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10767__I0 _05198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07388__A2 _02694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10358_ _04977_ _00842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13146_ _01025_ clknet_leaf_40_clock u2.mem\[63\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_5_26_0_clock_I clknet_4_13_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_201_clock clknet_5_31_0_clock clknet_leaf_201_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10551__S _05095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13077_ _00956_ clknet_leaf_22_clock u2.mem\[59\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10289_ _04937_ _00813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10519__I0 _05001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09385__I0 _04373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12028_ row_select_trans\[1\].A clknet_leaf_304_clock row_select_trans\[1\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06348__B1 _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_7_clock clknet_5_1_0_clock clknet_leaf_7_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_93_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_216_clock clknet_5_29_0_clock clknet_leaf_216_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_25_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09688__I1 u2.mem\[36\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06520_ _02004_ row_select_trans\[4\].data_sync _02005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06451_ _01923_ _01946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09787__S _04628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09170_ _04237_ _00394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06382_ u2.mem\[167\]\[5\] _01749_ _01750_ u2.mem\[183\]\[5\] _01884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08121_ _03512_ _03559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_147_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10726__S _05205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08052_ _01844_ _03504_ _03508_ _00005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__12843__CLK clknet_leaf_214_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07003_ _02477_ _02479_ _02481_ _02401_ _02482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_115_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10758__I0 _05227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12993__CLK clknet_leaf_253_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08954_ _03628_ _03539_ _03632_ _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_170_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07834__I _02558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09027__S _04141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09376__I0 _04366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07905_ u2.mem\[6\]\[13\] _02622_ _02624_ u2.mem\[47\]\[13\] _03371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_29_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08885_ _04054_ _00292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11183__I0 _05460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07836_ u2.mem\[29\]\[12\] _03301_ _03302_ u2.mem\[11\]\[12\] _03303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_3929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12223__CLK clknet_leaf_242_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10930__I0 _05305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input16_I data_in_a[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13349__CLK clknet_leaf_3_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07767_ u2.mem\[29\]\[11\] _03068_ _03069_ u2.mem\[11\]\[11\] _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11292__S _05559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09506_ _04449_ _00518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08665__I _03674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06718_ u2.mem\[176\]\[1\] _02002_ _02012_ u2.mem\[172\]\[1\] _02019_ u2.mem\[189\]\[1\]
+ _02202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_77_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07698_ u2.mem\[40\]\[10\] _03022_ _03023_ u2.mem\[30\]\[10\] _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11486__I1 u2.mem\[167\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09437_ _04378_ u2.mem\[30\]\[9\] _04406_ _04408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06649_ _02014_ _02033_ _02134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07854__A3 _03317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13499__CLK clknet_leaf_329_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11238__I1 u2.mem\[152\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06185__I _01691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09368_ _04131_ _04362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07067__A1 _02428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08319_ _03690_ _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09299_ _04265_ u2.mem\[27\]\[6\] _04318_ _04321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09851__I1 u2.mem\[40\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11330_ _05583_ u2.mem\[158\]\[0\] _05585_ _05586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08106__S _03546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06814__B2 u2.mem\[147\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06290__A2 _01708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11261_ _05542_ _01180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10212_ _04885_ u2.mem\[49\]\[0\] _04887_ _04888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13000_ _00879_ clknet_leaf_338_clock u2.mem\[54\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11192_ _05497_ _01156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10143_ _04792_ u2.mem\[47\]\[4\] _04846_ _04847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10074_ _04804_ u2.mem\[45\]\[9\] _04802_ _04805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11266__I _05545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08776__S _03977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07542__A2 _02927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06750__B1 _02147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10976_ _04224_ _05363_ _05364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_71_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12715_ _00594_ clknet_leaf_268_clock u2.mem\[37\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11930__S _05955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11229__I1 u2.mem\[151\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06095__I _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12646_ _00525_ clknet_leaf_94_clock u2.mem\[32\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12866__CLK clknet_leaf_154_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12577_ _00456_ clknet_leaf_182_clock u2.mem\[28\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09842__I1 u2.mem\[40\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10988__I0 _05352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06805__A1 u2.mem\[176\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11528_ _05667_ _05711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06805__B2 u2.mem\[189\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07073__A4 _02430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08007__B1 _03462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11459_ _05666_ _01254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_140_clock clknet_5_12_0_clock clknet_leaf_140_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_124_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13129_ _01008_ clknet_leaf_342_clock u2.mem\[62\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09358__I0 _04285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12246__CLK clknet_leaf_73_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07781__A2 _03238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input8_I data_in_a[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08670_ _03916_ u2.mem\[13\]\[5\] _03914_ _03917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08686__S _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_155_clock clknet_5_24_0_clock clknet_leaf_155_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_113_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10912__I0 _05301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07621_ u2.mem\[39\]\[8\] _03090_ _03091_ u2.mem\[48\]\[8\] _03092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_26_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12396__CLK clknet_leaf_193_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07552_ _02409_ _03023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06503_ row_select_trans\[2\].data_sync _01988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07483_ u2.mem\[57\]\[6\] _02904_ _02905_ u2.mem\[41\]\[6\] _02956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_34_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06219__B _01725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09222_ _04272_ u2.mem\[25\]\[9\] _04270_ _04273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06434_ _01923_ _01933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09310__S _04323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09153_ _04128_ u2.mem\[24\]\[1\] _04226_ _04228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_124_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06365_ u2.mem\[144\]\[4\] _01670_ _01672_ u2.mem\[182\]\[4\] _01868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_159_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_226_clock_I clknet_5_28_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08104_ _03547_ _00018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07829__I _02538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09084_ _04140_ u2.mem\[22\]\[4\] _04187_ _04188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11640__I1 u2.mem\[177\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06296_ u2.mem\[170\]\[2\] _01687_ _01689_ u2.mem\[156\]\[2\] _01801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07064__A4 _02406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08035_ data_in_trans\[1\].data_sync _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13021__CLK clknet_leaf_272_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06272__A2 _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09597__I0 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_108_clock clknet_5_11_0_clock clknet_leaf_108_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_162_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07221__A1 _01726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06024__A2 _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07221__B2 _02698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09986_ _04739_ _04750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_107_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07772__A2 _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09349__I0 _04276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09980__S _04745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13171__CLK clknet_leaf_281_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08937_ _04032_ u2.mem\[19\]\[8\] _04084_ _04085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11156__I0 _05464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12739__CLK clknet_leaf_29_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08868_ _04043_ _00286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10903__I0 _05307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07524__A2 _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07819_ _02504_ _03286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08799_ _03997_ _00263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10830_ _05269_ _01022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06908__I _02386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12889__CLK clknet_leaf_52_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10761_ _05229_ u2.mem\[61\]\[15\] _05223_ _05230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11750__S _05849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12500_ _00379_ clknet_leaf_108_clock u2.mem\[23\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13480_ _01359_ clknet_leaf_303_clock u2.mem\[183\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10692_ _05173_ _05184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_41_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12431_ _00310_ clknet_leaf_169_clock u2.mem\[19\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12119__CLK clknet_leaf_343_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12362_ _00241_ clknet_leaf_137_clock u2.mem\[14\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07055__A4 _02533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07460__A1 u2.mem\[32\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11313_ _05411_ _05566_ _05575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_12293_ _00172_ clknet_leaf_98_clock u2.mem\[10\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12269__CLK clknet_leaf_194_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09588__I0 _04467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11244_ _05511_ u2.mem\[152\]\[3\] _05529_ _05533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06799__B _01993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11175_ _05468_ u2.mem\[148\]\[3\] _05484_ _05488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10126_ _04813_ u2.mem\[46\]\[13\] _04835_ _04837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_72_clock clknet_5_8_0_clock clknet_leaf_72_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_79_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07763__A2 _03062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11147__I0 _05470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10057_ _04783_ _04793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_94_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_175_clock_I clknet_5_27_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_87_clock clknet_5_11_0_clock clknet_leaf_87_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11724__I _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07279__A1 u2.mem\[58\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07142__C _02450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10959_ _05353_ _01067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_10_clock clknet_5_3_0_clock clknet_leaf_10_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_149_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09130__S _04213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06981__C _02459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12629_ _00508_ clknet_leaf_96_clock u2.mem\[31\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13044__CLK clknet_leaf_33_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09815__I1 u2.mem\[39\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06150_ _01656_ _01657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_25_clock clknet_5_2_0_clock clknet_leaf_25_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_144_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07451__A1 u2.mem\[39\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06081_ _01587_ _01588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_172_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09579__I0 _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13194__CLK clknet_leaf_287_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10189__I1 u2.mem\[48\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09840_ _04224_ _04659_ _04660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09771_ _04573_ u2.mem\[38\]\[2\] _04618_ _04621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06983_ u2.mem\[1\]\[0\] _02457_ _02461_ u2.mem\[7\]\[0\] _02462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11138__I0 _05464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11835__S _05895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08722_ _03950_ _00233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11689__I1 u2.mem\[180\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09751__I0 _04605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08653_ _03904_ _03905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_27_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07604_ _02581_ _03075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08584_ _03810_ u2.mem\[11\]\[5\] _03861_ _03863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_81_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06190__A1 u2.mem\[147\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07535_ u2.mem\[17\]\[7\] _02846_ _02847_ u2.mem\[24\]\[7\] _03007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11570__S _05730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07466_ u2.mem\[16\]\[6\] _02800_ _02801_ u2.mem\[33\]\[6\] _02939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_167_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11861__I1 u2.mem\[191\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09040__S _04155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09205_ _04251_ _04261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_139_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06417_ _01911_ _01916_ _01918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07397_ _02419_ _02871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_377_clock_I clknet_5_0_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07559__I _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09975__S _04740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09136_ _04164_ u2.mem\[23\]\[11\] _04213_ _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06348_ u2.mem\[171\]\[4\] _01611_ _01774_ u2.mem\[157\]\[4\] _01851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12411__CLK clknet_leaf_190_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13537__CLK clknet_leaf_34_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09067_ data_in_trans\[15\].data_sync _04176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08490__I0 _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06279_ _01781_ _01782_ _01783_ _01784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10914__S _05319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07993__A2 _03446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08018_ _03478_ _03479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_150_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12561__CLK clknet_leaf_161_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07745__A2 _03030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_8_0_clock clknet_3_4_0_clock clknet_4_8_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_09969_ _04681_ u2.mem\[43\]\[0\] _04740_ _04741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_4202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12980_ _00859_ clknet_leaf_67_clock u2.mem\[53\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09742__I0 _04599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11931_ _05959_ _01433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10352__I1 u2.mem\[52\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11544__I _05721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06705__C2 u2.mem\[177\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06638__I _02122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06181__A1 _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11862_ _05919_ _01404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09014__I _04134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10813_ u2.mem\[63\]\[5\] _03510_ _05258_ _05260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11301__I0 _05544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11793_ _03678_ _05876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09949__I _04718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13532_ _01411_ clknet_leaf_349_clock u2.mem\[192\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08853__I _04014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10744_ _03699_ _05218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07681__A1 u2.mem\[17\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13463_ _01342_ clknet_leaf_360_clock u2.mem\[180\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10675_ _05093_ u2.mem\[60\]\[0\] _05174_ _05175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12414_ _00293_ clknet_leaf_191_clock u2.mem\[18\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12091__CLK clknet_2_2__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13394_ _01273_ clknet_leaf_328_clock u2.mem\[169\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12345_ _00224_ clknet_leaf_61_clock u2.mem\[13\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10824__S _05263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12904__CLK clknet_leaf_52_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12276_ _00155_ clknet_leaf_100_clock u2.mem\[9\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11227_ _05508_ u2.mem\[151\]\[2\] _05520_ _05523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10040__I0 _04716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07736__A2 _03202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11158_ _05466_ u2.mem\[147\]\[2\] _05475_ _05478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10109_ _04827_ _00743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11089_ _05434_ _05435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_49_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09125__S _04208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10343__I1 u2.mem\[52\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11454__I _03490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08964__S _04097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06172__A1 _01678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06992__B _02359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07320_ _02451_ _02795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09110__A1 _03751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09859__I _04660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12434__CLK clknet_leaf_171_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07251_ u2.mem\[28\]\[2\] _02580_ _02582_ u2.mem\[31\]\[2\] _02728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_32_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06475__A2 _01955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06202_ _01596_ _01635_ _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07182_ _02524_ _02660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_129_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07019__A4 _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06133_ _01639_ _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12584__CLK clknet_leaf_110_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09594__I _04500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06064_ _01547_ _01570_ _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_144_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11359__I0 _05595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08224__I0 _03572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07727__A2 _03148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10031__I0 _04707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09823_ _04650_ _00634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09754_ _04608_ _04609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06966_ _02444_ _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09035__S _04141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08705_ _03940_ _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_95_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09685_ _04489_ u2.mem\[36\]\[11\] _04554_ _04558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06897_ _02352_ _02375_ _02376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11364__I _05607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08636_ _03823_ u2.mem\[12\]\[11\] _03889_ _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06163__A1 _01612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08567_ _03830_ u2.mem\[10\]\[14\] _03850_ _03853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07518_ u2.mem\[44\]\[7\] _02889_ _02890_ u2.mem\[42\]\[7\] _02990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_126_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08498_ _03809_ _00150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07449_ _02628_ _02923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_168_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12927__CLK clknet_leaf_242_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10460_ _05044_ _00877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11598__I0 _05754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_123_clock_I clknet_5_15_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09119_ _04207_ _00373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10391_ _04999_ _00853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10270__I0 _04893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07966__A2 _03427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12130_ _01471_ clknet_leaf_35_clock u2.driver_mem\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08215__I0 _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10443__I _05029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12061_ net19 clknet_2_1__leaf_clock_a data_in_trans\[6\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10022__I0 _04698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09009__I _04130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07718__A2 _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09963__I0 _04714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11012_ _05342_ _05386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12307__CLK clknet_leaf_111_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11770__I0 _05833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12963_ _00842_ clknet_leaf_110_clock u2.mem\[52\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11914_ _05949_ _05950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_111_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12457__CLK clknet_leaf_128_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12894_ _00773_ clknet_leaf_224_clock u2.mem\[48\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_48_clock_I clknet_5_7_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11845_ _05907_ u2.mem\[190\]\[1\] _05905_ _05908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11776_ _03654_ _05864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13515_ _01394_ clknet_leaf_347_clock u2.mem\[189\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10727_ _05206_ _00982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13446_ _01325_ clknet_leaf_352_clock u2.mem\[177\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10658_ _05164_ _00955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11589__I0 _05746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10554__S _05095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13377_ _01256_ clknet_leaf_8_clock u2.mem\[166\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10589_ _03712_ _05124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12328_ _00207_ clknet_leaf_136_clock u2.mem\[12\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10961__A1 _05354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08206__I0 _03554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12259_ _00138_ clknet_leaf_23_clock u2.mem\[8\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10013__I0 _04689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09954__I0 _04705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07709__A2 _03044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_325_clock_I clknet_5_16_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13232__CLK clknet_leaf_302_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06820_ u2.mem\[144\]\[4\] _02115_ _02117_ u2.mem\[182\]\[4\] _02301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06393__A1 u2.mem\[166\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06393__B2 u2.mem\[161\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07662__I _02552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07590__B1 _03060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06751_ u2.mem\[179\]\[2\] _02150_ _02152_ u2.mem\[191\]\[2\] _02234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11513__I0 _05668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09470_ _04427_ _00504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06682_ u2.mem\[185\]\[1\] _02121_ _02123_ u2.mem\[173\]\[1\] _02166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_149_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13382__CLK clknet_leaf_319_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08421_ _03688_ u2.mem\[7\]\[7\] _03758_ _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06696__A2 _02050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10729__S _05205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08352_ _03717_ _03718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07303_ u2.mem\[39\]\[3\] _02617_ _02619_ u2.mem\[48\]\[3\] _02779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06448__A2 _01942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08283_ _03661_ _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07234_ u2.mem\[53\]\[2\] _02476_ _02483_ u2.mem\[56\]\[2\] _02711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07165_ u2.mem\[1\]\[1\] _02457_ _02461_ u2.mem\[7\]\[1\] _02643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10464__S _05045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07837__I _02571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07948__A2 _02622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06116_ _01622_ _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06605__C1 u2.mem\[193\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08070__A1 _01958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07096_ _02347_ _02575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_117_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10263__I _04922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06047_ _01553_ _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_160_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06620__A2 _02104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09945__I0 _04696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11752__I0 _05829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09806_ _04570_ u2.mem\[39\]\[1\] _04639_ _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06384__A1 u2.mem\[184\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07998_ _01547_ _03461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07581__B1 _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09737_ _04595_ _04596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06949_ _02348_ _02415_ _02428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09668_ _04548_ _00581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07479__A4 _02951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08619_ _03883_ _00197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10639__S _05152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09599_ _04478_ u2.mem\[34\]\[6\] _04506_ _04509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11630_ _05754_ u2.mem\[176\]\[3\] _05771_ _05775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06916__I _02394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08109__S _03546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07636__A1 u2.mem\[27\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11561_ _05732_ _01290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13300_ _01179_ clknet_leaf_383_clock u2.mem\[153\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10512_ _04992_ u2.mem\[56\]\[1\] _05073_ _05075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13105__CLK clknet_leaf_329_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11492_ _05680_ u2.mem\[167\]\[5\] _05682_ _05689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_274_clock_I clknet_5_23_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13231_ _01110_ clknet_leaf_302_clock u2.mem\[142\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10443_ _05029_ _05035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_137_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07747__I _02357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13162_ _01041_ clknet_leaf_279_clock u2.mem\[130\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08061__A1 _03514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10374_ _04117_ _04986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11269__I _05504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10173__I _04864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12113_ _01476_ clknet_leaf_345_clock u2.select_mem_row\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06611__A2 _02046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13255__CLK clknet_leaf_286_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13093_ _00972_ clknet_leaf_20_clock u2.mem\[60\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09936__I0 _04687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08739__I1 u2.mem\[14\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12044_ col_select_trans\[3\].A clknet_leaf_315_clock col_select_trans\[3\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11743__I0 _05835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_5_0_clock clknet_0_clock clknet_3_5_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_66_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07572__B1 _03042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06914__A3 _02392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12946_ _00825_ clknet_leaf_151_clock u2.mem\[51\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07875__A1 _03337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06678__A2 _02074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12877_ _00756_ clknet_leaf_224_clock u2.mem\[47\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11828_ _05897_ _01392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11997__CLK clknet_leaf_34_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07627__A1 _03066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11759_ _05854_ _01366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10284__S _04933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13429_ _01308_ clknet_leaf_350_clock u2.mem\[175\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06850__A2 _02120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10234__I0 _04902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08052__A1 _01844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11982__I0 _05225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10785__I1 u2.mem\[62\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10083__I _04783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08970_ _04104_ _00327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08689__S _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07921_ u2.mem\[53\]\[14\] _03274_ _03275_ u2.mem\[56\]\[14\] _03386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_29_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12622__CLK clknet_leaf_201_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07852_ _02605_ _03319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07392__I _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06366__B2 u2.mem\[185\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06803_ u2.mem\[165\]\[4\] _02076_ _02079_ u2.mem\[163\]\[4\] u2.mem\[145\]\[4\]
+ _02082_ _02284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput1 col_select_a[0] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_07783_ _02360_ _03250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09522_ _04442_ _04458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__12772__CLK clknet_leaf_64_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06734_ u2.mem\[159\]\[2\] _02174_ _02176_ u2.mem\[149\]\[2\] _02217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06118__A1 u2.mem\[167\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06118__B2 u2.mem\[183\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09453_ _04416_ _04417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10459__S _05040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06665_ _01998_ _02077_ _02150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_164_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08404_ _03479_ _03751_ _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_7_0_clock clknet_4_3_0_clock clknet_5_7_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_09384_ _04150_ _04373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13128__CLK clknet_leaf_39_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12002__CLK clknet_leaf_41_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06596_ _02023_ _02080_ _02081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_5_0_0_clock_I clknet_4_0_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08335_ _03703_ _03704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08266_ _03572_ u2.mem\[4\]\[12\] _03649_ _03650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12152__CLK clknet_leaf_65_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07217_ _02623_ _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_165_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13278__CLK clknet_leaf_8_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08197_ _03538_ u2.mem\[3\]\[0\] _03608_ _03609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10225__I0 _04895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08969__I1 u2.mem\[20\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07148_ _02626_ _02627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_173_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11089__I _05434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11973__I0 _05216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10776__I1 u2.mem\[62\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07079_ _02522_ _02523_ _02430_ _02506_ _02558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__10922__S _05327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10090_ _04815_ u2.mem\[45\]\[14\] _04811_ _04816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_121_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11725__I0 _05833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07149__A3 _02615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10721__I _04997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07554__B1 _02872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12800_ _00679_ clknet_leaf_166_clock u2.mem\[42\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10992_ _05335_ u2.mem\[137\]\[0\] _05373_ _05374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_16_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12731_ _00610_ clknet_leaf_266_clock u2.mem\[38\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12662_ _00541_ clknet_leaf_83_clock u2.mem\[33\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06646__I _02130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11613_ _05764_ _01310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08657__I0 _03907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12593_ _00472_ clknet_leaf_161_clock u2.mem\[29\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10464__I0 _05023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11544_ _05721_ _05722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_51_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11475_ _05678_ _01258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13214_ _01093_ clknet_leaf_297_clock u2.mem\[139\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10426_ _05024_ _00863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08034__A1 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12645__CLK clknet_leaf_94_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11964__I0 _05915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11928__S _05955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12035__D net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13145_ _01024_ clknet_leaf_40_clock u2.mem\[63\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10357_ _04904_ u2.mem\[52\]\[8\] _04976_ _04977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09909__I0 _04703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13076_ _00955_ clknet_leaf_26_clock u2.mem\[59\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10288_ _04911_ u2.mem\[50\]\[11\] _04933_ _04937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11716__I0 _05825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11727__I _03673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12795__CLK clknet_leaf_184_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12027_ net38 clknet_2_2__leaf_clock_a row_select_trans\[1\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06348__A1 u2.mem\[171\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07545__B1 _02995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12025__CLK clknet_2_3__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12929_ _00808_ clknet_leaf_151_clock u2.mem\[50\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10279__S _04928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06450_ u2.mem\[0\]\[6\] _01945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_107_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_370_clock clknet_5_1_0_clock clknet_leaf_370_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_15_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12175__CLK clknet_leaf_236_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06381_ u2.mem\[178\]\[5\] _01746_ _01747_ u2.mem\[164\]\[5\] _01883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08120_ _03558_ _00023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10455__I0 _05014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08051_ _03506_ _03507_ _03508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_174_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07002_ _02480_ _02481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__10207__I0 _04817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13570__CLK clknet_leaf_13_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11955__I0 _05907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08820__I0 _03938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07784__B1 _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09308__S _04323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08953_ _04093_ _00321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11707__I0 _05794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11637__I _05778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07904_ u2.mem\[8\]\[13\] _03326_ _03327_ u2.mem\[4\]\[13\] _03370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_44_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08884_ _04019_ u2.mem\[18\]\[2\] _04051_ _04054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06339__A1 _01809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11183__I1 u2.mem\[149\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_222_clock_I clknet_5_29_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07835_ _02563_ _03302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_323_clock clknet_5_16_0_clock clknet_leaf_323_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_42_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07766_ u2.mem\[26\]\[11\] _03141_ _03142_ u2.mem\[10\]\[11\] _03234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_25_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09505_ _04366_ u2.mem\[32\]\[4\] _04448_ _04449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_77_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06717_ u2.mem\[194\]\[1\] _02198_ _02199_ u2.mem\[190\]\[1\] _02200_ u2.mem\[160\]\[1\]
+ _02201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_37_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07697_ u2.mem\[32\]\[10\] _03019_ _03020_ u2.mem\[2\]\[10\] _03166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09978__S _04745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09436_ _04407_ _00490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08882__S _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_338_clock clknet_5_18_0_clock clknet_leaf_338_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_25_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06648_ _01992_ _02052_ _02133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07854__A4 _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09367_ _04361_ _00467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08639__I0 _03825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06579_ _02056_ _02064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10446__I0 _05005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08318_ data_in_trans\[8\].data_sync _03690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07067__A2 _02377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09298_ _04320_ _00439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12668__CLK clknet_leaf_217_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08249_ _03640_ _00070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11260_ _05514_ u2.mem\[153\]\[4\] _05536_ _05542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11946__I0 _05227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10211_ _04886_ _04887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_134_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08811__I0 _03929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11191_ _05470_ u2.mem\[149\]\[4\] _05491_ _05497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06578__A1 u2.mem\[167\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06578__B2 u2.mem\[183\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10142_ _04840_ _04846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_97_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10073_ _04595_ _04804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12048__CLK clknet_leaf_304_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07527__B1 _02905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08856__I _03696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06750__A1 u2.mem\[170\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06750__B2 u2.mem\[156\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10099__S _04820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12198__CLK clknet_leaf_22_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10975_ _05275_ _05363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__13443__CLK clknet_leaf_363_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_56_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12714_ _00593_ clknet_leaf_146_clock u2.mem\[36\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06376__I _01877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12645_ _00524_ clknet_leaf_94_clock u2.mem\[32\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09687__I _04543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10437__I0 _04992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12576_ _00455_ clknet_leaf_184_clock u2.mem\[28\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06266__B1 _01737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11527_ _05710_ _01278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10626__I _05130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_171_clock_I clknet_5_26_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11458_ _05663_ u2.mem\[166\]\[0\] _05665_ _05666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11937__I0 _05218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10409_ _05011_ u2.mem\[53\]\[8\] _05012_ _05013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08802__I0 _03920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11389_ _05595_ u2.mem\[161\]\[5\] _05615_ _05622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07766__B1 _03142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13128_ _01007_ clknet_leaf_39_clock u2.mem\[62\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07230__A2 _02470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07781__A3 _03243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13059_ _00938_ clknet_leaf_31_clock u2.mem\[58\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07518__B1 _02890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07620_ _02618_ _03091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06741__A1 u2.mem\[144\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06741__B2 u2.mem\[182\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_31_0_clock clknet_4_15_0_clock clknet_5_31_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_07551_ _02402_ _03022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_96_clock_I clknet_5_10_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09798__S _04633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06502_ _01985_ _01986_ _01987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07297__A2 _02682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07482_ u2.mem\[37\]\[6\] _02829_ _02830_ u2.mem\[59\]\[6\] _02955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09221_ _04157_ _04272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12810__CLK clknet_leaf_130_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06433_ u2.mem\[192\]\[2\] _01931_ _01932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10428__I0 _05025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09152_ _04227_ _00386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06364_ u2.mem\[154\]\[4\] _01699_ _01701_ u2.mem\[162\]\[4\] _01866_ _01867_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_08103_ _03538_ u2.mem\[1\]\[0\] _03546_ _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06257__C2 u2.mem\[181\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09083_ _04181_ _04187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10536__I _05072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06295_ u2.mem\[173\]\[2\] _01720_ _01722_ u2.mem\[185\]\[2\] _01800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_148_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12960__CLK clknet_leaf_168_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08034_ _01545_ _03489_ _03494_ _00001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_11_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11928__I0 _05209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11568__S _05730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10472__S _05051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07757__B1 _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07845__I _02585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13316__CLK clknet_leaf_316_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09985_ _04749_ _00697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08936_ _04073_ _04084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11156__I1 u2.mem\[147\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_262_clock clknet_5_22_0_clock clknet_leaf_262_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_135_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_373_clock_I clknet_5_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08867_ _04041_ u2.mem\[17\]\[12\] _04042_ _04043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12340__CLK clknet_leaf_94_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13466__CLK clknet_leaf_361_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07818_ u2.mem\[49\]\[12\] _03283_ _03284_ u2.mem\[46\]\[12\] _03285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_131_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07580__I _02531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08798_ _03916_ u2.mem\[16\]\[5\] _03995_ _03997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06732__A1 u2.mem\[187\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06732__B2 u2.mem\[192\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07749_ _03212_ _03213_ _03214_ _03216_ _03217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xclkbuf_leaf_277_clock clknet_5_23_0_clock clknet_leaf_277_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_72_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06196__I _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07288__A2 _02542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10760_ _03720_ _05229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12490__CLK clknet_leaf_127_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09419_ _04360_ u2.mem\[30\]\[1\] _04396_ _04398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_160_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_4_0_clock clknet_3_2_0_clock clknet_4_4_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_9_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10691_ _05183_ _00969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_200_clock clknet_5_31_0_clock clknet_leaf_200_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_12_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12430_ _00309_ clknet_leaf_191_clock u2.mem\[19\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06924__I _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08237__A1 _03629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11092__I0 _05424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12361_ _00240_ clknet_leaf_136_clock u2.mem\[14\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06799__A1 u2.mem\[184\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11312_ _05574_ _01199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_6_clock clknet_5_1_0_clock clknet_leaf_6_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12292_ _00171_ clknet_leaf_99_clock u2.mem\[10\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_215_clock clknet_5_29_0_clock clknet_leaf_215_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_5_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11919__I0 _05909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09588__I1 u2.mem\[34\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10382__S _04989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11243_ _05532_ _01172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11174_ _05487_ _01148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06420__B1 _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10125_ _04836_ _00750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08787__S _03990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11147__I1 u2.mem\[146\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10056_ _04578_ _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_169_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07704__B _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06723__A1 u2.mem\[167\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_118_clock_I clknet_5_14_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07920__B1 _02501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06723__B2 u2.mem\[183\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12833__CLK clknet_5_26_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07279__A2 _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10958_ _05352_ u2.mem\[134\]\[5\] _05336_ _05353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09411__S _04385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06487__B1 _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10557__S _05095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10889_ _05307_ u2.mem\[130\]\[5\] _05296_ _05308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12983__CLK clknet_leaf_149_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12628_ _00507_ clknet_leaf_95_clock u2.mem\[31\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09276__I0 _04281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10356__I _04965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12559_ _00438_ clknet_leaf_159_clock u2.mem\[27\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12213__CLK clknet_leaf_23_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06080_ _01550_ _01579_ _01587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_89_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13339__CLK clknet_leaf_1_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07739__B1 _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12363__CLK clknet_leaf_234_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13489__CLK clknet_leaf_306_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09770_ _04620_ _00611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06982_ _02460_ _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11138__I1 u2.mem\[146\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08721_ _03920_ u2.mem\[14\]\[7\] _03946_ _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08496__I _03798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08652_ _03479_ _03903_ _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10897__I0 _05301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09751__I1 u2.mem\[37\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07603_ _02579_ _03074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08583_ _03862_ _00182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06190__A2 _01676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07534_ u2.mem\[23\]\[7\] _02915_ _02916_ u2.mem\[22\]\[7\] _03006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06478__B1 _01948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07465_ u2.mem\[1\]\[6\] _02797_ _02798_ u2.mem\[7\]\[6\] _02938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09204_ _04139_ _04260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06416_ _01916_ _01917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09267__I0 _04272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07396_ u2.mem\[40\]\[5\] _02789_ _02790_ u2.mem\[30\]\[5\] _02870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09120__I _04202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09135_ _04216_ _00380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09967__A1 _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11074__I0 _05424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06347_ u2.mem\[167\]\[4\] _01749_ _01750_ u2.mem\[183\]\[4\] _01850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_147_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07978__B1 _02569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09066_ _04175_ _00352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06278_ u2.mem\[172\]\[2\] _01654_ _01666_ u2.mem\[150\]\[2\] _01783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06650__B1 _02134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08017_ _03477_ mem_address_trans\[5\].data_sync mem_address_trans\[6\].data_sync
+ mem_address_trans\[7\].data_sync _03478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__07993__A3 _03451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09991__S _04750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06402__B1 _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09968_ _04739_ _04740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_103_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10930__S _05326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08919_ _04010_ u2.mem\[19\]\[0\] _04074_ _04075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12856__CLK clknet_leaf_143_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09899_ _04696_ u2.mem\[41\]\[6\] _04692_ _04697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11930_ _05211_ u2.mem\[193\]\[7\] _05955_ _05959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06705__A1 u2.mem\[165\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07902__B1 _02629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06705__B2 u2.mem\[163\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11861_ _05903_ u2.mem\[191\]\[0\] _05918_ _05919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06181__A2 _01630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10812_ _05259_ _01014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06720__A4 _02203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11792_ _05875_ _01378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11301__I1 u2.mem\[156\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06469__B1 _01943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13531_ _01410_ clknet_leaf_348_clock u2.mem\[192\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10743_ _05217_ _00987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12236__CLK clknet_leaf_226_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13462_ _01341_ clknet_leaf_360_clock u2.mem\[180\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07681__A2 _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09258__I0 _04263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10674_ _05173_ _05174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09030__I _04147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12413_ _00292_ clknet_leaf_193_clock u2.mem\[18\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13393_ _01272_ clknet_leaf_327_clock u2.mem\[169\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_154_clock clknet_5_24_0_clock clknet_leaf_154_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12344_ _00223_ clknet_leaf_86_clock u2.mem\[13\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07433__A2 _02902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_44_clock_I clknet_5_6_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12275_ _00154_ clknet_leaf_111_clock u2.mem\[9\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11226_ _05522_ _01165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09430__I0 _04371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_169_clock clknet_5_26_0_clock clknet_leaf_169_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07736__A3 _03203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11157_ _05477_ _01141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10108_ _04795_ u2.mem\[46\]\[5\] _04825_ _04827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11088_ _04417_ _05402_ _05434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_114_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10039_ _04780_ _00720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_269_clock_I clknet_5_23_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09205__I _04251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13011__CLK clknet_leaf_30_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_107_clock clknet_5_11_0_clock clknet_leaf_107_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_63_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09141__S _04218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07121__A1 _02560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07250_ u2.mem\[9\]\[2\] _02572_ _02577_ u2.mem\[25\]\[2\] _02727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_143_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09249__I0 _04254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08980__S _04107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_321_clock_I clknet_5_16_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13161__CLK clknet_leaf_279_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11056__I0 _05380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06201_ _01707_ _01708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10086__I _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07181_ _02520_ _02659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_160_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12729__CLK clknet_leaf_45_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06132_ _01567_ _01576_ _01639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_145_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07424__A2 _02879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06063_ _01569_ _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11359__I1 u2.mem\[159\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12879__CLK clknet_leaf_243_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09421__I0 _04362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09822_ _04592_ u2.mem\[39\]\[8\] _04649_ _04650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09753_ data_in_trans\[13\].data_sync _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06965_ _02439_ _02440_ _02442_ _02443_ _02444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_171_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08704_ _03606_ _03725_ _03877_ _03940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_09684_ _04557_ _00588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06148__C1 u2.mem\[172\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06896_ _02341_ _02342_ _02375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08635_ _03892_ _00204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06163__A2 _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08566_ _03852_ _00175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12259__CLK clknet_leaf_23_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13504__CLK clknet_leaf_333_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07517_ _02985_ _02986_ _02987_ _02988_ _02989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_39_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08497_ _03807_ u2.mem\[9\]\[4\] _03808_ _03809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08160__I0 _03548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07448_ _02626_ _02922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_167_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_71_clock clknet_5_8_0_clock clknet_leaf_71_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_126_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11047__I0 _05388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07379_ u2.mem\[18\]\[4\] _02852_ _02853_ u2.mem\[19\]\[4\] _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_10_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11598__I1 u2.mem\[174\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09118_ _04136_ u2.mem\[23\]\[3\] _04203_ _04207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10390_ _04998_ u2.mem\[53\]\[3\] _04989_ _04999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06218__A3 _01724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09049_ _04162_ _00348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_86_clock clknet_5_9_0_clock clknet_leaf_86_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_108_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10724__I _05000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12060_ data_in_trans\[5\].A clknet_leaf_375_clock data_in_trans\[5\].data_sync vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11756__S _05849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11011_ _05385_ _01087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06387__C1 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11770__I1 u2.mem\[185\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13034__CLK clknet_leaf_51_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12962_ _00841_ clknet_leaf_168_clock u2.mem\[52\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_270_clock_I clknet_5_23_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09025__I _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11913_ _04013_ _05926_ _05949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_24_clock clknet_5_2_0_clock clknet_leaf_24_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12893_ _00772_ clknet_leaf_224_clock u2.mem\[48\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11844_ _03661_ _05907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13184__CLK clknet_leaf_294_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11286__I0 _05544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11775_ _05863_ _01373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08151__I0 _03579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11986__A1 _03534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13514_ _01393_ clknet_leaf_346_clock u2.mem\[189\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10726_ _05204_ u2.mem\[61\]\[4\] _05205_ _05206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_39_clock clknet_5_6_0_clock clknet_leaf_39_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07654__A2 _03122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_1_0_clock clknet_0_clock clknet_3_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_13445_ _01324_ clknet_leaf_352_clock u2.mem\[177\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10835__S _05268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10657_ _05115_ u2.mem\[59\]\[9\] _05162_ _05164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_167_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13376_ _01255_ clknet_leaf_8_clock u2.mem\[166\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10588_ _05123_ _00926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12327_ _00206_ clknet_leaf_138_clock u2.mem\[12\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12258_ _00137_ clknet_leaf_241_clock u2.mem\[8\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11209_ _03501_ _05510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10570__S _05104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12189_ _00068_ clknet_leaf_267_clock u2.mem\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06378__C1 _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09136__S _04213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11465__I _05670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06393__A2 _01592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07590__B2 u2.mem\[62\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06750_ u2.mem\[170\]\[2\] _02145_ _02147_ u2.mem\[156\]\[2\] _02233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_95_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06559__I _02022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12401__CLK clknet_leaf_172_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11513__I1 u2.mem\[169\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13527__CLK clknet_leaf_325_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06681_ u2.mem\[144\]\[1\] _02115_ _02117_ u2.mem\[182\]\[1\] _02165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08420_ _03761_ _00120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_0_0_clock_I clknet_3_0_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08351_ _03716_ _03717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12551__CLK clknet_leaf_123_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08142__I0 _03572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07302_ u2.mem\[5\]\[3\] _02689_ _02690_ u2.mem\[38\]\[3\] _02778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06508__B _01992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08282_ _03495_ _03661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07645__A2 _03113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07233_ u2.mem\[54\]\[2\] _02650_ _02651_ u2.mem\[55\]\[2\] _02710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06853__B1 _02157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07164_ u2.mem\[15\]\[1\] _02445_ _02452_ u2.mem\[13\]\[1\] _02642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08215__S _03618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06605__B1 _02087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06115_ _01580_ _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_173_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06605__C2 _02089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07095_ _02448_ _02574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__08070__A2 _03516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06046_ _01547_ _01549_ _01552_ _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_5_3_0_clock clknet_4_1_0_clock clknet_5_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_82_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11576__S _05739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13057__CLK clknet_leaf_256_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11752__I1 u2.mem\[184\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07030__B1 _02508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09805_ _04640_ _00626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input39_I row_select_a[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07997_ u2.active_mem\[4\] _03458_ _03459_ u2.active_mem\[5\] _03460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_47_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06384__A2 _01778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06948_ u2.mem\[27\]\[0\] _02420_ _02426_ u2.mem\[35\]\[0\] _02427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06923__A4 _02401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09736_ data_in_trans\[9\].data_sync _04595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12081__CLK clknet_leaf_304_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09667_ _04471_ u2.mem\[36\]\[3\] _04544_ _04548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06879_ _02357_ _02358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08618_ _03805_ u2.mem\[12\]\[3\] _03879_ _03883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09598_ _04508_ _00551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08549_ _03812_ u2.mem\[10\]\[6\] _03840_ _03843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_93_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11560_ _05707_ u2.mem\[172\]\[0\] _05731_ _05732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07636__A2 _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10511_ _05074_ _00898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06844__B1 _02116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11491_ _05688_ _01264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10655__S _05162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_217_clock_I clknet_5_29_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13230_ _01109_ clknet_leaf_290_clock u2.mem\[141\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10442_ _05034_ _00869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07939__A3 _03402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13161_ _01040_ clknet_leaf_279_clock u2.mem\[130\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10373_ _04985_ _00849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12112_ _01475_ clknet_leaf_347_clock u2.select_mem_row\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13092_ _00971_ clknet_leaf_26_clock u2.mem\[60\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11486__S _05683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10390__S _04989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12043_ net4 clknet_2_2__leaf_clock_a col_select_trans\[3\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08859__I _03700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11743__I1 u2.mem\[183\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12424__CLK clknet_leaf_121_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11285__I _05558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12945_ _00824_ clknet_leaf_151_clock u2.mem\[51\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12876_ _00755_ clknet_leaf_220_clock u2.mem\[47\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06678__A3 _02113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11827_ _05864_ u2.mem\[189\]\[0\] _05896_ _05897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07627__A2 _03077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11758_ _05835_ u2.mem\[184\]\[4\] _05848_ _05854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_18_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08824__A1 _03482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10709_ _05193_ _00977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11689_ _05790_ u2.mem\[180\]\[1\] _05810_ _05812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_146_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13428_ _01307_ clknet_leaf_352_clock u2.mem\[174\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_2_0__f_clock_a clknet_0_clock_a clknet_2_0__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_155_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13359_ _01238_ clknet_leaf_373_clock u2.mem\[163\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07260__B1 _02612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07920_ u2.mem\[54\]\[14\] _02499_ _02501_ u2.mem\[55\]\[14\] _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08769__I _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07012__B1 _02490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07851_ _02603_ _03318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11195__I _03490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06366__A2 _01719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06802_ u2.mem\[188\]\[4\] _02185_ _02186_ u2.mem\[187\]\[4\] _02187_ u2.mem\[192\]\[4\]
+ _02283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__12917__CLK clknet_leaf_88_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06905__A4 _02383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07782_ _01966_ _03017_ _03228_ _03249_ _01488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xinput2 col_select_a[1] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_56_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09521_ _04457_ _00525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06733_ u2.mem\[188\]\[2\] _02185_ _02177_ u2.mem\[175\]\[2\] _02216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_77_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06118__A2 _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11923__I _05949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_166_clock_I clknet_5_26_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09452_ _03747_ _03901_ _04416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_149_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06664_ u2.mem\[170\]\[0\] _02146_ _02148_ u2.mem\[156\]\[0\] _02149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07866__A2 _02432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08403_ _03750_ _03751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09383_ _04372_ _00472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06595_ _01991_ _02017_ _02080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08334_ data_in_trans\[11\].data_sync _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07618__A2 _02922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08265_ _03633_ _03649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_119_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07848__I _02598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_4_0_clock_I clknet_4_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07216_ _02621_ _02694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_153_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09615__I0 _04494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08196_ _03607_ _03608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07147_ _02560_ _02561_ _02474_ _02562_ _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_118_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_5_26_0_clock clknet_4_13_0_clock clknet_5_26_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11973__I1 u2.mem\[194\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12447__CLK clknet_leaf_168_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07251__B1 _02582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07078_ _02540_ _02545_ _02551_ _02556_ _02557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06029_ u2.driver_mem\[12\] _01522_ _01537_ _01519_ _01538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08679__I _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07583__I _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11725__I1 u2.mem\[182\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07149__A4 _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07554__A1 u2.mem\[27\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06420__C _01920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09719_ _04143_ _04582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10991_ _05372_ _05373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_16_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12730_ _00609_ clknet_leaf_47_clock u2.mem\[37\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10161__I0 _04810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09303__I _04312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12661_ _00540_ clknet_leaf_76_clock u2.mem\[33\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08106__I0 _03548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11612_ _05752_ u2.mem\[175\]\[2\] _05761_ _05764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_24_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12592_ _00471_ clknet_leaf_161_clock u2.mem\[29\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11543_ _04310_ _05690_ _05721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13222__CLK clknet_leaf_300_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_368_clock_I clknet_5_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06293__A1 u2.mem\[154\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07490__B1 _02916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09606__I0 _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06293__B2 u2.mem\[162\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11474_ _05677_ u2.mem\[166\]\[4\] _05664_ _05678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13213_ _01092_ clknet_leaf_296_clock u2.mem\[139\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10425_ _05023_ u2.mem\[53\]\[13\] _05021_ _05024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11413__I0 _05623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11964__I1 u2.mem\[194\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13144_ _01023_ clknet_leaf_41_clock u2.mem\[63\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10356_ _04965_ _04976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_151_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13372__CLK clknet_leaf_371_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06596__A2 _02080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13075_ _00954_ clknet_leaf_25_clock u2.mem\[59\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10287_ _04936_ _00812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12026_ row_select_trans\[0\].A clknet_leaf_304_clock row_select_trans\[0\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07545__A1 _01951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06348__A2 _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08593__I0 _03819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07545__B2 _03016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06330__C _01833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11944__S _05965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12928_ _00807_ clknet_leaf_243_clock u2.mem\[50\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10152__I0 _04801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12859_ _00738_ clknet_leaf_211_clock u2.mem\[46\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06520__A2 row_select_trans\[4\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06380_ _01879_ _01880_ _01881_ _01882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_33_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06808__B1 _02192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10295__S _04938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07668__I _02549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08050_ _03492_ _03507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06284__B2 u2.mem\[161\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06823__A3 _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07001_ _02372_ _02480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07233__B1 _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11955__I1 u2.mem\[194\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_92_clock_I clknet_5_10_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08952_ _04048_ u2.mem\[19\]\[15\] _04089_ _04093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08499__I _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11707__I1 u2.mem\[181\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07903_ u2.mem\[39\]\[13\] _03323_ _03324_ u2.mem\[48\]\[13\] _03369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08883_ _04053_ _00291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07536__A1 u2.mem\[52\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08584__I0 _03810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11854__S _05904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07834_ _02558_ _03301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07765_ _03229_ _03230_ _03231_ _03232_ _03233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_09504_ _04442_ _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06716_ _02137_ _02200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07696_ u2.mem\[45\]\[10\] _03099_ _03100_ u2.mem\[34\]\[10\] _03165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10143__I0 _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09435_ _04375_ u2.mem\[30\]\[8\] _04406_ _04407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06647_ u2.mem\[148\]\[0\] _02129_ _02131_ u2.mem\[152\]\[0\] _02132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13245__CLK clknet_leaf_307_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09366_ _04360_ u2.mem\[29\]\[1\] _04358_ _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_24_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06578_ u2.mem\[167\]\[0\] _02059_ _02062_ u2.mem\[183\]\[0\] _02063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08317_ _03689_ _00089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09297_ _04263_ u2.mem\[27\]\[5\] _04318_ _04320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07067__A3 _02429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08248_ _03554_ u2.mem\[4\]\[4\] _03639_ _03640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13395__CLK clknet_leaf_327_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08179_ _03597_ _00043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09793__I _04617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10210_ _04013_ _04863_ _04886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07224__B1 _02410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11190_ _05496_ _01155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07775__A1 _03239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10141_ _04845_ _00757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_0_0_clock clknet_3_0_0_clock clknet_4_0_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_10072_ _04803_ _00730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08575__I0 _03801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11764__S _05857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10382__I0 _04992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08327__I0 _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06750__A2 _02145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06657__I _02141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10134__I0 _04782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10974_ _05362_ _01073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09033__I data_in_trans\[7\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12713_ _00592_ clknet_leaf_146_clock u2.mem\[36\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09968__I _04739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08872__I _03717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12644_ _00523_ clknet_leaf_94_clock u2.mem\[32\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12612__CLK clknet_leaf_82_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11634__I0 _05758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12575_ _00454_ clknet_leaf_184_clock u2.mem\[28\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10907__I _05318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06266__A1 _01727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11526_ _05707_ u2.mem\[170\]\[0\] _05709_ _05710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_114_clock_I clknet_5_14_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08007__A2 _03461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11457_ _05664_ _05665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10843__S _05278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12762__CLK clknet_leaf_51_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07215__B1 _02612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10408_ _04988_ _05012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__11937__I1 u2.mem\[193\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11388_ _05621_ _01228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07766__A1 u2.mem\[26\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10339_ _04885_ u2.mem\[52\]\[0\] _04966_ _04967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13127_ _01006_ clknet_leaf_39_clock u2.mem\[62\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09208__I _04144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13118__CLK clknet_leaf_276_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13058_ _00937_ clknet_leaf_250_clock u2.mem\[58\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_152_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11674__S _05801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12009_ net26 clknet_2_1__leaf_clock_a mem_address_trans\[2\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12142__CLK clknet_leaf_230_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13268__CLK clknet_leaf_384_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07550_ u2.mem\[32\]\[8\] _03019_ _03020_ u2.mem\[2\]\[8\] _03021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_4_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_39_clock_I clknet_5_6_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06501_ row_select_trans\[1\].data_sync _01986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10089__I _04611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07481_ u2.mem\[60\]\[6\] _02826_ _02827_ u2.mem\[62\]\[6\] _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09220_ _04271_ _00410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06432_ _01919_ _01931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08782__I mem_address_trans\[7\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12292__CLK clknet_leaf_99_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09151_ _04119_ u2.mem\[24\]\[0\] _04226_ _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06363_ _01863_ _01864_ _01865_ _01866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_72_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07398__I _02425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08102_ _03545_ _03546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09082_ _04186_ _00357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06257__B2 u2.mem\[155\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11250__A1 _04248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06294_ u2.mem\[144\]\[2\] _01671_ _01673_ u2.mem\[182\]\[2\] _01799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_163_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08033_ _03491_ _03493_ _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_174_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07206__B1 _02683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10600__I1 u2.mem\[58\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09984_ _04698_ u2.mem\[43\]\[7\] _04745_ _04749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08935_ _04083_ _00313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_316_clock_I clknet_5_17_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11584__S _05738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08957__I _04096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08866_ _04014_ _04042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_170_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input21_I data_in_a[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06717__C1 _02200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07817_ _02531_ _03284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08797_ _03996_ _00262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_5_12_0_clock_I clknet_4_6_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09989__S _04750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11069__A1 _04394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07748_ u2.mem\[3\]\[11\] _03036_ _03215_ _03216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08893__S _04056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12635__CLK clknet_leaf_211_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07679_ _02595_ _03149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10928__S _05327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06496__A1 _01981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09418_ _04397_ _00482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08692__I _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10690_ _05110_ u2.mem\[60\]\[7\] _05179_ _05183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_16_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11616__I0 _05756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09349_ _04276_ u2.mem\[28\]\[11\] _04346_ _04350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_40_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08237__A2 _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12785__CLK clknet_leaf_336_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06248__A1 u2.mem\[184\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12360_ _00239_ clknet_leaf_137_clock u2.mem\[14\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07101__I _02579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06799__A2 _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11311_ _05556_ u2.mem\[156\]\[5\] _05567_ _05574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12291_ _00170_ clknet_leaf_110_clock u2.mem\[10\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06263__A4 _01768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12015__CLK clknet_2_3__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11919__I1 u2.mem\[193\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11242_ _05508_ u2.mem\[152\]\[2\] _05529_ _05532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_5_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08796__I0 _03913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11173_ _05466_ u2.mem\[148\]\[2\] _05484_ _05487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10124_ _04810_ u2.mem\[46\]\[12\] _04835_ _04836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06420__A1 u2.mem\[193\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06420__B2 u2.mem\[192\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10055_ _04791_ _00725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13410__CLK clknet_leaf_323_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_384_clock clknet_5_0_0_clock clknet_leaf_384_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_169_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_169_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_40_clock_I clknet_5_6_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13560__CLK clknet_leaf_32_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10957_ _05351_ _05352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11480__A1 _05354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10888_ _05004_ _05307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12627_ _00506_ clknet_leaf_111_clock u2.mem\[31\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07436__B1 _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12558_ _00437_ clknet_leaf_203_clock u2.mem\[27\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07011__I _02489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07987__A1 _03447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_322_clock clknet_5_16_0_clock clknet_leaf_322_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_265_clock_I clknet_5_22_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11509_ _04248_ _05690_ _05699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12489_ _00368_ clknet_leaf_125_clock u2.mem\[22\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09139__S _04218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08787__I0 _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11468__I _03501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07167__B _02359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08978__S _04107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_337_clock clknet_5_18_0_clock clknet_leaf_337_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_98_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06981_ _02439_ _02440_ _02458_ _02459_ _02460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_119_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13090__CLK clknet_leaf_256_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08720_ _03949_ _00232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11299__A1 _04333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12658__CLK clknet_leaf_235_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08651_ _03902_ _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07911__A1 u2.mem\[40\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07602_ u2.mem\[9\]\[8\] _03071_ _03072_ u2.mem\[25\]\[8\] _03073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07911__B2 u2.mem\[30\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08582_ _03807_ u2.mem\[11\]\[4\] _03861_ _03862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07533_ _03001_ _03002_ _03003_ _03004_ _03005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_23_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06478__A1 u2.mem\[193\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07675__B1 _03072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07464_ u2.mem\[15\]\[6\] _02794_ _02795_ u2.mem\[13\]\[6\] _02937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_62_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09401__I _04357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09203_ _04259_ _00405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06415_ _01912_ _01916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10547__I _05094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07395_ u2.mem\[32\]\[5\] _02786_ _02787_ u2.mem\[2\]\[5\] _02869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09267__I1 u2.mem\[26\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09134_ _04161_ u2.mem\[23\]\[10\] _04213_ _04216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12038__CLK clknet_leaf_316_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06346_ u2.mem\[178\]\[4\] _01746_ _01747_ u2.mem\[164\]\[4\] _01849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07427__B1 _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09967__A2 _04659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09065_ _04174_ u2.mem\[21\]\[14\] _04168_ _04175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06277_ u2.mem\[174\]\[2\] _01657_ _01659_ u2.mem\[155\]\[2\] _01661_ u2.mem\[181\]\[2\]
+ _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__10483__S _05056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07856__I _02616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08016_ mem_address_trans\[4\].data_sync _03477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_162_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06650__A1 u2.mem\[194\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12188__CLK clknet_leaf_267_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11378__I _05615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13433__CLK clknet_leaf_352_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09967_ _04311_ _04659_ _04739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08918_ _04073_ _04074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_135_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09898_ _04585_ _04696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07591__I _02536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08849_ _03687_ _04030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08950__I0 _04046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11860_ _05917_ _05918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11837__I0 _05876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10811_ u2.mem\[63\]\[4\] _03506_ _05258_ _05259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11791_ _05874_ u2.mem\[186\]\[4\] _05865_ _05875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08702__I0 _03938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11841__I _05904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06469__A1 u2.mem\[193\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13530_ _01409_ clknet_leaf_325_clock u2.mem\[191\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06469__B2 u2.mem\[194\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07666__B1 _03063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10742_ _05216_ u2.mem\[61\]\[9\] _05214_ _05217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13461_ _01340_ clknet_leaf_360_clock u2.mem\[180\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10673_ _04334_ _05172_ _05173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09258__I1 u2.mem\[26\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12412_ _00291_ clknet_leaf_192_clock u2.mem\[18\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13392_ _01271_ clknet_leaf_369_clock u2.mem\[168\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12343_ _00222_ clknet_leaf_139_clock u2.mem\[13\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12274_ _00153_ clknet_leaf_176_clock u2.mem\[9\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11225_ _05505_ u2.mem\[151\]\[1\] _05520_ _05522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09430__I1 u2.mem\[30\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11156_ _05464_ u2.mem\[147\]\[1\] _05475_ _05477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10107_ _04826_ _00742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10328__I0 _04913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11087_ _05433_ _01115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10038_ _04714_ u2.mem\[44\]\[14\] _04777_ _04780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08941__I0 _04037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12950__CLK clknet_leaf_63_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_3_0_0_clock_I clknet_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11989_ _00001_ clknet_leaf_335_clock u2.mem\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07657__B1 _03126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09221__I _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13306__CLK clknet_leaf_376_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07121__A2 _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09249__I1 u2.mem\[26\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06200_ _01556_ _01677_ _01593_ _01707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_07180_ u2.mem\[44\]\[1\] _02656_ _02657_ u2.mem\[42\]\[1\] _02658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_261_clock clknet_5_22_0_clock clknet_leaf_261_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06131_ u2.mem\[188\]\[0\] _01632_ _01634_ u2.mem\[187\]\[0\] _01637_ u2.mem\[192\]\[0\]
+ _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__12330__CLK clknet_leaf_136_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13456__CLK clknet_leaf_320_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07424__A3 _02888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06062_ _01558_ _01568_ _01569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11198__I _05501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_276_clock clknet_5_23_0_clock clknet_leaf_276_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_160_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09421__I1 u2.mem\[30\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10567__I0 _05108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12480__CLK clknet_leaf_176_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09821_ _04638_ _04649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_67_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06396__B1 _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09752_ _04607_ _00606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06964_ _02394_ _02443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__10319__I0 _04904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08703_ _03939_ _00225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08300__I _03658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06895_ _02373_ _02374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_09683_ _04487_ u2.mem\[36\]\[10\] _04554_ _04557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_66_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08932__I0 _04028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08634_ _03821_ u2.mem\[12\]\[10\] _03889_ _03892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_5_clock clknet_5_0_0_clock clknet_leaf_5_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_66_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_214_clock clknet_5_29_0_clock clknet_leaf_214_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11819__I0 _05872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08565_ _03828_ u2.mem\[10\]\[13\] _03850_ _03852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_78_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10478__S _05051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11661__I _05673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07648__B1 _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07516_ u2.mem\[58\]\[7\] _02811_ _02812_ u2.mem\[36\]\[7\] _02988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08496_ _03798_ _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_39_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08160__I1 u2.mem\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07447_ _02917_ _02918_ _02919_ _02920_ _02921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_161_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06320__B1 _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_229_clock clknet_5_19_0_clock clknet_leaf_229_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_7_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06871__A1 col_select_trans\[5\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07378_ _02605_ _02853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09117_ _04206_ _00372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06329_ _01830_ _01831_ _01832_ _01833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_136_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_8_clock_I clknet_5_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09048_ _04161_ u2.mem\[21\]\[10\] _04155_ _04162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12823__CLK clknet_leaf_129_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11010_ _05384_ u2.mem\[138\]\[1\] _05382_ _05385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06387__C2 u2.mem\[193\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_213_clock_I clknet_5_28_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12961_ _00840_ clknet_leaf_168_clock u2.mem\[52\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08923__I0 _04019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11912_ _01981_ _05929_ _05948_ _01425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07887__B1 _02555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12892_ _00771_ clknet_leaf_222_clock u2.mem\[48\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12203__CLK clknet_leaf_229_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13329__CLK clknet_leaf_1_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11843_ _05906_ _01398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07639__B1 _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11286__I1 u2.mem\[155\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11774_ _05837_ u2.mem\[185\]\[5\] _05856_ _05863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13513_ _01392_ clknet_leaf_354_clock u2.mem\[189\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11986__A2 _05972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10725_ _05195_ _05205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13479__CLK clknet_leaf_304_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06862__A1 col_select_trans\[5\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13444_ _01323_ clknet_leaf_364_clock u2.mem\[177\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10656_ _05163_ _00954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13375_ _01254_ clknet_leaf_367_clock u2.mem\[166\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10587_ _05121_ u2.mem\[57\]\[12\] _05122_ _05123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12326_ _00205_ clknet_leaf_93_clock u2.mem\[12\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12257_ _00136_ clknet_leaf_240_clock u2.mem\[8\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09417__S _04396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11208_ _05509_ _01160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12188_ _00067_ clknet_leaf_267_clock u2.mem\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06378__B1 _01658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06378__C2 u2.mem\[181\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11139_ _05465_ _01135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07590__A2 _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11682__S _05800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06680_ u2.mem\[169\]\[1\] _02142_ _02144_ u2.mem\[147\]\[1\] _02164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11481__I _05682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08350_ data_in_trans\[14\].data_sync _03716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11426__A1 _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07301_ _02773_ _02774_ _02775_ _02776_ _02777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_127_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08281_ _03660_ _00082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07232_ u2.mem\[50\]\[2\] _02647_ _02648_ u2.mem\[51\]\[2\] _02709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_4_4_0_clock_I clknet_3_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06853__A1 u2.mem\[146\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06853__B2 u2.mem\[186\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12846__CLK clknet_leaf_214_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07163_ _02635_ _02636_ _02637_ _02640_ _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06114_ _01571_ _01597_ _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06605__A1 u2.mem\[151\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_162_clock_I clknet_5_26_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07094_ _02446_ _02573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_12_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06605__B2 u2.mem\[158\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11857__S _05904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06045_ _01550_ _01551_ _01552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10761__S _05223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12996__CLK clknet_leaf_65_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09327__S _04336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06369__B1 _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09804_ _04565_ u2.mem\[39\]\[0\] _04639_ _04640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10560__I _05094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07030__B2 u2.mem\[20\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12226__CLK clknet_leaf_241_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07996_ _01614_ _03459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07581__A2 _03050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09735_ _04594_ _00602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08030__I _03490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06947_ _02425_ _02426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07869__B1 _02426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_153_clock clknet_5_24_0_clock clknet_leaf_153_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_27_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09666_ _04547_ _00580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06878_ _02347_ _02351_ _02356_ _02357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_08617_ _03882_ _00196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_5_22_0_clock clknet_4_11_0_clock clknet_5_22_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_76_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09597_ _04476_ u2.mem\[34\]\[5\] _04506_ _04508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11391__I _05499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_87_clock_I clknet_5_11_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08548_ _03842_ _00167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_168_clock clknet_5_26_0_clock clknet_leaf_168_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_24_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08479_ _03722_ u2.mem\[8\]\[15\] _03792_ _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10510_ _04987_ u2.mem\[56\]\[0\] _05073_ _05074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06844__A1 u2.mem\[144\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11490_ _05677_ u2.mem\[167\]\[4\] _05682_ _05688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06844__B2 u2.mem\[182\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08406__S _03753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10441_ _04998_ u2.mem\[54\]\[3\] _05030_ _05034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10372_ _04920_ u2.mem\[52\]\[15\] _04981_ _04985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08205__I _03607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13160_ _01039_ clknet_leaf_293_clock u2.mem\[130\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07939__A4 _03403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12111_ _01474_ clknet_leaf_348_clock u2.select_mem_row\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13001__CLK clknet_leaf_50_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13091_ _00970_ clknet_leaf_26_clock u2.mem\[60\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12042_ col_select_trans\[2\].A clknet_leaf_315_clock col_select_trans\[2\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_106_clock clknet_5_11_0_clock clknet_leaf_106_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07021__A1 _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07572__A2 _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13151__CLK clknet_leaf_260_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_364_clock_I clknet_5_4_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12719__CLK clknet_leaf_250_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08875__I _03721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12944_ _00823_ clknet_leaf_151_clock u2.mem\[51\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12875_ _00754_ clknet_leaf_228_clock u2.mem\[47\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06678__A4 _02162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11007__S _05382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11826_ _05895_ _05896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09700__S _04567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11757_ _05853_ _01365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07627__A3 _03088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06835__A1 u2.mem\[187\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10708_ _05128_ u2.mem\[60\]\[15\] _05189_ _05193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06835__B2 u2.mem\[192\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11688_ _05811_ _01338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13427_ _01306_ clknet_leaf_365_clock u2.mem\[174\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10645__I _05151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10639_ _05097_ u2.mem\[59\]\[1\] _05152_ _05154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08115__I _03545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13358_ _01237_ clknet_leaf_372_clock u2.mem\[163\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12309_ _00188_ clknet_leaf_98_clock u2.mem\[11\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13289_ _01168_ clknet_leaf_0_clock u2.mem\[151\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12249__CLK clknet_leaf_55_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11476__I _03509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07012__A1 u2.mem\[58\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10380__I _04126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07850_ u2.mem\[52\]\[12\] _03315_ _03316_ u2.mem\[21\]\[12\] _03317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10942__I0 _05340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_70_clock clknet_5_8_0_clock clknet_leaf_70_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_56_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06801_ u2.mem\[171\]\[4\] _02066_ _02068_ u2.mem\[157\]\[4\] _02281_ _02282_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_68_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07781_ _03233_ _03238_ _03243_ _03248_ _03249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12399__CLK clknet_leaf_172_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput3 col_select_a[2] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09520_ _04382_ u2.mem\[32\]\[11\] _04453_ _04457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06732_ u2.mem\[187\]\[2\] _02186_ _02187_ u2.mem\[192\]\[2\] _02215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_leaf_109_clock_I clknet_5_11_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09560__I0 _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09451_ _04415_ _00497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06663_ _02147_ _02148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_85_clock clknet_5_9_0_clock clknet_leaf_85_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_51_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08402_ _03747_ _03749_ _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09382_ _04371_ u2.mem\[29\]\[6\] _04367_ _04372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06594_ _02078_ _02079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07079__A1 _02522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09610__S _04511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08333_ _03702_ _00092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06826__A1 u2.mem\[164\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08264_ _03648_ _00077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08226__S _03623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07215_ u2.mem\[8\]\[1\] _02610_ _02612_ u2.mem\[4\]\[1\] _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08195_ _03480_ _03605_ _03482_ _03606_ _03607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__13024__CLK clknet_leaf_265_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07146_ u2.mem\[6\]\[0\] _02622_ _02624_ u2.mem\[47\]\[0\] _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_173_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_5_8_0_clock_I clknet_4_4_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_23_clock clknet_5_2_0_clock clknet_leaf_23_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_145_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07077_ u2.mem\[61\]\[0\] _02553_ _02555_ u2.mem\[63\]\[0\] _02556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_156_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09379__I0 _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09057__S _04168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13174__CLK clknet_leaf_279_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06028_ u2.driver_mem\[13\] _01517_ _01537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_134_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07003__A1 _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10290__I _04922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_38_clock clknet_5_6_0_clock clknet_leaf_38_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_130_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07554__A2 _02871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07979_ u2.mem\[29\]\[15\] _03301_ _03302_ u2.mem\[11\]\[15\] _03443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06762__B1 _02099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09718_ _04581_ _00598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08695__I _03713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10990_ _04249_ _05363_ _05372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_55_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09649_ _04521_ _04537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_76_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12660_ _00539_ clknet_leaf_83_clock u2.mem\[33\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09520__S _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11611_ _05763_ _01309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_169_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12591_ _00470_ clknet_leaf_181_clock u2.mem\[29\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11542_ _05720_ _01283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06293__A2 _01699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11473_ _05676_ _05677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_13_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13212_ _01091_ clknet_leaf_290_clock u2.mem\[138\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_167_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10424_ _03712_ _05023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11413__I1 u2.mem\[163\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13517__CLK clknet_leaf_325_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11497__S _05692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08290__I0 _03667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13143_ _01022_ clknet_leaf_40_clock u2.mem\[63\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10355_ _04975_ _00841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10286_ _04909_ u2.mem\[50\]\[10\] _04933_ _04936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13074_ _00953_ clknet_leaf_249_clock u2.mem\[59\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11177__I0 _05470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12541__CLK clknet_leaf_198_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12025_ net37 clknet_2_3__leaf_clock_a row_select_trans\[0\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10924__I0 _05299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_110_clock_I clknet_5_11_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12927_ _00806_ clknet_leaf_242_clock u2.mem\[50\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11960__S _05975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06339__B _01842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12858_ _00737_ clknet_leaf_143_clock u2.mem\[45\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07014__I _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11809_ _05885_ _01385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13047__CLK clknet_leaf_340_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12789_ _00668_ clknet_leaf_28_clock u2.mem\[41\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06808__A1 u2.mem\[155\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06808__B2 u2.mem\[150\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10375__I _04986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07000_ _02478_ _02479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__12071__CLK clknet_2_0__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13197__CLK clknet_leaf_294_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_35_clock_I clknet_5_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07784__A2 _03099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08951_ _04092_ _00320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07902_ u2.mem\[5\]\[13\] _02627_ _02629_ u2.mem\[38\]\[13\] _03368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08882_ _04017_ u2.mem\[18\]\[1\] _04051_ _04053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07833_ u2.mem\[26\]\[12\] _03141_ _03142_ u2.mem\[10\]\[12\] _03300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07764_ u2.mem\[57\]\[11\] _03137_ _03138_ u2.mem\[41\]\[11\] _03232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_84_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09404__I _04170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09503_ _04447_ _00517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06715_ _02134_ _02199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07695_ _01958_ _03017_ _03131_ _03164_ _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09434_ _04395_ _04406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_169_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06646_ _02130_ _02131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09365_ _04127_ _04360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06577_ _02061_ _02062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07859__I _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08316_ _03688_ u2.mem\[5\]\[7\] _03676_ _03689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_312_clock_I clknet_5_17_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12414__CLK clknet_leaf_191_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09296_ _04319_ _00438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07472__A1 u2.mem\[58\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08247_ _03633_ _03639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06275__A2 _01776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08178_ _03566_ u2.mem\[2\]\[9\] _03595_ _03597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07224__A1 u2.mem\[40\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07129_ _02592_ _02597_ _02602_ _02607_ _02608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__12564__CLK clknet_leaf_90_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07224__B2 u2.mem\[30\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08272__I0 _03579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11110__S _05445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10140_ _04790_ u2.mem\[47\]\[3\] _04841_ _04845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06983__B1 _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10071_ _04801_ u2.mem\[45\]\[8\] _04802_ _04803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11859__A1 _04416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07527__A2 _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06003__I _01511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11844__I _03661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08327__I1 u2.mem\[5\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10973_ _05352_ u2.mem\[135\]\[5\] _05355_ _05362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12712_ _00591_ clknet_leaf_146_clock u2.mem\[36\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12643_ _00522_ clknet_leaf_93_clock u2.mem\[32\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12094__CLK clknet_leaf_337_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06673__I _02157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12574_ _00453_ clknet_leaf_200_clock u2.mem\[28\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11634__I1 u2.mem\[176\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10598__A1 _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07463__A1 _02932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11525_ _05708_ _05709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_11_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06266__A2 _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12907__CLK clknet_leaf_207_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11456_ _04179_ _05645_ _05664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10407_ _03690_ _05011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08263__I0 _03570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11387_ _05593_ u2.mem\[161\]\[4\] _05615_ _05621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07766__A2 _03141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13126_ _01005_ clknet_leaf_21_clock u2.mem\[62\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10338_ _04965_ _04966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_113_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06974__B1 _02452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11955__S _05972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13057_ _00936_ clknet_leaf_256_clock u2.mem\[58\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10269_ _04926_ _00804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07518__A2 _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12008_ mem_address_trans\[1\].A clknet_leaf_315_clock mem_address_trans\[1\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09763__I0 _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11570__I0 _05719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_261_clock_I clknet_5_22_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09224__I _04160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06500_ _01984_ _01985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07480_ u2.mem\[61\]\[6\] _02899_ _02900_ u2.mem\[63\]\[6\] _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_62_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12437__CLK clknet_leaf_102_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07151__B1 _02629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06431_ _01727_ _01915_ _01926_ _01930_ _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_61_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07679__I _02595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09150_ _04225_ _04226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06362_ u2.mem\[152\]\[4\] _01713_ _01715_ u2.mem\[148\]\[4\] _01865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_163_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08101_ _03482_ _03541_ _03544_ _03545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_09081_ _04136_ u2.mem\[22\]\[3\] _04182_ _04186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12587__CLK clknet_leaf_205_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06293_ u2.mem\[154\]\[2\] _01699_ _01701_ u2.mem\[162\]\[2\] _01797_ _01798_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_174_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08032_ _03492_ _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11389__I0 _05595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06009__A2 _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08254__I0 _03561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07757__A2 _03050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10061__I0 _04795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08303__I _03509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09983_ _04748_ _00696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11865__S _05918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08934_ _04030_ u2.mem\[19\]\[7\] _04079_ _04083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08865_ _03708_ _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06717__C2 u2.mem\[160\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07816_ _02527_ _03283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08796_ _03913_ u2.mem\[16\]\[4\] _03995_ _03996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06193__A1 _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input14_I data_in_a[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07747_ _02357_ _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07678_ _02593_ _03148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_5_16_0_clock_I clknet_4_8_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09417_ _04356_ u2.mem\[30\]\[0\] _04396_ _04397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06629_ _02045_ _02001_ _02114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06496__A2 _01927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07589__I _02543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09348_ _04349_ _00460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11616__I1 u2.mem\[175\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08237__A3 _03632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06248__A2 _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07445__A1 u2.mem\[52\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08493__I0 _03805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09279_ _04308_ _00432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11310_ _05573_ _01198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12290_ _00169_ clknet_leaf_179_clock u2.mem\[10\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11839__I _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08245__I0 _03552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11241_ _05531_ _01171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07748__A2 _03036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09993__I0 _04707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11172_ _05486_ _01147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10123_ _04819_ _04835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_121_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10054_ _04790_ u2.mem\[45\]\[3\] _04784_ _04791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_121_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06668__I _02152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06184__A1 _01566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07381__B1 _02690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07920__A2 _02499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10956_ _04143_ _05351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11480__A2 _05645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10887_ _05306_ _01042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12626_ _00505_ clknet_leaf_180_clock u2.mem\[31\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07436__A1 u2.mem\[26\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08484__I0 _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12557_ _00436_ clknet_leaf_202_clock u2.mem\[27\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_208_clock_I clknet_5_30_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10291__I0 _04913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11508_ _05698_ _01271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12488_ _00367_ clknet_leaf_125_clock u2.mem\[22\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11749__I _05848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11439_ _05653_ _01247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07739__A2 _03099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09984__I0 _04698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11791__I0 _05874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13235__CLK clknet_leaf_288_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13109_ _00988_ clknet_leaf_21_clock u2.mem\[61\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06980_ _02394_ _02459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09155__S _04226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input6_I col_select_a[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09361__A1 _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08650_ _03900_ _03901_ _03902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_94_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07601_ _02576_ _03072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13385__CLK clknet_leaf_323_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08581_ _03855_ _03861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_78_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07532_ u2.mem\[28\]\[7\] _02841_ _02842_ u2.mem\[31\]\[7\] _03004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07463_ _02932_ _02933_ _02934_ _02935_ _02936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_39_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06478__A2 _01960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10828__I _05252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07675__B2 u2.mem\[25\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09202_ _04258_ u2.mem\[25\]\[3\] _04252_ _04259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06414_ _01914_ _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07394_ u2.mem\[45\]\[5\] _02866_ _02867_ u2.mem\[34\]\[5\] _02868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_33_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09133_ _04215_ _00379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07427__A1 u2.mem\[61\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08475__I0 _03714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06345_ _01845_ _01846_ _01847_ _01848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_163_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07978__A2 _02567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10282__I0 _04904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09064_ _04173_ _04174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06276_ u2.mem\[189\]\[2\] _01650_ _01663_ u2.mem\[180\]\[2\] _01652_ u2.mem\[176\]\[2\]
+ _01781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_135_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08015_ u3.data _03476_ net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06650__A2 _02133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10563__I _05004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09129__I _04202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10034__I0 _04709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09975__I0 _04689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11782__I0 _05868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06402__A2 _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09966_ _04738_ _00689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09065__S _04168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12602__CLK clknet_leaf_116_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08917_ _04072_ _03988_ _04073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09897_ _04695_ _00663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08848_ _04029_ _00280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07902__A2 _02627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08779_ mem_address_trans\[4\].data_sync _03983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA_clkbuf_leaf_4_clock_I clknet_5_0_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_157_clock_I clknet_5_25_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12752__CLK clknet_leaf_247_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10810_ _05252_ _05258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_2858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11837__I1 u2.mem\[189\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11790_ _03673_ _05874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06469__A2 _01960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10738__I _05195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10741_ _03695_ _05216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13460_ _01339_ clknet_leaf_360_clock u2.mem\[180\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10672_ _04862_ _05172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07112__I _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12411_ _00290_ clknet_leaf_190_clock u2.mem\[18\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08466__I0 _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13391_ _01270_ clknet_leaf_367_clock u2.mem\[168\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10273__I0 _04895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12342_ _00221_ clknet_leaf_92_clock u2.mem\[13\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07433__A4 _02906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13258__CLK clknet_leaf_285_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12273_ _00152_ clknet_leaf_176_clock u2.mem\[9\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06641__A2 _02125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09039__I _04123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10025__I0 _04700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_17_0_clock clknet_4_8_0_clock clknet_5_17_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_88_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11224_ _05521_ _01164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11155_ _05476_ _01140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10106_ _04792_ u2.mem\[46\]\[4\] _04825_ _04826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11086_ _05432_ u2.mem\[142\]\[5\] _05421_ _05433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10037_ _04779_ _00719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10849__S _05278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11988_ _00000_ clknet_leaf_380_clock u3.data vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10939_ _05338_ _01062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_3_4_0_clock_I clknet_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08118__I _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07022__I _02500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12609_ _00488_ clknet_leaf_155_clock u2.mem\[30\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08457__I0 _03680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_359_clock_I clknet_5_5_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10264__I0 _04885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06130_ _01636_ _01637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07424__A4 _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06061_ col_select_trans\[3\].data_sync _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10016__I0 _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11764__I0 _05825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09820_ _04648_ _00633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07593__B1 _03063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09751_ _04605_ u2.mem\[37\]\[12\] _04606_ _04607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06963_ _02441_ _02429_ _02416_ _02442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_171_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08702_ _03938_ u2.mem\[13\]\[15\] _03932_ _03939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12775__CLK clknet_leaf_141_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09682_ _04556_ _00587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06148__A1 u2.mem\[189\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06894_ _02372_ _02373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06148__B2 u2.mem\[176\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09613__S _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08633_ _03891_ _00203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07896__A1 _03358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07641__B _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08564_ _03851_ _00174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12005__CLK clknet_2_0__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11819__I1 u2.mem\[188\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07515_ u2.mem\[53\]\[7\] _02808_ _02809_ u2.mem\[56\]\[7\] _02987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08696__I0 _03934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08495_ _03674_ _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07446_ u2.mem\[18\]\[5\] _02852_ _02853_ u2.mem\[19\]\[5\] _02920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_126_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08028__I _03488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06320__A1 u2.mem\[187\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06320__B2 u2.mem\[192\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12155__CLK clknet_leaf_231_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10494__S _05061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08448__I0 _03663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07377_ _02603_ _02852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09116_ _04132_ u2.mem\[23\]\[2\] _04203_ _04206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06328_ u2.mem\[152\]\[3\] _01712_ _01714_ u2.mem\[148\]\[3\] _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08073__A1 _01962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09047_ _04160_ _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06623__A2 _02104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_383_clock clknet_5_0_0_clock clknet_leaf_383_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06259_ u2.mem\[152\]\[1\] _01713_ _01708_ u2.mem\[153\]\[1\] _01765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_159_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10007__I0 _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_83_clock_I clknet_5_9_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13550__CLK clknet_leaf_8_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08698__I _03717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06387__A1 u2.mem\[158\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07584__B1 _03054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06387__B2 u2.mem\[151\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09949_ _04718_ _04729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_89_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11507__I0 _05680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12960_ _00839_ clknet_leaf_168_clock u2.mem\[52\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07107__I _02585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09523__S _04458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11911_ _03534_ _05929_ _05948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12891_ _00770_ clknet_leaf_224_clock u2.mem\[48\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_321_clock clknet_5_16_0_clock clknet_leaf_321_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_72_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07887__B2 u2.mem\[63\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11842_ _05903_ u2.mem\[190\]\[0\] _05905_ _05906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09322__I _04333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11773_ _05862_ _01372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10494__I0 _05016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13512_ _01391_ clknet_leaf_354_clock u2.mem\[188\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10724_ _05000_ _05204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06311__A1 u2.mem\[155\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_336_clock clknet_5_18_0_clock clknet_leaf_336_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08439__I0 _03722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13443_ _01322_ clknet_leaf_363_clock u2.mem\[177\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10655_ _05112_ u2.mem\[59\]\[8\] _05162_ _05163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_360_clock_I clknet_5_5_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12648__CLK clknet_leaf_114_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13374_ _01253_ clknet_leaf_369_clock u2.mem\[165\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10586_ _05094_ _05122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_154_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12325_ _00204_ clknet_leaf_91_clock u2.mem\[12\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12256_ _00135_ clknet_leaf_229_clock u2.mem\[8\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08602__S _03871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11207_ _05508_ u2.mem\[150\]\[2\] _05502_ _05509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12798__CLK clknet_leaf_208_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12187_ _00066_ clknet_leaf_266_clock u2.mem\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07575__B1 _03045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06378__B2 u2.mem\[155\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_11_0_clock_I clknet_3_5_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11138_ _05464_ u2.mem\[146\]\[1\] _05462_ _05465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12070__D data_in_trans\[10\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12028__CLK clknet_leaf_304_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11069_ _04394_ _05402_ _05421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_76_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12178__CLK clknet_leaf_239_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11426__A2 _05645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07300_ u2.mem\[18\]\[3\] _02604_ _02606_ u2.mem\[19\]\[3\] _02776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__13423__CLK clknet_leaf_361_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10485__I0 _05007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08280_ _03656_ u2.mem\[5\]\[0\] _03659_ _03660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06302__A1 _01780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07231_ _02704_ _02705_ _02706_ _02707_ _02708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06853__A2 _02155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11203__S _05502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06591__I _02075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07162_ u2.mem\[27\]\[1\] _02638_ _02639_ u2.mem\[35\]\[1\] _02640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08055__A1 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13573__CLK clknet_leaf_16_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_105_clock_I clknet_5_11_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06113_ u2.mem\[178\]\[0\] _01617_ _01619_ u2.mem\[164\]\[0\] _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_172_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07093_ _02571_ _02572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_4_8_0_clock_I clknet_3_4_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08850__I0 _04030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09608__S _04511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06044_ col_select_trans\[4\].data_sync _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_160_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11737__I0 _05829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08602__I0 _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06369__A1 u2.mem\[146\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06369__B2 u2.mem\[186\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09407__I _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09803_ _04638_ _04639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07030__A2 _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06032__S _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07995_ _01562_ _01575_ _03458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09734_ _04592_ u2.mem\[37\]\[8\] _04593_ _04594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06946_ _02421_ _02422_ _02423_ _02424_ _02425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_39_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09343__S _04346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07869__A1 u2.mem\[27\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09665_ _04469_ u2.mem\[36\]\[2\] _04544_ _04547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06877_ _02352_ _02353_ _02355_ _02356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_08616_ _03803_ u2.mem\[12\]\[2\] _03879_ _03882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09596_ _04507_ _00550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08547_ _03810_ u2.mem\[10\]\[5\] _03840_ _03842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_93_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10476__I0 _04995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08478_ _03795_ _00144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07429_ u2.mem\[37\]\[5\] _02829_ _02830_ u2.mem\[59\]\[5\] _02903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06844__A2 _02114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07597__I _02558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10228__I0 _04898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08046__A1 _01809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10440_ _05033_ _00868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11976__I0 _05218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08841__I0 _04023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10371_ _04984_ _00848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12940__CLK clknet_leaf_221_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12110_ _05992_ clknet_leaf_381_clock u2.driver_enable vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09518__S _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13090_ _00969_ clknet_leaf_256_clock u2.mem\[60\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11728__I0 _05835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11847__I _03665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12041_ net3 clknet_2_2__leaf_clock_a col_select_trans\[2\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10751__I _05195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_307_clock_I clknet_5_20_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06780__A1 u2.mem\[155\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_260_clock clknet_5_22_0_clock clknet_leaf_260_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09253__S _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12943_ _00822_ clknet_leaf_242_clock u2.mem\[51\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10399__S _05002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12320__CLK clknet_leaf_167_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13446__CLK clknet_leaf_352_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12874_ _00753_ clknet_leaf_133_clock u2.mem\[46\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11825_ _05411_ _05886_ _05895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_275_clock clknet_5_23_0_clock clknet_leaf_275_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11756_ _05833_ u2.mem\[184\]\[3\] _05849_ _05853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12470__CLK clknet_leaf_103_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08824__A3 _03544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10707_ _05192_ _00976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06835__A2 _02100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11687_ _05786_ u2.mem\[180\]\[0\] _05810_ _05811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_174_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13426_ _01305_ clknet_leaf_365_clock u2.mem\[174\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08037__A1 _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10638_ _05153_ _00946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11967__I0 _05209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11958__S _05975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13357_ _01236_ clknet_leaf_373_clock u2.mem\[163\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10862__S _05287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10569_ _03686_ _05110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_4_clock clknet_5_0_0_clock clknet_leaf_4_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12308_ _00187_ clknet_leaf_96_clock u2.mem\[11\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07260__A2 _02610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08332__S _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13288_ _01167_ clknet_leaf_383_clock u2.mem\[151\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_213_clock clknet_5_28_0_clock clknet_leaf_213_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11719__I0 _05829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12239_ _00118_ clknet_leaf_239_clock u2.mem\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09227__I _04163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07012__A2 _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08131__I _03520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11693__S _05810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06800_ _02278_ _02279_ _02280_ _02281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xclkbuf_leaf_228_clock clknet_5_28_0_clock clknet_leaf_228_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07780_ _03244_ _03245_ _03246_ _03247_ _03248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_84_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06771__A1 u2.mem\[171\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06771__B2 u2.mem\[157\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput4 col_select_a[3] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_06731_ _02210_ _02211_ _02212_ _02213_ _02214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_76_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09450_ _04391_ u2.mem\[30\]\[15\] _04411_ _04415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_25_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06662_ _02044_ _02011_ _02147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07720__B1 _03138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_31_clock_I clknet_5_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08401_ _03748_ _03631_ _03749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12813__CLK clknet_leaf_206_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09381_ _04147_ _04371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06593_ _02006_ _02077_ _02078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_127_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08332_ _03701_ u2.mem\[5\]\[10\] _03693_ _03702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06287__B1 _01734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08263_ _03570_ u2.mem\[4\]\[11\] _03644_ _03648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12963__CLK clknet_leaf_110_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07214_ u2.mem\[39\]\[1\] _02617_ _02619_ u2.mem\[48\]\[1\] _02692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08194_ _03540_ _03606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_146_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11958__I0 _05909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07145_ _02623_ _02624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_256_clock_I clknet_5_19_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07251__A2 _02580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07076_ _02554_ _02555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06027_ u2.driver_mem\[14\] _01522_ _01535_ _01536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_161_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07539__B1 _02923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13469__CLK clknet_leaf_360_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07978_ u2.mem\[26\]\[15\] _02567_ _02569_ u2.mem\[10\]\[15\] _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_74_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06762__B2 u2.mem\[161\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09717_ _04579_ u2.mem\[37\]\[4\] _04580_ _04581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06929_ _02407_ _02408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_28_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11108__S _05445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10697__I0 _05117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09648_ _04536_ _00573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12493__CLK clknet_leaf_197_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07711__B1 _03123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09579_ _04496_ u2.mem\[33\]\[14\] _04492_ _04497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11610_ _05750_ u2.mem\[175\]\[1\] _05761_ _05763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12590_ _00469_ clknet_leaf_201_clock u2.mem\[29\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11110__I1 u2.mem\[144\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06278__B1 _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11541_ _05719_ u2.mem\[170\]\[5\] _05708_ _05720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06817__A2 _02129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11472_ _03505_ _05676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07490__A2 _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07120__I _02598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13211_ _01090_ clknet_leaf_301_clock u2.mem\[138\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10423_ _05022_ _00862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13142_ _01021_ clknet_leaf_19_clock u2.mem\[63\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10354_ _04902_ u2.mem\[52\]\[7\] _04971_ _04975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07242__A2 _02708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13073_ _00952_ clknet_leaf_335_clock u2.mem\[59\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10285_ _04935_ _00811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09047__I _04160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12024_ mem_address_trans\[9\].A clknet_leaf_321_clock mem_address_trans\[9\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_152_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12836__CLK clknet_leaf_88_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10688__I0 _05108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12926_ _00805_ clknet_leaf_221_clock u2.mem\[50\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07702__B1 _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12857_ _00736_ clknet_5_13_0_clock u2.mem\[45\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12986__CLK clknet_leaf_50_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11808_ _05876_ u2.mem\[187\]\[5\] _05878_ _05885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08327__S _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12788_ _00667_ clknet_leaf_28_clock u2.mem\[41\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11739_ _05831_ u2.mem\[183\]\[2\] _05840_ _05843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12216__CLK clknet_leaf_54_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10860__I0 _05198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08805__I0 _03922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13409_ _01288_ clknet_leaf_319_clock u2.mem\[171\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07769__B1 _03075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_152_clock clknet_5_24_0_clock clknet_leaf_152_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_157_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07233__A2 _02650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12366__CLK clknet_leaf_209_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08950_ _04046_ u2.mem\[19\]\[14\] _04089_ _04092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07901_ _03363_ _03364_ _03365_ _03366_ _03367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_44_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08881_ _04052_ _00290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_167_clock clknet_5_26_0_clock clknet_leaf_167_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_116_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09930__A1 _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07832_ _03291_ _03294_ _03297_ _03298_ _03299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_170_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06744__A1 u2.mem\[194\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07763_ u2.mem\[37\]\[11\] _03062_ _03063_ u2.mem\[59\]\[11\] _03231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09502_ _04364_ u2.mem\[32\]\[3\] _04443_ _04447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06714_ _02133_ _02198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10679__I0 _05099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07694_ _03140_ _03147_ _03154_ _03163_ _03164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07205__I _02595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09433_ _04405_ _00489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06645_ _02107_ _02070_ _02130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10767__S _05232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09364_ _04359_ _00466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09297__I0 _04263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06576_ _02057_ _02060_ _02061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_105_clock clknet_5_11_0_clock clknet_leaf_105_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_90_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08315_ _03687_ _03688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10566__I _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09295_ _04260_ u2.mem\[27\]\[4\] _04318_ _04319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10851__I0 _05204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08246_ _03638_ _00069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08036__I _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13141__CLK clknet_leaf_20_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08177_ _03596_ _00042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12709__CLK clknet_leaf_64_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07128_ u2.mem\[18\]\[0\] _02604_ _02606_ u2.mem\[19\]\[0\] _02607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07224__A2 _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08272__I1 u2.mem\[4\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10007__S _04762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07059_ _02463_ _02515_ _02516_ _02417_ _02538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12859__CLK clknet_leaf_211_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10070_ _04783_ _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_138_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06735__A1 _02215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10972_ _05361_ _01072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07115__I _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12711_ _00590_ clknet_leaf_142_clock u2.mem\[36\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10677__S _05174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12642_ _00521_ clknet_leaf_159_clock u2.mem\[32\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09288__I0 _04254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12239__CLK clknet_leaf_239_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12573_ _00452_ clknet_leaf_201_clock u2.mem\[28\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11524_ _04287_ _05690_ _05708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12389__CLK clknet_leaf_79_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11455_ _05662_ _05663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_171_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07785__I _02384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10406_ _05010_ _00857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07215__A2 _02610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09460__I0 _04362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11386_ _05620_ _01227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08263__I1 u2.mem\[4\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13125_ _01004_ clknet_leaf_21_clock u2.mem\[62\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_84_clock clknet_5_9_0_clock clknet_leaf_84_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10337_ _04095_ _04964_ _04965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13056_ _00935_ clknet_leaf_256_clock u2.mem\[58\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09212__I0 _04265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10268_ _04891_ u2.mem\[50\]\[2\] _04923_ _04926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12007_ net25 clknet_2_1__leaf_clock_a mem_address_trans\[1\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10199_ _04879_ _00781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06726__A1 _02205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_99_clock clknet_5_10_0_clock clknet_leaf_99_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11570__I1 u2.mem\[172\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_204_clock_I clknet_5_31_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11971__S _05980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09441__S _04406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12909_ _00788_ clknet_leaf_202_clock u2.mem\[49\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_22_clock clknet_5_2_0_clock clknet_leaf_22_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_146_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06430_ u2.mem\[193\]\[1\] _01928_ _01929_ u2.mem\[192\]\[1\] _01914_ _01930_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_34_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09240__I _04176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13164__CLK clknet_leaf_285_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11086__I0 _05432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06361_ u2.mem\[153\]\[4\] _01708_ _01710_ u2.mem\[160\]\[4\] _01864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_33_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08100_ _03542_ _03543_ _03544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_147_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_37_clock clknet_5_6_0_clock clknet_leaf_37_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09080_ _04185_ _00356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06292_ _01794_ _01795_ _01796_ _01797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_124_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_147_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08031_ _03487_ _03492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput40 row_select_a[3] net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_159_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11211__S _05502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11389__I1 u2.mem\[161\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07206__A2 _02682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10210__A1 _04013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09982_ _04696_ u2.mem\[43\]\[6\] _04745_ _04748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06965__A1 _02439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08933_ _04082_ _00312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06104__I _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11010__I0 _05384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08864_ _04040_ _00285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06717__A1 u2.mem\[194\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07815_ u2.mem\[14\]\[12\] _03125_ _03126_ u2.mem\[12\]\[12\] _03282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_123_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08795_ _03989_ _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07390__A1 _02833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06193__A2 _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07746_ u2.mem\[16\]\[11\] _03033_ _03034_ u2.mem\[33\]\[11\] _03214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07677_ _03143_ _03144_ _03145_ _03146_ _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_129_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09416_ _04395_ _04396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_77_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06628_ _02083_ _02090_ _02095_ _02112_ _02113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_90_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09150__I _04225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09347_ _04274_ u2.mem\[28\]\[10\] _04346_ _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06559_ _02022_ _02044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12531__CLK clknet_leaf_111_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11777__A1 _04287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09278_ _04283_ u2.mem\[26\]\[14\] _04305_ _04308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09690__I0 _04494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08229_ _03626_ _00064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06653__B1 _02137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_0_clock_I clknet_5_0_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11240_ _05505_ u2.mem\[152\]\[1\] _05529_ _05531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_153_clock_I clknet_5_24_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11171_ _05464_ u2.mem\[148\]\[1\] _05484_ _05486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06956__A1 _02421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10122_ _04834_ _00749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13037__CLK clknet_leaf_282_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10053_ _04575_ _04790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07905__B1 _02624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06184__A2 _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11791__S _05865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12061__CLK clknet_2_1__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13187__CLK clknet_leaf_292_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_13_0_clock clknet_4_6_0_clock clknet_5_13_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_17_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10955_ _05350_ _01066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_78_clock_I clknet_5_8_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10886_ _05305_ u2.mem\[130\]\[4\] _05296_ _05306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09060__I _04170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12625_ _00504_ clknet_leaf_181_clock u2.mem\[31\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09995__I _04739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07436__A2 _02908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12556_ _00435_ clknet_leaf_202_clock u2.mem\[27\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09681__I0 _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11507_ _05680_ u2.mem\[168\]\[5\] _05691_ _05698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07987__A3 _03449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10934__I _04117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12487_ _00366_ clknet_leaf_125_clock u2.mem\[22\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05998__A2 row_col_select_trans.data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11438_ _05635_ u2.mem\[164\]\[5\] _05646_ _05653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_172_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11240__I0 _05505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11369_ _05589_ u2.mem\[160\]\[2\] _05608_ _05611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11791__I1 u2.mem\[186\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13108_ _00987_ clknet_leaf_17_clock u2.mem\[61\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13039_ _00918_ clknet_leaf_335_clock u2.mem\[57\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12404__CLK clknet_leaf_103_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07600_ _02571_ _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08580_ _03860_ _00181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09171__S _04236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07531_ u2.mem\[9\]\[7\] _02838_ _02839_ u2.mem\[25\]\[7\] _03003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_19_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07124__A1 _02522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12554__CLK clknet_leaf_123_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07462_ u2.mem\[27\]\[6\] _02871_ _02872_ u2.mem\[35\]\[6\] _02935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06594__I _02078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07675__A2 _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09201_ _04135_ _04258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06413_ _01913_ _01914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07393_ _02435_ _02867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09132_ _04158_ u2.mem\[23\]\[9\] _04213_ _04215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10806__I0 u2.mem\[63\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06344_ u2.mem\[172\]\[4\] _01654_ _01667_ u2.mem\[150\]\[4\] _01847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_31_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07427__A2 _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09672__I0 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09063_ data_in_trans\[14\].data_sync _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06275_ _01775_ _01776_ _01777_ _01779_ _01780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_8_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08014_ u3.enable _03476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08314__I _03686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10780__S _05237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06938__A1 _02390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11782__I1 u2.mem\[186\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09965_ _04716_ u2.mem\[42\]\[15\] _04734_ _04738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08916_ _04071_ _04072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_4206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12084__CLK clknet_leaf_381_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09896_ _04694_ u2.mem\[41\]\[5\] _04692_ _04695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_4217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08847_ _04028_ u2.mem\[17\]\[6\] _04024_ _04029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08984__I _04096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08778_ _03485_ _03982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09081__S _04182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07729_ u2.mem\[52\]\[10\] _03082_ _03083_ u2.mem\[21\]\[10\] _03198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11116__S _05444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10020__S _04767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10740_ _05215_ _00986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07666__A2 _03062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_31_0_clock_I clknet_4_15_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10671_ _05171_ _00961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12410_ _00289_ clknet_leaf_124_clock u2.mem\[17\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13390_ _01269_ clknet_leaf_364_clock u2.mem\[168\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09663__I0 _04467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12341_ _00220_ clknet_leaf_94_clock u2.mem\[13\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11470__I0 _05674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10754__I _03712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12272_ _00151_ clknet_leaf_179_clock u2.mem\[9\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11223_ _05500_ u2.mem\[151\]\[0\] _05520_ _05521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10690__S _05179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12427__CLK clknet_leaf_190_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08160__S _03585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11154_ _05460_ u2.mem\[147\]\[0\] _05475_ _05476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10105_ _04819_ _04825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_122_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11085_ _05351_ _05432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09055__I _04166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10036_ _04712_ u2.mem\[44\]\[13\] _04777_ _04779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11987_ _01979_ _05972_ _05991_ _01457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11026__S _05395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07657__A2 _03125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10938_ _05335_ u2.mem\[134\]\[0\] _05337_ _05338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12068__D data_in_trans\[9\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10869_ _05293_ _01037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12608_ _00487_ clknet_leaf_157_clock u2.mem\[30\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09654__I0 _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10264__I1 u2.mem\[50\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12539_ _00418_ clknet_leaf_187_clock u2.mem\[26\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13202__CLK clknet_leaf_297_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06060_ _01566_ _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08134__I _03522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07290__B1 _02672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11913__A1 _04013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11764__I1 u2.mem\[185\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13352__CLK clknet_leaf_377_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06396__A2 _01707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06962_ _02404_ _02441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_09750_ _04566_ _04606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_171_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08701_ _03721_ _03938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09681_ _04485_ u2.mem\[36\]\[9\] _04554_ _04556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06893_ _02364_ _02371_ _02353_ _02372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_66_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08393__I0 _03714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08632_ _03819_ u2.mem\[12\]\[9\] _03889_ _03891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_101_clock_I clknet_5_10_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08563_ _03825_ u2.mem\[10\]\[12\] _03850_ _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08145__I0 _03575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07514_ u2.mem\[54\]\[7\] _02883_ _02884_ u2.mem\[55\]\[7\] _02986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08494_ _03806_ _00149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07648__A2 _03116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08309__I _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09893__I0 _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07445_ u2.mem\[52\]\[5\] _02849_ _02850_ u2.mem\[21\]\[5\] _02919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_17_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07376_ u2.mem\[52\]\[4\] _02849_ _02850_ u2.mem\[21\]\[4\] _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_104_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08245__S _03634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09645__I0 _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09115_ _04205_ _00371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11452__I0 _05635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06327_ u2.mem\[153\]\[3\] _01707_ _01709_ u2.mem\[160\]\[3\] _01831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_109_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08073__A2 _03516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07281__B1 _02657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09046_ data_in_trans\[10\].data_sync _04160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06258_ u2.mem\[180\]\[1\] _01664_ _01667_ u2.mem\[150\]\[1\] _01764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08044__I _03501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_26_clock_I clknet_5_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06189_ _01685_ _01690_ _01695_ _01696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_150_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06499__I row_select_trans\[0\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09948_ _04728_ _00681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11507__I1 u2.mem\[168\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09804__S _04639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09879_ _04682_ _04683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_4047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08384__I0 _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11910_ _05947_ _01424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12890_ _00769_ clknet_leaf_57_clock u2.mem\[47\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07887__A2 _02553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09603__I _04500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10891__A1 _04072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11841_ _05904_ _05905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_166_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07639__A2 _03030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11772_ _05835_ u2.mem\[185\]\[4\] _05856_ _05862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06847__B1 _02130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13511_ _01390_ clknet_leaf_332_clock u2.mem\[188\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10723_ _05203_ _00981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11691__I0 _05792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13225__CLK clknet_leaf_301_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06962__I _02404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13442_ _01321_ clknet_leaf_364_clock u2.mem\[177\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10654_ _05151_ _05162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09636__I0 _04478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_303_clock_I clknet_5_20_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13373_ _01252_ clknet_leaf_371_clock u2.mem\[165\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10585_ _03707_ _05121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12324_ _00203_ clknet_leaf_95_clock u2.mem\[12\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07272__B1 _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13375__CLK clknet_leaf_367_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12255_ _00134_ clknet_leaf_241_clock u2.mem\[8\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07793__I _02444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11206_ _05507_ _05508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12186_ _00065_ clknet_leaf_59_clock u2.mem\[3\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07575__A1 u2.mem\[58\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06378__A2 _01656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11137_ _05339_ _05464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_1_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11068_ _05334_ _05420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08375__I0 _03680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10019_ _04769_ _00711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_4_15_0_clock_I clknet_3_7_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09513__I _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09875__I0 _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11682__I0 _05798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07230_ u2.mem\[3\]\[2\] _02470_ _02359_ _02707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09627__I0 _04469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07161_ _02425_ _02639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10394__I _04988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11434__I0 _05631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06112_ _01618_ _01607_ _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07092_ _02439_ _02440_ _02546_ _02443_ _02571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_69_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08850__I1 u2.mem\[17\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06043_ col_select_trans\[5\].data_sync _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07917__B _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12742__CLK clknet_leaf_24_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11737__I1 u2.mem\[183\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06369__A2 _01691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09802_ _03751_ _04542_ _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07994_ _01980_ _03250_ _03436_ _03457_ _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06945_ _02377_ _02391_ _02416_ _02424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA__12892__CLK clknet_leaf_222_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09733_ _04566_ _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_132_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08366__I0 _03663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07869__A2 _02420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09664_ _04546_ _00579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06876_ _02339_ _02354_ _02355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_252_clock_I clknet_5_19_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08615_ _03881_ _00195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09595_ _04473_ u2.mem\[34\]\[4\] _04506_ _04507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10569__I _03686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12122__CLK clknet_leaf_343_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13248__CLK clknet_leaf_308_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08546_ _03841_ _00166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08039__I data_in_trans\[2\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09866__I0 _04602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08477_ _03718_ u2.mem\[8\]\[14\] _03792_ _03795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_168_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07428_ u2.mem\[60\]\[5\] _02826_ _02827_ u2.mem\[62\]\[5\] _02902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_168_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12272__CLK clknet_leaf_179_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13398__CLK clknet_leaf_325_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07359_ u2.mem\[26\]\[4\] _02675_ _02676_ u2.mem\[10\]\[4\] _02834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_149_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07254__B1 _02591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11976__I1 u2.mem\[194\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10370_ _04918_ u2.mem\[52\]\[14\] _04981_ _04984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09029_ data_in_trans\[6\].data_sync _04147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12040_ col_select_trans\[1\].A clknet_leaf_316_clock col_select_trans\[1\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08502__I _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09534__S _04465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06780__A2 _02029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06957__I _02435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12942_ _00821_ clknet_leaf_220_clock u2.mem\[51\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09333__I _04335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12873_ _00752_ clknet_leaf_132_clock u2.mem\[46\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08109__I0 _03550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11824_ _05894_ _01391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09857__I0 _04589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12615__CLK clknet_leaf_137_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11755_ _05852_ _01364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07788__I _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06296__A1 u2.mem\[170\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06296__B2 u2.mem\[156\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10706_ _05126_ u2.mem\[60\]\[14\] _05189_ _05192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11686_ _05809_ _05810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_14_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13425_ _01304_ clknet_leaf_365_clock u2.mem\[174\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10637_ _05093_ u2.mem\[59\]\[0\] _05152_ _05153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12765__CLK clknet_leaf_219_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11103__I _05442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07245__B1 _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13356_ _01235_ clknet_leaf_377_clock u2.mem\[162\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10568_ _05109_ _00920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12307_ _00186_ clknet_leaf_111_clock u2.mem\[11\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10499_ _05020_ u2.mem\[55\]\[12\] _05066_ _05067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13287_ _01166_ clknet_leaf_382_clock u2.mem\[151\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11719__I1 u2.mem\[182\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12238_ _00117_ clknet_leaf_230_clock u2.mem\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12169_ _00048_ clknet_leaf_60_clock u2.mem\[2\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12145__CLK clknet_leaf_230_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08348__I0 _03714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06771__A2 _02065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06730_ u2.mem\[180\]\[2\] _02043_ _02013_ u2.mem\[172\]\[2\] _02213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xinput5 col_select_a[4] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_65_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06661_ _02145_ _02146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10389__I _04997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_382_clock clknet_5_0_0_clock clknet_leaf_382_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08400_ _03483_ _03748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09380_ _04370_ _00471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12295__CLK clknet_leaf_117_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06592_ _02026_ _01991_ _02077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09848__I0 _04576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08331_ _03700_ _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13540__CLK clknet_leaf_12_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06287__A1 u2.mem\[193\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08262_ _03647_ _00076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06287__B2 u2.mem\[177\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07213_ u2.mem\[5\]\[1\] _02689_ _02690_ u2.mem\[38\]\[1\] _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_140_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08193_ _03481_ _03605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_158_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06039__A1 col_select_trans\[0\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09619__S _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07144_ _02443_ _02614_ _02615_ _02442_ _02623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__11958__I1 u2.mem\[194\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07787__A1 u2.mem\[32\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_320_clock clknet_5_16_0_clock clknet_leaf_320_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_156_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07075_ _02463_ _02515_ _02516_ _02442_ _02554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_133_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06026_ u2.driver_mem\[15\] _01508_ _01535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07539__A1 u2.mem\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_335_clock clknet_5_18_0_clock clknet_leaf_335_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09354__S _04351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input37_I row_select_a[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06211__A1 u2.mem\[154\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06211__B2 u2.mem\[162\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07977_ _03437_ _03438_ _03439_ _03440_ _03441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06762__A2 _02097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09716_ _04566_ _04580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06928_ _02346_ _02407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12638__CLK clknet_leaf_215_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09647_ _04489_ u2.mem\[35\]\[11\] _04532_ _04536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06859_ _02008_ row_select_trans\[4\].data_sync _02338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_55_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09578_ _04173_ _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08529_ _03830_ u2.mem\[9\]\[14\] _03826_ _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11646__I0 _05756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11124__S _05453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07475__B1 _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06278__B2 u2.mem\[150\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11540_ _05679_ _05719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_169_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11471_ _05675_ _01257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10963__S _05356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09529__S _04458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07227__B1 _02452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10422_ _05020_ u2.mem\[53\]\[12\] _05021_ _05022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13210_ _01089_ clknet_leaf_298_clock u2.mem\[138\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12018__CLK clknet_leaf_315_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08433__S _03768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08814__I1 u2.mem\[16\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07778__B2 u2.mem\[4\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10353_ _04974_ _00840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13141_ _01020_ clknet_leaf_20_clock u2.mem\[63\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07242__A3 _02713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13072_ _00951_ clknet_leaf_335_clock u2.mem\[59\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10284_ _04907_ u2.mem\[50\]\[9\] _04933_ _04935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12168__CLK clknet_leaf_62_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12023_ net33 clknet_2_2__leaf_clock_a mem_address_trans\[9\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11794__S _05865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13413__CLK clknet_5_5_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06738__C1 u2.mem\[168\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06202__A1 _01596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07950__A1 _03399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09063__I data_in_trans\[14\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13563__CLK clknet_leaf_10_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12925_ _00804_ clknet_leaf_221_clock u2.mem\[50\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11885__I0 u2.mem\[192\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06505__A2 _01989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_148_clock_I clknet_5_13_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12856_ _00735_ clknet_leaf_143_clock u2.mem\[45\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11807_ _05884_ _01384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10937__I _05336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12787_ _00666_ clknet_leaf_31_clock u2.mem\[41\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11034__S _05394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11738_ _05842_ _01357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07311__I _02384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11969__S _05980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12076__D data_in_trans\[13\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11669_ _05799_ _01331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_200_clock_I clknet_5_31_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09439__S _04406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07218__B1 _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13408_ _01287_ clknet_leaf_319_clock u2.mem\[171\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10672__I _04862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07467__B _02749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13339_ _01218_ clknet_leaf_1_clock u2.mem\[160\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08569__I0 _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06992__A2 _02470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07900_ u2.mem\[18\]\[13\] _03318_ _03319_ u2.mem\[19\]\[13\] _03366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_97_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13093__CLK clknet_leaf_20_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08880_ _04010_ u2.mem\[18\]\[0\] _04051_ _04052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09930__A2 _04659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07831_ u2.mem\[57\]\[12\] _03137_ _03138_ u2.mem\[41\]\[12\] _03298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06597__I _02081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10128__I0 _04815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07762_ u2.mem\[60\]\[11\] _03059_ _03060_ u2.mem\[62\]\[11\] _03230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09501_ _04446_ _00516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06713_ u2.mem\[153\]\[1\] _02196_ _02131_ u2.mem\[152\]\[1\] _02197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07693_ _03157_ _03158_ _03159_ _03162_ _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_38_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09432_ _04373_ u2.mem\[30\]\[7\] _04401_ _04405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12930__CLK clknet_leaf_151_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06644_ _02128_ _02129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11628__I0 _05752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09363_ _04356_ u2.mem\[29\]\[0\] _04358_ _04359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06575_ _01998_ _02060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09297__I1 u2.mem\[27\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08314_ _03686_ _03687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09294_ _04312_ _04318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_166_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08245_ _03552_ u2.mem\[4\]\[3\] _03634_ _03638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10783__S _05242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07209__B1 _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09349__S _04346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06680__A1 u2.mem\[169\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11005__A1 _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08176_ _03563_ u2.mem\[2\]\[8\] _03595_ _03596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06680__B2 u2.mem\[147\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07127_ _02605_ _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11800__I0 _05868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10582__I _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09148__I _04223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07058_ _02536_ _02537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07775__A4 _03242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06983__A2 _02457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06009_ u2.driver_mem\[1\] _01517_ _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xclkbuf_leaf_274_clock clknet_5_23_0_clock clknet_leaf_274_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_121_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09084__S _04187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08980__I0 _04037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07932__B2 u2.mem\[59\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10119__I0 _04806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_289_clock clknet_5_21_0_clock clknet_leaf_289_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_1_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11867__I0 _05911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10971_ _05349_ u2.mem\[135\]\[4\] _05355_ _05361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10958__S _05336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12710_ _00589_ clknet_leaf_65_clock u2.mem\[36\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07696__B1 _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_3_clock clknet_5_0_0_clock clknet_leaf_3_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_71_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12641_ _00520_ clknet_leaf_157_clock u2.mem\[32\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10757__I _03716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09288__I1 u2.mem\[27\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12572_ _00451_ clknet_leaf_201_clock u2.mem\[28\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07131__I _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11523_ _05662_ _05707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10693__S _05184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_227_clock clknet_5_22_0_clock clknet_leaf_227_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_89_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06970__I _02448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11454_ _03490_ _05662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11588__I _05747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10405_ _05009_ u2.mem\[53\]\[7\] _05002_ _05010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11385_ _05591_ u2.mem\[161\]\[3\] _05616_ _05620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13124_ _01003_ clknet_leaf_20_clock u2.mem\[62\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10336_ _04862_ _04964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12803__CLK clknet_leaf_113_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_74_clock_I clknet_5_8_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06974__A2 _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08897__I _04050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10267_ _04925_ _00803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13055_ _00934_ clknet_leaf_254_clock u2.mem\[58\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12006_ mem_address_trans\[0\].A clknet_leaf_315_clock mem_address_trans\[0\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06411__S _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10198_ _04808_ u2.mem\[48\]\[11\] _04875_ _04879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08971__I0 _04028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12953__CLK clknet_leaf_148_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10868__S _05286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_299_clock_I clknet_5_21_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12908_ _00787_ clknet_leaf_202_clock u2.mem\[49\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07687__B1 _03156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10530__I0 _05014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07151__A2 _02627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13309__CLK clknet_leaf_363_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12839_ _00718_ clknet_leaf_131_clock u2.mem\[44\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06360_ u2.mem\[190\]\[4\] _01703_ _01705_ u2.mem\[194\]\[4\] _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_61_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08137__I _03524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06291_ u2.mem\[152\]\[2\] _01713_ _01715_ u2.mem\[148\]\[2\] _01796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10833__I1 _03532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13459__CLK clknet_leaf_362_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_351_clock_I clknet_5_4_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08030_ _03490_ _03491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09169__S _04236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06880__I _02358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput30 mem_address_a[6] net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput41 row_select_a[4] net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_174_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12483__CLK clknet_leaf_119_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10210__A2 _04863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09981_ _04747_ _00695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08954__A3 _03632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08932_ _04028_ u2.mem\[19\]\[6\] _04079_ _04082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08863_ _04039_ u2.mem\[17\]\[11\] _04033_ _04040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08962__I0 _04019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07814_ u2.mem\[44\]\[12\] _03122_ _03123_ u2.mem\[42\]\[12\] _03281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_3709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08794_ _03994_ _00261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07216__I _02621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07390__A2 _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07745_ u2.mem\[1\]\[11\] _03030_ _03031_ u2.mem\[7\]\[11\] _03213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_42_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10778__S _05237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07676_ u2.mem\[28\]\[9\] _03074_ _03075_ u2.mem\[31\]\[9\] _03146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10521__I0 _05005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09415_ _04394_ _04011_ _04395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06627_ u2.mem\[166\]\[0\] _02097_ _02099_ u2.mem\[161\]\[0\] _02111_ _02112_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_80_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07693__A3 _03159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09346_ _04348_ _00459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06558_ _02042_ _02043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08047__I _03488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11777__A2 _05847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10824__I1 _03522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09277_ _04307_ _00431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06489_ u2.mem\[0\]\[14\] _01976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_103_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09690__I1 u2.mem\[36\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09079__S _04182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06653__A1 u2.mem\[153\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08228_ _03577_ u2.mem\[3\]\[14\] _03623_ _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06653__B2 u2.mem\[160\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12826__CLK clknet_leaf_129_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10018__S _04767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08159_ _03586_ _00034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11201__I _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07602__B1 _03072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11170_ _05485_ _01146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06956__A2 _02433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10121_ _04808_ u2.mem\[46\]\[11\] _04830_ _04834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12976__CLK clknet_leaf_264_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10052_ _04789_ _00724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07905__A1 u2.mem\[6\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07905__B2 u2.mem\[47\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07381__A2 _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10688__S _05179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_151_clock clknet_5_24_0_clock clknet_leaf_151_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_28_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07669__B1 _03138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08158__S _03585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10512__I0 _04992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10954_ _05349_ u2.mem\[134\]\[4\] _05336_ _05350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12356__CLK clknet_leaf_93_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10885_ _05000_ _05305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12624_ _00503_ clknet_leaf_183_clock u2.mem\[31\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06892__A1 _02339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09130__I0 _04154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_166_clock clknet_5_26_0_clock clknet_leaf_166_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12555_ _00434_ clknet_leaf_206_clock u2.mem\[27\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10815__I1 _03512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07796__I _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11506_ _05697_ _01270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12486_ _00365_ clknet_leaf_107_clock u2.mem\[22\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07987__A4 _03450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11437_ _05652_ _01246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11240__I1 u2.mem\[152\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11368_ _05610_ _01219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13107_ _00986_ clknet_leaf_17_clock u2.mem\[61\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10319_ _04904_ u2.mem\[51\]\[8\] _04954_ _04955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11299_ _04333_ _05566_ _05567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_65_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_104_clock clknet_5_10_0_clock clknet_leaf_104_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13038_ _00917_ clknet_leaf_263_clock u2.mem\[57\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11982__S _05985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11781__I _03661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_119_clock clknet_5_14_0_clock clknet_leaf_119_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07530_ u2.mem\[29\]\[7\] _02835_ _02836_ u2.mem\[11\]\[7\] _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11456__A1 _04179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10503__I0 _05025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07461_ u2.mem\[40\]\[6\] _02789_ _02790_ u2.mem\[30\]\[6\] _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_34_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10397__I _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13281__CLK clknet_leaf_384_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09200_ _04257_ _00404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06412_ _01911_ _01912_ _01913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__06883__A1 _02338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07392_ _02431_ _02866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12849__CLK clknet_leaf_154_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09121__I0 _04140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09131_ _04214_ _00378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06343_ u2.mem\[174\]\[4\] _01657_ _01658_ u2.mem\[155\]\[4\] _01661_ u2.mem\[181\]\[4\]
+ _01846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_124_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10806__I1 _03499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06824__B _02304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09062_ _04172_ _00351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06274_ u2.mem\[184\]\[2\] _01778_ _01753_ _01779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_147_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08013_ _03468_ _03475_ _05992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12999__CLK clknet_leaf_149_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11021__I _05351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09627__S _04522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06115__I _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11231__I1 u2.mem\[151\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06938__A2 _02400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09964_ _04737_ _00688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12229__CLK clknet_leaf_73_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08330__I _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08915_ _03484_ _03747_ _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_09895_ _04582_ _04694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11892__S _05937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08846_ _03683_ _04028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10742__I0 _05216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08777_ _03981_ _00257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07728_ u2.mem\[17\]\[10\] _03079_ _03080_ u2.mem\[24\]\[10\] _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10301__S _04944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_22_clock_I clknet_5_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07659_ u2.mem\[43\]\[9\] _03053_ _03054_ u2.mem\[20\]\[9\] _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_26_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_83_clock clknet_5_9_0_clock clknet_leaf_83_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06874__A1 _01989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10670_ _05128_ u2.mem\[59\]\[15\] _05167_ _05171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_159_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08706__S _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09112__I0 _04119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09329_ _04256_ u2.mem\[28\]\[2\] _04336_ _04339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12340_ _00219_ clknet_leaf_94_clock u2.mem\[13\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08505__I _03687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_98_clock clknet_5_10_0_clock clknet_leaf_98_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_33_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_247_clock_I clknet_5_18_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12271_ _00150_ clknet_leaf_177_clock u2.mem\[9\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10971__S _05355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09537__S _04465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11222_ _05519_ _05520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_134_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_21_clock clknet_5_2_0_clock clknet_leaf_21_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_107_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11153_ _05474_ _05475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_110_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10104_ _04824_ _00741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13154__CLK clknet_leaf_281_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11084_ _05431_ _01114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10035_ _04778_ _00718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08000__B1 _03462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_36_clock clknet_5_3_0_clock clknet_leaf_36_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11986_ _03534_ _05972_ _05991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_17_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10937_ _05336_ _05337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_44_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06314__B1 _01664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06865__A1 _02340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08616__S _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10868_ _05207_ u2.mem\[129\]\[5\] _05286_ _05293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12607_ _00486_ clknet_leaf_159_clock u2.mem\[30\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10945__I _05342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10799_ _05251_ _01009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06617__A1 u2.mem\[187\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12538_ _00417_ clknet_leaf_117_clock u2.mem\[25\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07814__B1 _03123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06617__B2 u2.mem\[192\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12469_ _00348_ clknet_leaf_104_clock u2.mem\[21\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11776__I _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11913__A2 _05926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09246__I _04289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07593__A2 _03062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08150__I _03534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06961_ _02388_ _02440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_41_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08700_ _03937_ _00224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12521__CLK clknet_leaf_125_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09680_ _04555_ _00586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06892_ _02339_ _02338_ _02344_ _02371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09182__S _04241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09590__I0 _04469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08393__I1 u2.mem\[6\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08631_ _03890_ _00202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07896__A3 _03360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08562_ _03834_ _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10121__S _04830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07513_ u2.mem\[50\]\[7\] _02880_ _02881_ u2.mem\[51\]\[7\] _02985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_39_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_196_clock_I clknet_5_31_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08493_ _03805_ u2.mem\[9\]\[3\] _03799_ _03806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_1_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09893__I1 u2.mem\[41\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06856__A1 _02324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07444_ u2.mem\[17\]\[5\] _02846_ _02847_ u2.mem\[24\]\[5\] _02918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07375_ _02600_ _02850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13027__CLK clknet_leaf_30_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09114_ _04128_ u2.mem\[23\]\[1\] _04203_ _04205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06608__A1 _02031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07805__B1 _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08325__I _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06326_ u2.mem\[190\]\[3\] _01702_ _01704_ u2.mem\[194\]\[3\] _01830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11452__I1 u2.mem\[165\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11887__S _05932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09045_ _04159_ _00347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06257_ u2.mem\[174\]\[1\] _01657_ _01659_ u2.mem\[155\]\[1\] _01661_ u2.mem\[181\]\[1\]
+ _01763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_50_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12051__CLK clknet_2_1__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13177__CLK clknet_leaf_292_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08261__S _03644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06188_ u2.mem\[146\]\[0\] _01692_ _01694_ u2.mem\[186\]\[0\] _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_104_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11686__I _05809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07033__A1 _02441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10963__I0 _05335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07584__A2 _03053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08060__I data_in_trans\[7\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09947_ _04698_ u2.mem\[42\]\[7\] _04724_ _04728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06792__B1 _02086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06792__C2 _02093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08995__I _04118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09878_ _04249_ _04659_ _04682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08384__I1 u2.mem\[6\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08829_ _04016_ _00274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10031__S _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11840_ _04393_ _05886_ _05904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_166_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06448__C _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11771_ _05861_ _01371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13510_ _01389_ clknet_leaf_347_clock u2.mem\[188\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10722_ _05202_ u2.mem\[61\]\[3\] _05196_ _05203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06847__B2 u2.mem\[152\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11840__A1 _04393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11691__I1 u2.mem\[180\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13441_ _01320_ clknet_leaf_363_clock u2.mem\[177\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10653_ _05161_ _00953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13372_ _01251_ clknet_leaf_371_clock u2.mem\[165\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10584_ _05120_ _00925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12323_ _00202_ clknet_leaf_113_clock u2.mem\[12\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07272__B2 u2.mem\[33\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09267__S _04300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12254_ _00133_ clknet_leaf_227_clock u2.mem\[8\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11205_ _03498_ _05507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12544__CLK clknet_leaf_188_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12185_ _00064_ clknet_leaf_59_clock u2.mem\[3\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07575__A2 _03044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11136_ _05463_ _01134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11067_ _05419_ _01109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10706__I0 _05126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12694__CLK clknet_leaf_82_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10018_ _04694_ u2.mem\[44\]\[5\] _04767_ _04769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07314__I _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06358__C _01860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11969_ _05211_ u2.mem\[194\]\[7\] _05980_ _05982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_17_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06302__A3 _01793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06374__B _01876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07160_ _02419_ _02638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12074__CLK clknet_leaf_362_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11434__I1 u2.mem\[164\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06111_ _01558_ _01568_ _01585_ _01618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_157_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07263__A1 _02724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07091_ u2.mem\[26\]\[0\] _02567_ _02569_ u2.mem\[10\]\[0\] _02570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06042_ _01548_ _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07015__A1 _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07566__A2 _03036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09801_ _04637_ _00625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07993_ _03441_ _03446_ _03451_ _03456_ _03457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_115_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09732_ _04591_ _04592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06944_ _02373_ _02423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_80_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09563__I0 _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09663_ _04467_ u2.mem\[36\]\[1\] _04544_ _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06875_ row_select_trans\[1\].data_sync _02009_ _02354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08614_ _03801_ u2.mem\[12\]\[1\] _03879_ _03881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09594_ _04500_ _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_82_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09315__I0 _04281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08545_ _03807_ u2.mem\[10\]\[4\] _03840_ _03841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11122__I0 _05424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09866__I1 u2.mem\[40\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12417__CLK clknet_leaf_171_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08476_ _03794_ _00143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09491__A2 mem_address_trans\[5\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07427_ u2.mem\[61\]\[5\] _02899_ _02900_ u2.mem\[63\]\[5\] _02901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10585__I _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07358_ _02825_ _02828_ _02831_ _02832_ _02833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_136_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06309_ u2.mem\[184\]\[3\] _01778_ _01753_ _01813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__12567__CLK clknet_leaf_116_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07289_ u2.mem\[37\]\[3\] _02537_ _02539_ u2.mem\[59\]\[3\] _02765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_163_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09028_ _04146_ _00343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11189__I0 _05468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07006__A1 _02377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07021__A4 _02458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06765__B1 _02200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12941_ _00820_ clknet_leaf_221_clock u2.mem\[51\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12872_ _00751_ clknet_leaf_133_clock u2.mem\[46\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07190__B1 _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09306__I0 _04272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09550__S _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11823_ _05876_ u2.mem\[188\]\[5\] _05887_ _05894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09857__I1 u2.mem\[40\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06973__I _02451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12097__CLK clknet_leaf_246_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11754_ _05831_ u2.mem\[184\]\[2\] _05849_ _05852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13342__CLK clknet_leaf_2_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10705_ _05191_ _00975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11685_ _04094_ _05808_ _05809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13424_ _01303_ clknet_leaf_361_clock u2.mem\[174\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10636_ _05151_ _05152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_70_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13355_ _01234_ clknet_leaf_370_clock u2.mem\[162\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13492__CLK clknet_leaf_307_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10567_ _05108_ u2.mem\[57\]\[6\] _05104_ _05109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12306_ _00185_ clknet_leaf_173_clock u2.mem\[11\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_144_clock_I clknet_5_13_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13286_ _01165_ clknet_leaf_381_clock u2.mem\[151\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10498_ _05050_ _05066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_29_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12237_ _00116_ clknet_leaf_226_clock u2.mem\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07309__I _02360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06213__I _01719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12168_ _00047_ clknet_leaf_62_clock u2.mem\[2\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11119_ _05452_ _05453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_12099_ _01497_ clknet_leaf_247_clock u2.active_mem\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput6 col_select_a[5] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_76_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06660_ _02005_ _02125_ _02145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_37_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07044__I _02448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09460__S _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07720__A2 _03137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06591_ _02075_ _02076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09848__I1 u2.mem\[40\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_69_clock_I clknet_5_9_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08330_ _03699_ _03700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08261_ _03568_ u2.mem\[4\]\[10\] _03644_ _03647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07212_ _02628_ _02690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08192_ _03604_ _00049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07236__A1 _02709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06039__A2 col_select_trans\[1\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07143_ _02621_ _02622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_146_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07074_ _02552_ _02553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_145_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06025_ _01516_ _01533_ _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10918__I0 _05307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07539__A2 _02922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07003__A4 _02401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06211__A2 _01699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07976_ u2.mem\[57\]\[15\] _02548_ _02550_ u2.mem\[41\]\[15\] _03440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09434__I _04395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09715_ _04578_ _04579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06927_ _02405_ _02400_ _02392_ _02406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA_clkbuf_leaf_346_clock_I clknet_5_5_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09646_ _04535_ _00572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06858_ _01878_ _01996_ _02337_ _01479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_3_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11894__I1 _03514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07711__A2 _03122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09577_ _04495_ _00543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06789_ _02255_ _02260_ _02265_ _02270_ _02271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08528_ _03717_ _03830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11646__I1 u2.mem\[177\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08459_ _03684_ u2.mem\[8\]\[6\] _03782_ _03785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11470_ _05674_ u2.mem\[166\]\[3\] _05665_ _05675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10421_ _04988_ _05021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_51_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13140_ _01019_ clknet_leaf_17_clock u2.mem\[63\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10352_ _04900_ u2.mem\[52\]\[6\] _04971_ _04974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07242__A4 _02718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13071_ _00950_ clknet_leaf_250_clock u2.mem\[59\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10283_ _04934_ _00810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12022_ mem_address_trans\[8\].A clknet_leaf_321_clock mem_address_trans\[8\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06738__B1 _02087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11582__I0 _05717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06202__A2 _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06968__I _02446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09527__I0 _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07950__A2 _03404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12924_ _00803_ clknet_leaf_221_clock u2.mem\[50\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11885__I1 _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07702__A2 _03030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12855_ _00734_ clknet_leaf_143_clock u2.mem\[45\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06917__B _02393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07799__I _02464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_70_clock_I clknet_5_8_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12732__CLK clknet_leaf_271_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11315__S _05576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11806_ _05874_ u2.mem\[187\]\[4\] _05878_ _05884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12786_ _00665_ clknet_leaf_338_clock u2.mem\[41\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11737_ _05829_ u2.mem\[183\]\[1\] _05840_ _05842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06208__I _01714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11668_ _05798_ u2.mem\[178\]\[5\] _05787_ _05799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12882__CLK clknet_leaf_243_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13407_ _01286_ clknet_leaf_320_clock u2.mem\[171\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08266__I0 _03572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10953__I _05348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10619_ _05142_ _00938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07748__B _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11599_ _05755_ _01305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07769__A2 _03074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08423__I _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13338_ _01217_ clknet_leaf_6_clock u2.mem\[159\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_295_clock_I clknet_5_21_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12092__D inverter_select_trans.A vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12112__CLK clknet_leaf_347_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13238__CLK clknet_leaf_302_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13269_ _01148_ clknet_leaf_384_clock u2.mem\[148\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07039__I _02517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11784__I _03665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07830_ u2.mem\[37\]\[12\] _03295_ _03296_ u2.mem\[59\]\[12\] _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_42_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12262__CLK clknet_leaf_72_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09518__I0 _04380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13388__CLK clknet_leaf_372_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07761_ u2.mem\[61\]\[11\] _03132_ _03133_ u2.mem\[63\]\[11\] _03229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11325__I0 _05556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09500_ _04362_ u2.mem\[32\]\[2\] _04443_ _04446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06712_ _02136_ _02196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07692_ u2.mem\[6\]\[9\] _03160_ _03161_ u2.mem\[47\]\[9\] _03162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07154__B1 _02535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09431_ _04404_ _00488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06643_ _02107_ _02041_ _02128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11225__S _05520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09362_ _04357_ _04358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_40_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06574_ _02058_ _02059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11628__I1 u2.mem\[176\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08313_ data_in_trans\[7\].data_sync _03686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07457__A1 _02907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09293_ _04317_ _00437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08244_ _03637_ _00068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08257__I0 _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08175_ _03584_ _03595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_146_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10064__I0 _04797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07126_ _02587_ _02588_ _02424_ _02589_ _02605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__11800__I1 u2.mem\[187\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07057_ _02455_ _02510_ _02511_ _02474_ _02536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_134_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06008_ _01507_ _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12605__CLK clknet_leaf_216_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11564__I0 _05713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09509__I0 _04371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07959_ u2.mem\[16\]\[15\] _03266_ _03267_ u2.mem\[33\]\[15\] _03423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_101_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_2_0__f_clock_a_I clknet_0_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10970_ _05360_ _01071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11867__I1 u2.mem\[191\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09629_ _04471_ u2.mem\[35\]\[3\] _04522_ _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11135__S _05462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12640_ _00519_ clknet_leaf_157_clock u2.mem\[32\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08508__I _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12571_ _00450_ clknet_leaf_186_clock u2.mem\[28\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11522_ _05706_ _01277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06120__A1 u2.mem\[184\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12135__CLK clknet_leaf_38_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08248__I0 _03554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11453_ _05661_ _01253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10773__I _05231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09996__I0 _04709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10404_ _03686_ _05009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11384_ _05619_ _01226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13123_ _01002_ clknet_leaf_21_clock u2.mem\[62\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_152_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10335_ _04963_ _00833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_17_clock_I clknet_5_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_381_clock clknet_5_0_0_clock clknet_leaf_381_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12285__CLK clknet_leaf_194_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13054_ _00933_ clknet_leaf_274_clock u2.mem\[58\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10266_ _04889_ u2.mem\[50\]\[1\] _04923_ _04925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13530__CLK clknet_leaf_325_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11555__I0 _05719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12005_ net24 clknet_2_0__leaf_clock_a mem_address_trans\[0\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10197_ _04878_ _00780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09074__I _04181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07923__A2 _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08971__I1 u2.mem\[20\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11307__I0 _05552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12907_ _00786_ clknet_leaf_207_clock u2.mem\[49\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07687__A1 u2.mem\[5\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10948__I _04134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11045__S _05404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12838_ _00717_ clknet_leaf_87_clock u2.mem\[44\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07322__I _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07439__A1 u2.mem\[28\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08487__I0 _03801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12087__D net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12769_ _00648_ clknet_leaf_152_clock u2.mem\[40\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06290_ u2.mem\[153\]\[2\] _01708_ _01710_ u2.mem\[160\]\[2\] _01795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_334_clock clknet_5_18_0_clock clknet_leaf_334_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_30_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08239__I0 _03538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput20 data_in_a[7] net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__10683__I _05173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13060__CLK clknet_leaf_29_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput31 mem_address_a[7] net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__06662__A2 _02011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput42 row_select_a[5] net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_50_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09987__I0 _04700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12628__CLK clknet_leaf_95_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11794__I0 _05876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_349_clock clknet_5_6_0_clock clknet_leaf_349_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09980_ _04694_ u2.mem\[43\]\[5\] _04745_ _04747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08931_ _04081_ _00311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12778__CLK clknet_leaf_141_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08862_ _03704_ _04039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10124__S _04835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06178__A1 u2.mem\[191\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06178__B2 u2.mem\[179\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08962__I1 u2.mem\[20\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07813_ _03272_ _03273_ _03276_ _03279_ _03280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_97_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08793_ _03911_ u2.mem\[16\]\[3\] _03990_ _03994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07390__A3 _02855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07744_ u2.mem\[15\]\[11\] _03027_ _03028_ u2.mem\[13\]\[11\] _03212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12008__CLK clknet_leaf_315_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07675_ u2.mem\[9\]\[9\] _03071_ _03072_ u2.mem\[25\]\[9\] _03145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_129_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09414_ _04393_ _04394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06626_ _02102_ _02106_ _02110_ _02111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09345_ _04272_ u2.mem\[28\]\[9\] _04346_ _04348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12158__CLK clknet_leaf_219_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06557_ _02041_ _02015_ _02042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10794__S _05247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09276_ _04281_ u2.mem\[26\]\[13\] _04305_ _04307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06102__A1 _01547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06488_ _01973_ _01970_ _01974_ _01975_ _01462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_21_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08227_ _03625_ _00063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06653__A2 _02136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09159__I _04225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09978__I0 _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08158_ _03538_ u2.mem\[2\]\[0\] _03585_ _03586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08063__I _03488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13553__CLK clknet_leaf_10_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11785__I0 _05870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07109_ _02413_ _02588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_88_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08998__I _03987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08089_ _03534_ _03528_ _03535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09095__S _04192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10120_ _04833_ _00748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10034__S _04777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10051_ _04788_ u2.mem\[45\]\[2\] _04784_ _04789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08012__B _03474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07905__A2 _02622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10969__S _05356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07118__B1 _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_243_clock_I clknet_5_24_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08439__S _03768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09622__I _04521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09902__I0 _04698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10953_ _05348_ _05349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08238__I _03633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10884_ _05304_ _01041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07684__A4 _03153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12623_ _00502_ clknet_leaf_182_clock u2.mem\[31\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06892__A2 _02338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12554_ _00433_ clknet_leaf_123_clock u2.mem\[26\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10976__A1 _04224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11505_ _05677_ u2.mem\[168\]\[4\] _05691_ _05697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12485_ _00364_ clknet_leaf_109_clock u2.mem\[22\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09969__I0 _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11436_ _05633_ u2.mem\[164\]\[4\] _05646_ _05652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08902__S _04061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08641__I0 _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11367_ _05587_ u2.mem\[160\]\[1\] _05608_ _05610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06930__B _02406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13106_ _00985_ clknet_leaf_330_clock u2.mem\[61\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10318_ _04943_ _04954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08701__I _03721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11298_ _05442_ _05566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_80_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13037_ _00916_ clknet_leaf_282_clock u2.mem\[57\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_152_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10249_ _04604_ _04913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07357__B1 _02672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06221__I _01726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11456__A2 _05645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13426__CLK clknet_leaf_365_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07460_ u2.mem\[32\]\[6\] _02786_ _02787_ u2.mem\[2\]\[6\] _02933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_39_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06332__A1 u2.mem\[170\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06332__B2 u2.mem\[156\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06411_ u2.select_mem_row\[4\] u2.select_mem_col\[4\] _01515_ _01912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07391_ _01843_ _02784_ _02824_ _02865_ _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_273_clock clknet_5_23_0_clock clknet_leaf_273_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_37_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11503__S _05692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09130_ _04154_ u2.mem\[23\]\[8\] _04213_ _04214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06342_ u2.mem\[189\]\[4\] _01650_ _01663_ u2.mem\[180\]\[4\] _01651_ u2.mem\[176\]\[4\]
+ _01845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__12450__CLK clknet_leaf_169_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13576__CLK clknet_leaf_32_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09061_ _04171_ u2.mem\[21\]\[13\] _04168_ _04172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10119__S _04830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06273_ _01626_ _01778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07832__A1 _03291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08880__I0 _04010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08012_ _01613_ _03471_ _03474_ _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_288_clock clknet_5_20_0_clock clknet_leaf_288_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_128_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08632__I0 _03819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_192_clock_I clknet_5_30_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07596__B1 _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06399__B2 u2.mem\[162\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11392__A1 _05295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_2_clock clknet_5_0_0_clock clknet_leaf_2_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_171_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06938__A3 _02416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09963_ _04714_ u2.mem\[42\]\[14\] _04734_ _04737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08611__I _03878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_211_clock clknet_5_28_0_clock clknet_leaf_211_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11519__I0 _05677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08914_ _04070_ _00305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09894_ _04693_ _00662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09643__S _04532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08845_ _04027_ _00279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10789__S _05242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10742__I1 u2.mem\[61\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08776_ _03938_ u2.mem\[15\]\[15\] _03977_ _03981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_226_clock clknet_5_28_0_clock clknet_leaf_226_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_113_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08259__S _03644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input12_I data_in_a[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07727_ u2.mem\[23\]\[10\] _03148_ _03149_ u2.mem\[22\]\[10\] _03196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_150_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08699__I0 _03936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07658_ u2.mem\[49\]\[9\] _03050_ _03051_ u2.mem\[46\]\[9\] _03128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_144_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06323__B2 u2.mem\[161\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06609_ _02093_ _02094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06874__A2 row_select_trans\[5\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07589_ _02543_ _03060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11413__S _05638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09328_ _04338_ _00451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08076__A1 _01966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09259_ _04297_ _00423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10029__S _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12943__CLK clknet_leaf_242_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12270_ _00149_ clknet_leaf_199_clock u2.mem\[9\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11758__I0 _05835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11221_ _05354_ _05482_ _05519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_49_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08623__I0 _03810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07587__B1 _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08521__I _03708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11152_ _04071_ _05443_ _05474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10103_ _04790_ u2.mem\[46\]\[3\] _04820_ _04824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11083_ _05430_ u2.mem\[142\]\[4\] _05421_ _05431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09553__S _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10034_ _04709_ u2.mem\[44\]\[12\] _04777_ _04778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10699__S _05184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11930__I0 _05211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11882__I _05928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12323__CLK clknet_leaf_113_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06976__I _02362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10498__I _05050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11985_ _05990_ _01456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10936_ _04180_ _05317_ _05336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06314__A1 u2.mem\[172\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12473__CLK clknet_leaf_169_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06314__B2 u2.mem\[180\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10867_ _05292_ _01036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11323__S _05575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12606_ _00485_ clknet_leaf_202_clock u2.mem\[30\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08067__A1 _01954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10798_ _05229_ u2.mem\[62\]\[15\] _05247_ _05251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07600__I _02571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12537_ _00416_ clknet_leaf_118_clock u2.mem\[25\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06617__A2 _02100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12468_ _00347_ clknet_leaf_106_clock u2.mem\[21\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08632__S _03889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07290__A2 _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11419_ _05631_ u2.mem\[163\]\[3\] _05638_ _05642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08614__I0 _03801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12399_ _00278_ clknet_leaf_172_clock u2.mem\[17\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07578__B1 _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06960_ _02386_ _02439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_113_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input4_I col_select_a[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06891_ _02369_ _02370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_95_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11921__I0 _05911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08630_ _03816_ u2.mem\[12\]\[8\] _03889_ _03890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06886__I _02364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10402__S _05002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06553__A1 _01999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07750__B1 _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07896__A4 _03361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12816__CLK clknet_leaf_167_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06819__C _02299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08561_ _03849_ _00173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07512_ _02979_ _02980_ _02981_ _02983_ _02984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_63_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_139_clock_I clknet_5_12_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08492_ _03670_ _03805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08807__S _04000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07502__B1 _02867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07443_ u2.mem\[23\]\[5\] _02915_ _02916_ u2.mem\[22\]\[5\] _02917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_165_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06856__A2 _02329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11233__S _05519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12966__CLK clknet_leaf_105_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08058__A1 _03512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07374_ _02598_ _02849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07510__I _02358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09113_ _04204_ _00370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06325_ u2.mem\[144\]\[3\] _01671_ _01673_ u2.mem\[182\]\[3\] _01829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_31_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06608__A2 _02070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09044_ _04158_ u2.mem\[21\]\[9\] _04155_ _04159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07281__A2 _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06256_ _01756_ _01759_ _01760_ _01761_ _01762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__08542__S _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11990__CLK clknet_leaf_334_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06187_ _01693_ _01694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_150_clock clknet_5_24_0_clock clknet_leaf_150_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07569__B1 _02884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10412__I0 _05014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07033__A2 _02429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08341__I _03708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09946_ _04727_ _00680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06792__A1 u2.mem\[151\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06792__B2 u2.mem\[158\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09877_ _04564_ _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08828_ _04010_ u2.mem\[17\]\[0\] _04015_ _04016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10312__S _04949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12496__CLK clknet_leaf_175_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08759_ _03971_ _00249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11770_ _05833_ u2.mem\[185\]\[3\] _05857_ _05861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10721_ _04997_ _05202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06847__A2 _02128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13440_ _01319_ clknet_leaf_354_clock u2.mem\[176\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09097__I0 _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10652_ _05110_ u2.mem\[59\]\[7\] _05157_ _05161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_103_clock clknet_5_10_0_clock clknet_leaf_103_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_70_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06464__C _01949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13371_ _01250_ clknet_leaf_375_clock u2.mem\[165\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10982__S _05365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08844__I0 _04026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10583_ _05119_ u2.mem\[57\]\[11\] _05113_ _05120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12322_ _00201_ clknet_leaf_167_clock u2.mem\[12\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07272__A2 _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08452__S _03777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13121__CLK clknet_leaf_330_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11877__I _05928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12253_ _00132_ clknet_leaf_227_clock u2.mem\[8\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_118_clock clknet_5_14_0_clock clknet_leaf_118_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_154_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11204_ _05506_ _01159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12184_ _00063_ clknet_leaf_62_clock u2.mem\[3\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13271__CLK clknet_leaf_4_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11135_ _05460_ u2.mem\[146\]\[0\] _05462_ _05463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11066_ _05392_ u2.mem\[141\]\[5\] _05412_ _05419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10706__I1 u2.mem\[60\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10017_ _04768_ _00710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07732__B1 _03156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_140_clock_I clknet_5_12_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12989__CLK clknet_leaf_274_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11968_ _05981_ _01448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10095__A1 _04394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10956__I _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10919_ _05325_ _01055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11899_ _05941_ _01419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12219__CLK clknet_leaf_229_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06302__A4 _01806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09088__I0 _04148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12095__D _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13569_ _01448_ clknet_leaf_12_clock u2.mem\[194\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09458__S _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06110_ _01616_ _01582_ _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07090_ _02568_ _02569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07263__A2 _02729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11787__I _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12369__CLK clknet_leaf_184_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06041_ col_select_trans\[2\].data_sync col_select_trans\[3\].data_sync _01548_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_173_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11347__A1 _04417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09260__I0 _04265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_65_clock_I clknet_5_9_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09800_ _04615_ u2.mem\[38\]\[15\] _04633_ _04637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_82_clock clknet_5_8_0_clock clknet_leaf_82_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_113_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07992_ _03452_ _03453_ _03454_ _03455_ _03456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_119_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06774__A1 u2.mem\[168\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09193__S _04252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06943_ _02369_ _02422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_09731_ data_in_trans\[8\].data_sync _04591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09563__I1 u2.mem\[33\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09662_ _04545_ _00578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06874_ _01989_ row_select_trans\[5\].data_sync _02353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_67_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07723__B1 _03069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08613_ _03880_ _00194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_97_clock clknet_5_10_0_clock clknet_leaf_97_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_132_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09593_ _04505_ _00549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08544_ _03834_ _03840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09315__I1 u2.mem\[27\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11122__I1 u2.mem\[145\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08475_ _03714_ u2.mem\[8\]\[13\] _03792_ _03794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06829__A2 _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_20_clock clknet_5_2_0_clock clknet_leaf_20_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_126_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07426_ _02554_ _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09079__I0 _04132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08336__I _03704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13144__CLK clknet_leaf_41_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11898__S _05937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07357_ u2.mem\[57\]\[4\] _02671_ _02672_ u2.mem\[41\]\[4\] _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_13_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_342_clock_I clknet_5_7_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06308_ u2.mem\[171\]\[3\] _01610_ _01774_ u2.mem\[157\]\[3\] _01812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_35_clock clknet_5_3_0_clock clknet_leaf_35_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10633__I0 _05128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07254__A2 _02586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07288_ u2.mem\[60\]\[3\] _02542_ _02544_ u2.mem\[62\]\[3\] _02764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09027_ _04145_ u2.mem\[21\]\[5\] _04141_ _04146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13294__CLK clknet_leaf_383_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06239_ _01738_ _01739_ _01744_ _01745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_151_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10307__S _04944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11189__I1 u2.mem\[149\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07006__A2 _02400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08071__I data_in_trans\[10\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09251__I0 _04256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06765__A1 u2.mem\[153\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07962__B1 _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06765__B2 u2.mem\[160\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09929_ _04717_ _00673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11138__S _05462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12940_ _00819_ clknet_leaf_221_clock u2.mem\[51\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06517__A1 _01999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07714__B1 _03054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07415__I _02513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09831__S _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06459__C _01949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12871_ _00750_ clknet_leaf_134_clock u2.mem\[46\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09306__I1 u2.mem\[27\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11822_ _05893_ _01390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11753_ _05851_ _01363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10704_ _05124_ u2.mem\[60\]\[13\] _05189_ _05191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11684_ _05768_ _05808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07150__I _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13423_ _01302_ clknet_leaf_361_clock u2.mem\[174\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10635_ _04311_ _05071_ _05151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12511__CLK clknet_leaf_176_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11601__S _05747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10624__I0 _05119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13354_ _01233_ clknet_leaf_377_clock u2.mem\[162\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08182__S _03595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08442__A1 mem_address_trans\[2\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10566_ _03682_ _05108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07245__A2 _02537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12305_ _00184_ clknet_leaf_161_clock u2.mem\[11\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13285_ _01164_ clknet_leaf_381_clock u2.mem\[151\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10497_ _05065_ _00893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12236_ _00115_ clknet_leaf_226_clock u2.mem\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12661__CLK clknet_leaf_76_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12167_ _00046_ clknet_leaf_62_clock u2.mem\[2\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06756__A1 _02209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11118_ _05285_ _05443_ _05452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_7_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12098_ _01496_ clknet_leaf_246_clock u2.active_mem\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13017__CLK clknet_leaf_50_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11049_ _05390_ u2.mem\[140\]\[4\] _05403_ _05409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput7 data_in_a[0] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__07325__I _02464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_291_clock_I clknet_5_21_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12041__CLK clknet_2_2__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06590_ _02031_ _02037_ _02075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13167__CLK clknet_leaf_277_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08260_ _03646_ _00075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07484__A2 _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07060__I _02538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07211_ _02626_ _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08191_ _03579_ u2.mem\[2\]\[15\] _03600_ _03604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11511__S _05700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07142_ _02573_ _02574_ _02497_ _02450_ _02621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10615__I0 _05110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07236__A2 _02710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07073_ _02418_ _02510_ _02511_ _02430_ _02552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_12_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06995__A1 _02428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06024_ u2.driver_mem\[8\] _01512_ _01532_ _01519_ _01533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_114_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07975_ u2.mem\[37\]\[15\] _03295_ _03296_ u2.mem\[59\]\[15\] _03439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_60_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09714_ _04138_ _04578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06926_ _02404_ _02405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_28_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09645_ _04487_ u2.mem\[35\]\[10\] _04532_ _04535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06857_ _02309_ _02314_ _02323_ _02336_ _02337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_28_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09576_ _04494_ u2.mem\[33\]\[13\] _04492_ _04495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06788_ _02266_ _02267_ _02268_ _02269_ _02270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08527_ _03829_ _00159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08458_ _03784_ _00135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07475__A2 _02892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07409_ _02498_ _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_17_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06683__B1 _02148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08389_ _03741_ _00109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11421__S _05637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10420_ _03707_ _05020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10606__I0 _05101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07227__A2 _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12684__CLK clknet_leaf_216_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10351_ _04973_ _00839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09826__S _04649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13070_ _00949_ clknet_leaf_269_clock u2.mem\[59\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08730__S _03951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10282_ _04904_ u2.mem\[50\]\[8\] _04933_ _04934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_2_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12021_ net32 clknet_2_3__leaf_clock_a mem_address_trans\[8\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06738__A1 u2.mem\[151\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07935__B1 _02569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06738__B2 u2.mem\[158\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09527__I1 u2.mem\[32\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07950__A3 _03409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12064__CLK clknet_leaf_374_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07145__I _02623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12923_ _00802_ clknet_leaf_225_clock u2.mem\[50\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06984__I _02407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12854_ _00733_ clknet_leaf_86_clock u2.mem\[45\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09360__I _04118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_13_clock_I clknet_5_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06917__C _02395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11805_ _05883_ _01383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12785_ _00664_ clknet_leaf_336_clock u2.mem\[41\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10845__I0 _05198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11736_ _05841_ _01356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10470__A1 _03751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11667_ _05679_ _05798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13406_ _01285_ clknet_leaf_319_clock u2.mem\[171\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_174_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07218__A2 _02694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10618_ _05112_ u2.mem\[58\]\[8\] _05141_ _05142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11598_ _05754_ u2.mem\[174\]\[3\] _05748_ _05755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11270__I0 _05548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_238_clock_I clknet_5_25_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13337_ _01216_ clknet_leaf_4_clock u2.mem\[159\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10549_ _05096_ _00914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06977__A1 _02412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09215__I0 _04267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13268_ _01147_ clknet_leaf_384_clock u2.mem\[148\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11022__I0 _05392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12219_ _00098_ clknet_leaf_229_clock u2.mem\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13199_ _01078_ clknet_leaf_292_clock u2.mem\[136\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06729__A1 u2.mem\[176\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06729__B2 u2.mem\[189\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12407__CLK clknet_leaf_121_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09518__I1 u2.mem\[32\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07760_ _03211_ _03217_ _03222_ _03227_ _03228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_110_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06711_ u2.mem\[154\]\[1\] _02126_ _02129_ u2.mem\[148\]\[1\] _02127_ u2.mem\[162\]\[1\]
+ _02195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_49_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07691_ _02623_ _03161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07154__A1 _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12557__CLK clknet_leaf_202_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09430_ _04371_ u2.mem\[30\]\[6\] _04401_ _04404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06894__I _02372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06642_ _02064_ _02052_ _02127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_92_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09361_ _03903_ _04250_ _04357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06573_ _02056_ _02057_ _02058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_90_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08312_ _03685_ _00088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09292_ _04258_ u2.mem\[27\]\[3\] _04313_ _04317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07457__A2 _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08243_ _03550_ u2.mem\[4\]\[2\] _03634_ _03637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07209__A2 _02604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08174_ _03594_ _00041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07125_ _02603_ _02604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11040__I _05403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_161_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07056_ _02438_ _02472_ _02503_ _02534_ _02535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__09206__I0 _04260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11975__I _05970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11013__I0 _05386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06007_ u2.select_mem_row\[2\] u2.select_mem_col\[2\] _01515_ _01516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12087__CLK clknet_2_3__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input42_I row_select_a[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13332__CLK clknet_leaf_6_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09509__I1 u2.mem\[32\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07958_ u2.mem\[1\]\[15\] _03263_ _03264_ u2.mem\[7\]\[15\] _03422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_169_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06909_ _02365_ _02366_ _02367_ _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_99_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07889_ u2.mem\[37\]\[13\] _03295_ _03296_ u2.mem\[59\]\[13\] _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13482__CLK clknet_leaf_306_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09628_ _04525_ _00564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07696__A2 _03099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_187_clock_I clknet_5_30_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09559_ _04464_ _04483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12570_ _00449_ clknet_leaf_128_clock u2.mem\[27\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11521_ _05680_ u2.mem\[169\]\[5\] _05699_ _05706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_169_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06120__A2 _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11452_ _05635_ u2.mem\[165\]\[5\] _05654_ _05661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10403_ _05008_ _00856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11383_ _05589_ u2.mem\[161\]\[2\] _05616_ _05619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09556__S _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10334_ _04920_ u2.mem\[51\]\[15\] _04959_ _04963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06044__I col_select_trans\[4\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13122_ _01001_ clknet_leaf_257_clock u2.mem\[62\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13053_ _00932_ clknet_leaf_274_clock u2.mem\[58\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10265_ _04924_ _00802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07908__B1 _03352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11555__I1 u2.mem\[171\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12004_ _00016_ clknet_leaf_41_clock u2.mem\[0\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10196_ _04806_ u2.mem\[48\]\[10\] _04875_ _04878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11307__I1 u2.mem\[156\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12906_ _00785_ clknet_leaf_52_clock u2.mem\[48\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07687__A2 _03155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07603__I _02579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12837_ _00716_ clknet_leaf_88_clock u2.mem\[44\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12768_ _00647_ clknet_leaf_156_clock u2.mem\[40\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11719_ _05829_ u2.mem\[182\]\[1\] _05827_ _05830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_159_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13205__CLK clknet_leaf_292_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12699_ _00578_ clknet_leaf_227_clock u2.mem\[36\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput10 data_in_a[12] net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput21 data_in_a[8] net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput32 mem_address_a[8] net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_116_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11794__I1 u2.mem\[186\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07072__B1 _02550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08370__S _03727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13355__CLK clknet_leaf_370_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08930_ _04026_ u2.mem\[19\]\[5\] _04079_ _04081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10405__S _05002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08861_ _04038_ _00284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07812_ u2.mem\[58\]\[12\] _03277_ _03278_ u2.mem\[36\]\[12\] _03279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08792_ _03993_ _00260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07743_ _03207_ _03208_ _03209_ _03210_ _03211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_38_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07674_ u2.mem\[29\]\[9\] _03068_ _03069_ u2.mem\[11\]\[9\] _03144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10140__S _04841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06625_ u2.mem\[159\]\[0\] _02108_ _02109_ u2.mem\[149\]\[0\] _02110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09413_ _03581_ _03901_ _04393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__06350__A2 _01850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09344_ _04347_ _00458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06556_ _02036_ _02000_ _02041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08545__S _03840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09275_ _04306_ _00430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11482__I0 _05663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06487_ u2.mem\[193\]\[13\] _01917_ _01919_ u2.mem\[192\]\[13\] _01964_ _01975_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08226_ _03575_ u2.mem\[3\]\[13\] _03623_ _03625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08157_ _03584_ _03585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_107_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07108_ _02412_ _02587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__11785__I1 u2.mem\[186\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07602__A2 _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08280__S _03659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08088_ data_in_trans\[15\].data_sync _03534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07039_ _02517_ _02518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06956__A4 _02393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10050_ _04572_ _04788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10114__I _04819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10952_ _04138_ _05348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07669__A2 _03137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10673__A1 _04334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12102__CLK clknet_leaf_43_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10883_ _05303_ u2.mem\[130\]\[3\] _05297_ _05304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12622_ _00501_ clknet_leaf_201_clock u2.mem\[31\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08455__S _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06892__A3 _02344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12553_ _00432_ clknet_leaf_123_clock u2.mem\[26\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11504_ _05696_ _01269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12252__CLK clknet_leaf_266_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12484_ _00363_ clknet_leaf_107_clock u2.mem\[22\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11225__I0 _05505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11435_ _05651_ _01245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09286__S _04313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07054__B1 _02532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11366_ _05609_ _01218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08641__I1 u2.mem\[12\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06930__C _02408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10317_ _04953_ _00825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06801__B1 _02068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13105_ _00984_ clknet_leaf_329_clock u2.mem\[61\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10225__S _04896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11297_ _05565_ _01193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10248_ _04912_ _00797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13036_ _00915_ clknet_leaf_276_clock u2.mem\[57\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07357__B2 u2.mem\[41\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10024__I _04761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10179_ _04868_ _00772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11056__S _05413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06580__A2 _02028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07333__I _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10895__S _05310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06410_ u2.select_mem_row\[5\] u2.select_mem_col\[5\] _01515_ _01911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07390_ _02833_ _02844_ _02855_ _02864_ _02865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_34_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06341_ _01843_ _01844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06096__A1 _01566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09060_ _04170_ _04171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07293__B1 _02564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06272_ u2.mem\[167\]\[2\] _01621_ _01624_ u2.mem\[183\]\[2\] _01777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08011_ _03472_ _03473_ _01549_ _03474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_162_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12745__CLK clknet_leaf_44_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09196__S _04252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_135_clock_I clknet_5_15_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06399__A2 _01699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09962_ _04736_ _00687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08913_ _04048_ u2.mem\[18\]\[15\] _04066_ _04070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09893_ _04691_ u2.mem\[41\]\[4\] _04692_ _04693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08844_ _04026_ u2.mem\[17\]\[5\] _04024_ _04027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09723__I data_in_trans\[6\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06020__A1 u2.driver_mem\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08775_ _03980_ _00256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12125__CLK clknet_leaf_349_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08148__I0 _03577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07726_ _03191_ _03192_ _03193_ _03194_ _03195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08339__I data_in_trans\[12\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09896__I0 _04694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07657_ u2.mem\[14\]\[9\] _03125_ _03126_ u2.mem\[12\]\[9\] _03127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_380_clock clknet_5_0_0_clock clknet_leaf_380_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_40_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06608_ _02031_ _02070_ _02093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12275__CLK clknet_leaf_111_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07588_ _02541_ _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13520__CLK clknet_leaf_5_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09327_ _04254_ u2.mem\[28\]\[1\] _04336_ _04338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06539_ row_select_trans\[1\].data_sync _02024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_139_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08076__A2 _03516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07284__B1 _02508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08074__I data_in_trans\[11\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09258_ _04263_ u2.mem\[26\]\[5\] _04295_ _04297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07823__A2 _03271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11207__I0 _05508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08209_ _03615_ _00055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09189_ _04248_ _04249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_4_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11758__I1 u2.mem\[184\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11220_ _05518_ _01163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08623__I1 u2.mem\[12\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07587__A1 u2.mem\[61\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11151_ _05473_ _01139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10045__S _04784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07418__I _02520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10102_ _04823_ _00740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11082_ _05348_ _05430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07339__A1 _02806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10033_ _04761_ _04777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_103_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10194__I0 _04804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08000__A2 _03461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_333_clock clknet_5_18_0_clock clknet_leaf_333_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_75_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_337_clock_I clknet_5_18_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06562__A2 _02046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13050__CLK clknet_leaf_337_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11984_ _05227_ u2.mem\[194\]\[14\] _05971_ _05990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12618__CLK clknet_leaf_137_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10935_ _05334_ _05335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_348_clock clknet_5_7_0_clock clknet_leaf_348_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_95_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11604__S _05747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08185__S _03600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10866_ _05204_ u2.mem\[129\]\[4\] _05286_ _05292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12605_ _00484_ clknet_leaf_216_clock u2.mem\[30\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11446__I0 _05629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08067__A2 _03516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08311__I0 _03684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10797_ _05250_ _01008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12536_ _00415_ clknet_leaf_109_clock u2.mem\[25\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07102__B _02442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08913__S _04066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07814__A2 _03122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12467_ _00346_ clknet_leaf_108_clock u2.mem\[21\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11418_ _05641_ _01238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08614__I1 u2.mem\[12\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12398_ _00277_ clknet_leaf_191_clock u2.mem\[17\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07578__A1 u2.mem\[14\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11349_ _05583_ u2.mem\[159\]\[0\] _05598_ _05599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06786__C1 u2.mem\[144\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07328__I _02469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06250__A1 u2.mem\[159\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06250__B2 u2.mem\[149\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12148__CLK clknet_leaf_74_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13019_ _00898_ clknet_leaf_266_clock u2.mem\[56\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06890_ _02368_ _02369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10185__I0 _04795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11921__I1 u2.mem\[193\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06553__A2 _02037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08560_ _03823_ u2.mem\[10\]\[11\] _03845_ _03849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_63_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07063__I _02541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07511_ u2.mem\[3\]\[7\] _02803_ _02982_ _02983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13543__CLK clknet_leaf_40_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08491_ _03804_ _00148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07998__I _01547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07442_ _02595_ _02916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_61_clock_I clknet_5_9_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07373_ u2.mem\[17\]\[4\] _02846_ _02847_ u2.mem\[24\]\[4\] _02848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_17_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09112_ _04119_ u2.mem\[23\]\[0\] _04203_ _04204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06324_ _01820_ _01821_ _01822_ _01827_ _01828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__07266__B1 _02397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09919__S _04710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07805__A2 _03113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09043_ _04157_ _04158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06255_ u2.mem\[175\]\[1\] _01602_ _01632_ u2.mem\[188\]\[1\] _01761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_163_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06186_ _01563_ _01677_ _01580_ _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA_clkbuf_leaf_286_clock_I clknet_5_20_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_13_0_clock clknet_3_6_0_clock clknet_4_13_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_116_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07033__A3 _02382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09945_ _04696_ u2.mem\[42\]\[6\] _04724_ _04727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06792__A2 _02084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13073__CLK clknet_leaf_335_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09876_ _04680_ _00657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10176__I0 _04786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09453__I _04416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08827_ _04014_ _04015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_3305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10599__I _05130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07741__A1 u2.mem\[40\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06544__A2 _02028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07741__B2 u2.mem\[30\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08758_ _03920_ u2.mem\[15\]\[7\] _03967_ _03971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09869__I0 _04605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07709_ u2.mem\[58\]\[10\] _03044_ _03045_ u2.mem\[36\]\[10\] _03178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11676__I0 _05792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08689_ _03929_ u2.mem\[13\]\[11\] _03923_ _03930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09494__A1 _03982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12910__CLK clknet_leaf_202_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10720_ _05201_ _00980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11428__I0 _05623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10651_ _05160_ _00952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_166_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13370_ _01249_ clknet_leaf_375_clock u2.mem\[165\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10582_ _03703_ _05119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12321_ _00200_ clknet_leaf_167_clock u2.mem\[12\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10800__A1 _04416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12252_ _00131_ clknet_leaf_266_clock u2.mem\[8\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11203_ _05505_ u2.mem\[150\]\[1\] _05502_ _05506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12183_ _00062_ clknet_leaf_62_clock u2.mem\[3\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07148__I _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06232__A1 u2.mem\[144\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06232__B2 u2.mem\[182\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06052__I col_select_trans\[3\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11134_ _05461_ _05462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_95_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_272_clock clknet_5_23_0_clock clknet_leaf_272_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_27_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11065_ _05418_ _01108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10167__I0 _04817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10503__S _05066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12440__CLK clknet_leaf_119_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10016_ _04691_ u2.mem\[44\]\[4\] _04767_ _04768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11903__I1 _03524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13566__CLK clknet_leaf_13_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07732__A1 u2.mem\[5\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_287_clock clknet_5_20_0_clock clknet_leaf_287_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_45_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11967_ _05209_ u2.mem\[194\]\[6\] _05980_ _05981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08532__I0 _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12590__CLK clknet_leaf_201_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10095__A2 _04760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_1_clock clknet_5_0_0_clock clknet_leaf_1_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10918_ _05307_ u2.mem\[132\]\[5\] _05318_ _05325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07611__I _02598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11898_ u2.mem\[192\]\[9\] _03520_ _05937_ _05941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_210_clock clknet_5_28_0_clock clknet_leaf_210_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11419__I0 _05631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10849_ _05202_ u2.mem\[128\]\[3\] _05278_ _05282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07248__B1 _02676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08643__S _03894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13568_ _01447_ clknet_leaf_13_clock u2.mem\[194\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_173_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12519_ _00398_ clknet_leaf_125_clock u2.mem\[24\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07263__A3 _02734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13499_ _01378_ clknet_leaf_329_clock u2.mem\[186\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_225_clock clknet_5_29_0_clock clknet_leaf_225_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_12_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06040_ _01546_ _01547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07058__I _02536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09474__S _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07420__B1 _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_21_0_clock_I clknet_4_10_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07991_ u2.mem\[6\]\[15\] _02622_ _02624_ u2.mem\[47\]\[15\] _03455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07971__A1 _03431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06774__A2 _02093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09730_ _04590_ _00601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06942_ _02362_ _02421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__10158__I0 _04808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09273__I _04289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09661_ _04463_ u2.mem\[36\]\[0\] _04544_ _04545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06873_ _02340_ _02352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_94_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08612_ _03797_ u2.mem\[12\]\[0\] _03879_ _03880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12933__CLK clknet_leaf_63_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09592_ _04471_ u2.mem\[34\]\[3\] _04501_ _04505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08543_ _03839_ _00165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08523__I0 _03825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11244__S _05529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10330__I0 _04916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08474_ _03793_ _00142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07425_ _02552_ _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07239__B1 _02532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07356_ u2.mem\[37\]\[4\] _02829_ _02830_ u2.mem\[59\]\[4\] _02831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_104_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06307_ u2.mem\[167\]\[3\] _01749_ _01750_ u2.mem\[183\]\[3\] _01811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10882__I _04997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12313__CLK clknet_leaf_116_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07287_ u2.mem\[61\]\[3\] _02666_ _02667_ u2.mem\[63\]\[3\] _02763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10633__I1 u2.mem\[58\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09026_ _04144_ _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06238_ u2.mem\[147\]\[1\] _01676_ _01680_ u2.mem\[169\]\[1\] _01743_ _01744_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_156_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08352__I _03717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06169_ _01675_ _01676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07006__A3 _02392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09251__I1 u2.mem\[26\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06214__A1 _01678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12463__CLK clknet_leaf_174_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07411__B1 _02884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11419__S _05638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10323__S _04954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09928_ _04716_ u2.mem\[41\]\[15\] _04710_ _04717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10149__I0 _04799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06600__I _02084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09859_ _04660_ _04671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_3102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06517__A2 _02001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12870_ _00749_ clknet_leaf_85_clock u2.mem\[46\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08728__S _03951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09911__I _04598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07190__A2 _02666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11821_ _05874_ u2.mem\[188\]\[4\] _05887_ _05893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11154__S _05475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11752_ _05829_ u2.mem\[184\]\[1\] _05849_ _05851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10321__I0 _04907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07431__I _02549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10703_ _05190_ _00974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11683_ _05807_ _01337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13422_ _01301_ clknet_leaf_326_clock u2.mem\[173\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10634_ _05150_ _00945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06047__I _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10624__I1 u2.mem\[58\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13353_ _01232_ clknet_leaf_376_clock u2.mem\[162\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11821__I0 _05874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10565_ _05107_ _00919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12304_ _00183_ clknet_leaf_174_clock u2.mem\[11\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07650__B1 _03045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13284_ _01163_ clknet_leaf_370_clock u2.mem\[150\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12806__CLK clknet_leaf_87_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10496_ _05018_ u2.mem\[55\]\[11\] _05061_ _05065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12235_ _00114_ clknet_leaf_230_clock u2.mem\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06205__A1 _01566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12166_ _00045_ clknet_leaf_79_clock u2.mem\[2\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07953__A1 u2.mem\[32\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11117_ _05451_ _01127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12956__CLK clknet_leaf_197_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12097_ _01495_ clknet_leaf_246_clock u2.active_mem\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11048_ _05408_ _01101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07705__A1 _03170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput8 data_in_a[10] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_36_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_234_clock_I clknet_5_28_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09821__I _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12999_ _00878_ clknet_leaf_149_clock u2.mem\[54\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11064__S _05412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11265__A1 _04287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07469__B1 _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10312__I0 _04898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12336__CLK clknet_leaf_159_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07210_ _02684_ _02685_ _02686_ _02687_ _02688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_08190_ _03603_ _00048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_164_clock clknet_5_26_0_clock clknet_leaf_164_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07141_ u2.mem\[39\]\[0\] _02617_ _02619_ u2.mem\[48\]\[0\] _02620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10615__I1 u2.mem\[58\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06444__A1 _01844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12486__CLK clknet_leaf_107_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07072_ u2.mem\[57\]\[0\] _02548_ _02550_ u2.mem\[41\]\[0\] _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_173_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06995__A2 _02441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06023_ u2.driver_mem\[9\] _01517_ _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_160_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_179_clock clknet_5_27_0_clock clknet_leaf_179_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_114_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07944__A1 _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10143__S _04846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07974_ u2.mem\[60\]\[15\] _03292_ _03293_ u2.mem\[62\]\[15\] _03438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_102_clock clknet_5_10_0_clock clknet_leaf_102_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09932__S _04719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09713_ _04577_ _00597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06925_ _02352_ _02375_ _02404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_45_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11038__I _05275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09644_ _04534_ _00571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07960__B _02358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06856_ _02324_ _02329_ _02330_ _02335_ _02336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_56_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10551__I0 _05097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09731__I data_in_trans\[8\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13111__CLK clknet_leaf_39_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09575_ _04170_ _04494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06787_ u2.mem\[146\]\[3\] _02156_ _02122_ u2.mem\[173\]\[3\] _02269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_117_clock clknet_5_14_0_clock clknet_leaf_117_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08526_ _03828_ u2.mem\[9\]\[13\] _03826_ _03829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_24_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10303__I0 _04889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08347__I _03713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08457_ _03680_ u2.mem\[8\]\[5\] _03782_ _03784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_168_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13261__CLK clknet_leaf_286_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07408_ u2.mem\[50\]\[5\] _02880_ _02881_ u2.mem\[51\]\[5\] _02882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06683__A1 u2.mem\[170\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06683__B2 u2.mem\[156\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08388_ _03705_ u2.mem\[6\]\[11\] _03737_ _03741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12829__CLK clknet_leaf_203_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07339_ _02806_ _02807_ _02810_ _02813_ _02814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__10606__I1 u2.mem\[58\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09621__A1 _04072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08082__I data_in_trans\[13\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10350_ _04898_ u2.mem\[52\]\[5\] _04971_ _04973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07632__B1 _03020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09009_ _04130_ _04131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10281_ _04922_ _04933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_69_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12979__CLK clknet_leaf_30_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_183_clock_I clknet_5_27_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12020_ mem_address_trans\[7\].A clknet_leaf_315_clock mem_address_trans\[7\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07426__I _02554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09842__S _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10988__S _05364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08735__I0 _03934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12922_ _00801_ clknet_leaf_132_clock u2.mem\[49\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11495__A1 _04223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07699__B1 _03105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12853_ _00732_ clknet_leaf_84_clock u2.mem\[45\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06371__B1 _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11804_ _05872_ u2.mem\[187\]\[3\] _05879_ _05883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12784_ _00663_ clknet_leaf_336_clock u2.mem\[41\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07161__I _02425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09160__I0 _04140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11735_ _05825_ u2.mem\[183\]\[0\] _05840_ _05841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_81_clock clknet_5_8_0_clock clknet_leaf_81_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_14_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11612__S _05761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06674__A1 u2.mem\[146\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11666_ _05797_ _01330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_174_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13405_ _01284_ clknet_leaf_320_clock u2.mem\[171\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10617_ _05130_ _05141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_161_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10228__S _04896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11597_ _05673_ _05754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06426__A1 u2.mem\[194\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13336_ _01215_ clknet_leaf_14_clock u2.mem\[159\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08921__S _04074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_96_clock clknet_5_10_0_clock clknet_leaf_96_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11270__I1 u2.mem\[154\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10548_ _05093_ u2.mem\[57\]\[0\] _05095_ _05096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_170_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06977__A2 _02413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13267_ _01146_ clknet_leaf_384_clock u2.mem\[148\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10479_ _05055_ _00885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12218_ _00097_ clknet_leaf_54_clock u2.mem\[5\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13198_ _01077_ clknet_leaf_293_clock u2.mem\[136\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07926__A1 u2.mem\[49\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12149_ _00028_ clknet_leaf_74_clock u2.mem\[1\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07336__I _02486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06240__I _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08726__I0 _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06710_ _02191_ _02193_ _02194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07690_ _02621_ _03160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08368__S _03727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_34_clock clknet_5_3_0_clock clknet_leaf_34_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_92_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06641_ _02023_ _02125_ _02126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_168_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06362__B1 _01715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06901__A2 _02379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13284__CLK clknet_leaf_370_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09360_ _04118_ _04356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06572_ _02026_ _02036_ _02057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07071__I _02549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09151__I0 _04119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08311_ _03684_ u2.mem\[5\]\[6\] _03676_ _03685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_75_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09291_ _04316_ _00436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_49_clock clknet_5_7_0_clock clknet_leaf_49_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_127_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07457__A3 _02921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09199__S _04252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08242_ _03636_ _00067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07862__B1 _03161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08173_ _03561_ u2.mem\[2\]\[7\] _03590_ _03594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10138__S _04841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06417__A1 _01911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07124_ _02522_ _02523_ _02393_ _02506_ _02603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_118_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08831__S _04015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06415__I _01912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07055_ _02509_ _02519_ _02526_ _02533_ _02534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__09206__I1 u2.mem\[25\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06006_ _01502_ _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_114_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06150__I _01656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input35_I output_active_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07957_ u2.mem\[15\]\[15\] _03260_ _03261_ u2.mem\[13\]\[15\] _03421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_29_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08717__I0 _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12501__CLK clknet_leaf_119_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06908_ _02386_ _02387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_101_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07888_ u2.mem\[60\]\[13\] _03292_ _03293_ u2.mem\[62\]\[13\] _03354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_28_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09627_ _04469_ u2.mem\[35\]\[2\] _04522_ _04525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06839_ u2.mem\[166\]\[5\] _02097_ _02099_ u2.mem\[161\]\[5\] _02318_ _02319_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_43_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06353__B1 _01734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09558_ _04153_ _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08077__I _03488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08509_ _03798_ _03817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09489_ _04391_ u2.mem\[31\]\[15\] _04434_ _04438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11432__S _05647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11520_ _05705_ _01276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11451_ _05660_ _01252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10048__S _04784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09837__S _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10402_ _05007_ u2.mem\[53\]\[6\] _05002_ _05008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07605__B1 _03075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11252__I1 u2.mem\[153\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11382_ _05618_ _01225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13121_ _01000_ clknet_leaf_330_clock u2.mem\[62\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_152_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10333_ _04962_ _00832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12031__CLK clknet_2_3__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13157__CLK clknet_leaf_285_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13052_ _00931_ clknet_leaf_274_clock u2.mem\[58\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10264_ _04885_ u2.mem\[50\]\[0\] _04923_ _04924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_121_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07908__A1 _01973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12003_ _00015_ clknet_leaf_41_clock u2.mem\[0\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10195_ _04877_ _00779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07156__I _02435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06060__I _01566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08708__I0 _03907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09371__I _04135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12905_ _00784_ clknet_leaf_52_clock u2.mem\[48\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06344__B1 _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12836_ _00715_ clknet_leaf_88_clock u2.mem\[44\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12767_ _00646_ clknet_leaf_237_clock u2.mem\[40\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11342__S _05584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07844__B1 _03149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06647__B2 u2.mem\[152\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11718_ _03661_ _05829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12698_ _00577_ clknet_leaf_140_clock u2.mem\[35\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput11 data_in_a[13] net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_11649_ _05785_ _01325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput22 data_in_a[9] net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_156_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput33 mem_address_a[9] net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_7_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13319_ _01198_ clknet_leaf_312_clock u2.mem\[156\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09546__I _04464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12524__CLK clknet_leaf_198_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08860_ _04037_ u2.mem\[17\]\[10\] _04033_ _04038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07811_ _02489_ _03278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08791_ _03909_ u2.mem\[16\]\[2\] _03990_ _03993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11517__S _05700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07742_ u2.mem\[27\]\[11\] _03104_ _03105_ u2.mem\[35\]\[11\] _03210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09372__I0 _04364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07673_ u2.mem\[26\]\[9\] _03141_ _03142_ u2.mem\[10\]\[9\] _03143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_65_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09412_ _04392_ _00481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_131_clock_I clknet_5_15_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06624_ _02107_ _02037_ _02109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09343_ _04269_ u2.mem\[28\]\[8\] _04346_ _04347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06555_ u2.mem\[155\]\[0\] _02030_ _02035_ u2.mem\[174\]\[0\] u2.mem\[181\]\[0\]
+ _02039_ _02040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_34_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11252__S _05537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09274_ _04278_ u2.mem\[26\]\[12\] _04305_ _04306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11482__I1 u2.mem\[167\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06486_ u2.mem\[194\]\[13\] _01933_ _01974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08225_ _03624_ _00062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12054__CLK clknet_leaf_379_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08156_ _03479_ _03583_ _03584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07107_ _02585_ _02586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08087_ _01976_ _03526_ _03533_ _00015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_173_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06810__A1 u2.mem\[146\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07038_ _02395_ _02515_ _02516_ _02485_ _02517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__06810__B2 u2.mem\[186\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_56_clock_I clknet_5_12_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10745__I0 _05218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09392__S _04376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08989_ _04046_ u2.mem\[20\]\[14\] _04112_ _04115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07118__A2 _02594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09363__I0 _04356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06748__C _02230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10951_ _05347_ _01065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06326__B1 _01704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06877__A1 _02352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10882_ _04997_ _05303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12621_ _00500_ clknet_leaf_201_clock u2.mem\[31\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12552_ _00431_ clknet_leaf_122_clock u2.mem\[26\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08535__I _03834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11622__A1 _03486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06483__C _01964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11503_ _05674_ u2.mem\[168\]\[3\] _05692_ _05696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12483_ _00362_ clknet_leaf_119_clock u2.mem\[22\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_333_clock_I clknet_5_18_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11434_ _05631_ u2.mem\[164\]\[3\] _05647_ _05651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11225__I1 u2.mem\[151\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06055__I col_select_trans\[0\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12547__CLK clknet_leaf_110_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11365_ _05583_ u2.mem\[160\]\[0\] _05608_ _05609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06262__C1 u2.mem\[172\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13104_ _00983_ clknet_leaf_259_clock u2.mem\[61\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10316_ _04902_ u2.mem\[51\]\[7\] _04949_ _04953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06801__A1 u2.mem\[171\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11296_ _05556_ u2.mem\[155\]\[5\] _05558_ _05565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13035_ _00914_ clknet_leaf_264_clock u2.mem\[57\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08003__B1 _03459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10247_ _04911_ u2.mem\[49\]\[11\] _04905_ _04912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07357__A2 _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12697__CLK clknet_leaf_143_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10178_ _04788_ u2.mem\[48\]\[2\] _04865_ _04868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10241__S _04905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07614__I _02603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09354__I0 _04281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06317__C2 u2.mem\[193\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09106__I0 _04174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12819_ _00698_ clknet_leaf_113_clock u2.mem\[43\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10975__I _05275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12077__CLK clknet_2_1__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06340_ u2.mem\[0\]\[4\] _01843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08445__I _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13322__CLK clknet_leaf_322_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06393__C _01894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06271_ u2.mem\[178\]\[2\] _01617_ _01619_ u2.mem\[164\]\[2\] _01776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_8_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08010_ u2.active_mem\[0\] _03458_ _03459_ u2.active_mem\[1\] _03473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_159_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07045__A1 _02522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13472__CLK clknet_leaf_308_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07596__A2 _02908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09961_ _04712_ u2.mem\[42\]\[13\] _04734_ _04736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08912_ _04069_ _00304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09892_ _04682_ _04692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_97_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08843_ _03679_ _04026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06020__A2 _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08774_ _03936_ u2.mem\[15\]\[14\] _03977_ _03980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09345__I0 _04272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07725_ u2.mem\[28\]\[10\] _03074_ _03075_ u2.mem\[31\]\[10\] _03194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06308__B1 _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_282_clock_I clknet_5_22_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07656_ _02524_ _03126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08556__S _03845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06607_ _02091_ _02092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10885__I _05000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07587_ u2.mem\[61\]\[8\] _02899_ _02900_ u2.mem\[63\]\[8\] _03058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_94_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09326_ _04337_ _00450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06538_ _02022_ _02023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08355__I data_in_trans\[15\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_146_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09257_ _04296_ _00422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06469_ u2.mem\[193\]\[9\] _01960_ _01943_ u2.mem\[194\]\[9\] _01949_ _01961_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__07823__A3 _03280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08208_ _03557_ u2.mem\[3\]\[5\] _03613_ _03615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11207__I1 u2.mem\[150\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09188_ _03900_ _04247_ _04248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_120_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08139_ _03571_ _00029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09186__I _04118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07587__A2 _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11150_ _05472_ u2.mem\[146\]\[5\] _05461_ _05473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06795__B1 _02177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10101_ _04788_ u2.mem\[46\]\[2\] _04820_ _04823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11081_ _05429_ _01113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07339__A2 _02807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09914__I _04601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10032_ _04776_ _00717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10194__I1 u2.mem\[48\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06011__A2 _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07434__I _02566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09336__I0 _04263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06478__C _01964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10996__S _05373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11983_ _05989_ _01455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10934_ _04117_ _05334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13345__CLK clknet_leaf_3_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10865_ _05291_ _01035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12604_ _00483_ clknet_leaf_216_clock u2.mem\[30\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08265__I _03633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11446__I1 u2.mem\[165\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10796_ _05227_ u2.mem\[62\]\[14\] _05247_ _05250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12535_ _00414_ clknet_leaf_110_clock u2.mem\[25\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09297__S _04318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12466_ _00345_ clknet_leaf_174_clock u2.mem\[21\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11417_ _05629_ u2.mem\[163\]\[2\] _05638_ _05641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12397_ _00276_ clknet_leaf_193_clock u2.mem\[17\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07609__I _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07578__A2 _02892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11348_ _05597_ _05598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_152_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06786__B1 _02116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06786__C2 _02114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11279_ _05554_ u2.mem\[154\]\[4\] _05545_ _05555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13018_ _00897_ clknet_leaf_149_clock u2.mem\[55\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09327__I0 _04254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07750__A2 _03113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07510_ _02358_ _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08490_ _03803_ u2.mem\[9\]\[2\] _03799_ _03804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_81_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07502__A2 _02866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07441_ _02593_ _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12712__CLK clknet_leaf_146_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07372_ _02590_ _02847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08175__I _03584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09111_ _04202_ _04203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_17_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07266__A1 u2.mem\[32\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06323_ u2.mem\[166\]\[3\] _01757_ _01758_ u2.mem\[161\]\[3\] _01826_ _01827_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_104_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09042_ data_in_trans\[9\].data_sync _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06254_ u2.mem\[187\]\[1\] _01634_ _01637_ u2.mem\[192\]\[1\] _01760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_229_clock_I clknet_5_19_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06185_ _01691_ _01692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07569__A2 _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06423__I _01923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06777__B1 _02091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09944_ _04726_ _00679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09566__I0 _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09875_ _04615_ u2.mem\[40\]\[15\] _04676_ _04680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09191__A1 _04249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08826_ _04011_ _04013_ _04014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12242__CLK clknet_leaf_239_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13368__CLK clknet_leaf_372_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08757_ _03970_ _00248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11705__S _05818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07708_ u2.mem\[53\]\[10\] _03041_ _03042_ u2.mem\[56\]\[10\] _03177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11825__A1 _05411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08688_ _03704_ _03929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11676__I1 u2.mem\[179\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07639_ u2.mem\[1\]\[9\] _03030_ _03031_ u2.mem\[7\]\[9\] _03109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_81_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12392__CLK clknet_leaf_140_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11428__I1 u2.mem\[164\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08085__I data_in_trans\[14\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10650_ _05108_ u2.mem\[59\]\[6\] _05157_ _05160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09309_ _04326_ _00444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10581_ _05118_ _00924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12320_ _00199_ clknet_leaf_167_clock u2.mem\[12\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_167_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08813__I _03989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07009__A1 _02441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12251_ _00130_ clknet_leaf_228_clock u2.mem\[8\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11202_ _05504_ _05505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12182_ _00061_ clknet_leaf_76_clock u2.mem\[3\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07024__A4 _02502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06768__C2 u2.mem\[186\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11133_ _05295_ _05443_ _05461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11064_ _05390_ u2.mem\[141\]\[4\] _05412_ _05418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10015_ _04761_ _04767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_7_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07732__A2 _03155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11116__I0 _05432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11966_ _05971_ _05980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_3884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10917_ _05324_ _01054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_178_clock_I clknet_5_27_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11897_ _05940_ _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11419__I1 u2.mem\[163\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10848_ _05281_ _01028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07248__A1 u2.mem\[26\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13567_ _01446_ clknet_leaf_14_clock u2.mem\[194\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10779_ _05240_ _01000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12518_ _00397_ clknet_leaf_106_clock u2.mem\[24\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08723__I _03940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13498_ _01377_ clknet_leaf_329_clock u2.mem\[186\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_230_clock_I clknet_5_28_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12449_ _00328_ clknet_leaf_169_clock u2.mem\[20\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09796__I0 _04609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09755__S _04606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06243__I _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07015__A4 _02424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07420__B2 u2.mem\[12\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07990_ u2.mem\[8\]\[15\] _03326_ _03327_ u2.mem\[4\]\[15\] _03454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12265__CLK clknet_leaf_55_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06941_ _02419_ _02420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13510__CLK clknet_leaf_347_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11355__I0 _05591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09660_ _04543_ _04544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_clkbuf_5_25_0_clock_I clknet_4_12_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06872_ _02349_ _02350_ _02351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07184__B1 _02532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07074__I _02552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07723__A2 _03068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08611_ _03878_ _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09591_ _04504_ _00548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08542_ _03805_ u2.mem\[10\]\[3\] _03835_ _03839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07802__I _02469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08473_ _03709_ u2.mem\[8\]\[12\] _03792_ _03793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07424_ _02874_ _02879_ _02888_ _02897_ _02898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__08834__S _04015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07239__A1 u2.mem\[49\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07355_ _02538_ _02830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11260__S _05536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06306_ u2.mem\[178\]\[3\] _01746_ _01747_ u2.mem\[164\]\[3\] _01810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_332_clock clknet_5_18_0_clock clknet_leaf_332_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07286_ _02745_ _02751_ _02756_ _02761_ _02762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_163_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09025_ _04143_ _04144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06237_ _01740_ _01741_ _01742_ _01743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__13040__CLK clknet_leaf_336_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09665__S _04544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09787__I0 _04596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12608__CLK clknet_leaf_157_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06168_ _01612_ _01641_ _01675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10546__A1 _04249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_347_clock clknet_5_5_0_clock clknet_leaf_347_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06214__A2 _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10604__S _05131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06099_ _01578_ _01590_ _01599_ _01605_ _01606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__09464__I _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07962__A2 _02493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13190__CLK clknet_leaf_297_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09927_ _04614_ _04716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12758__CLK clknet_leaf_71_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09858_ _04670_ _00649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07175__B1 _02483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07714__A2 _03053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08809_ _03927_ u2.mem\[16\]\[10\] _04000_ _04003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_74_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09789_ _04599_ u2.mem\[38\]\[10\] _04628_ _04631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11820_ _05892_ _01389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11751_ _05850_ _01362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10702_ _05121_ u2.mem\[60\]\[12\] _05189_ _05190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11682_ _05798_ u2.mem\[179\]\[5\] _05800_ _05807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13421_ _01300_ clknet_leaf_312_clock u2.mem\[173\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12138__CLK clknet_leaf_38_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10633_ _05128_ u2.mem\[58\]\[15\] _05146_ _05150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13352_ _01231_ clknet_leaf_377_clock u2.mem\[162\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10564_ _05106_ u2.mem\[57\]\[5\] _05104_ _05107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11821__I1 u2.mem\[188\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06989__B1 _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12303_ _00182_ clknet_leaf_179_clock u2.mem\[11\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06491__C _01920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07650__A1 u2.mem\[58\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13283_ _01162_ clknet_leaf_384_clock u2.mem\[150\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10495_ _05064_ _00892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12288__CLK clknet_leaf_179_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09778__I0 _04583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12234_ _00113_ clknet_leaf_53_clock u2.mem\[6\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13533__CLK clknet_leaf_333_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06205__A2 _01586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12165_ _00044_ clknet_leaf_78_clock u2.mem\[2\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06998__I _02407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07402__B2 u2.mem\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08450__I0 _03667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10514__S _05073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09374__I _04139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06756__A3 _02223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11116_ _05432_ u2.mem\[144\]\[5\] _05444_ _05451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_123_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12096_ _01494_ clknet_leaf_246_clock u2.active_mem\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11047_ _05388_ u2.mem\[140\]\[3\] _05404_ _05408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08919__S _04074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07166__B1 _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09950__I0 _04700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput9 data_in_a[11] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_65_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11345__S _05584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12998_ _00877_ clknet_leaf_66_clock u2.mem\[54\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07622__I _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11949_ _05969_ _01441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08654__S _03905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06141__A1 _01606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07484__A4 _02956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13063__CLK clknet_leaf_47_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11080__S _05422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09549__I _04144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07140_ _02618_ _02619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_381_clock_I clknet_5_0_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06444__A2 _01938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07071_ _02549_ _02550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_161_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07069__I _02547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09769__I0 _04570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06022_ _01504_ _01529_ _01530_ _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_160_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06995__A3 _02381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11576__I0 _05711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07973_ u2.mem\[61\]\[15\] _02553_ _02555_ u2.mem\[63\]\[15\] _03437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_141_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09712_ _04576_ u2.mem\[37\]\[3\] _04567_ _04577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06924_ _02402_ _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07157__B1 _02634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10000__I0 _04714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09941__I0 _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09643_ _04485_ u2.mem\[35\]\[9\] _04532_ _04534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06855_ u2.mem\[169\]\[5\] _02141_ _02143_ u2.mem\[147\]\[5\] _02334_ _02335_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_23_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09574_ _04493_ _00542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06786_ u2.mem\[185\]\[3\] _02120_ _02116_ u2.mem\[182\]\[3\] u2.mem\[144\]\[3\]
+ _02114_ _02268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08525_ _03713_ _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13406__CLK clknet_leaf_319_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08456_ _03783_ _00134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06132__A1 _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07407_ _02494_ _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08387_ _03740_ _00108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_271_clock clknet_5_23_0_clock clknet_leaf_271_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06683__A2 _02146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10067__I0 _04799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07338_ u2.mem\[58\]\[4\] _02811_ _02812_ u2.mem\[36\]\[4\] _02813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08363__I _03726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12430__CLK clknet_leaf_191_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13556__CLK clknet_leaf_14_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07632__A1 u2.mem\[32\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08680__I0 _03922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07269_ _02741_ _02742_ _02743_ _02744_ _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09395__S _04376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09008_ data_in_trans\[2\].data_sync _04130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06840__C1 _02092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_286_clock clknet_5_20_0_clock clknet_leaf_286_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_151_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10280_ _04932_ _00809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_126_clock_I clknet_5_15_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10334__S _04959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06199__B2 u2.mem\[194\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07935__A2 _02567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_0_clock clknet_5_0_0_clock clknet_leaf_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_104_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11319__I0 _05550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10133__I _04840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09932__I0 _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08735__I1 u2.mem\[14\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12921_ _00800_ clknet_leaf_132_clock u2.mem\[49\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07699__A1 u2.mem\[27\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11495__A2 _05690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_224_clock clknet_5_29_0_clock clknet_leaf_224_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12852_ _00731_ clknet_leaf_84_clock u2.mem\[45\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06371__A1 u2.mem\[147\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07442__I _02595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11803_ _05882_ _01382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12783_ _00662_ clknet_leaf_249_clock u2.mem\[41\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13086__CLK clknet_leaf_274_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09160__I1 u2.mem\[24\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11734_ _05839_ _05840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_239_clock clknet_5_25_0_clock clknet_leaf_239_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_41_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11665_ _05796_ u2.mem\[178\]\[4\] _05787_ _05797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06674__A2 _02156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10058__I0 _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13404_ _01283_ clknet_leaf_326_clock u2.mem\[170\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10616_ _05140_ _00937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11596_ _05753_ _01304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13335_ _01214_ clknet_leaf_14_clock u2.mem\[159\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06426__A2 _01924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10547_ _05094_ _05095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_143_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12923__CLK clknet_leaf_225_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06831__C1 u2.mem\[181\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13266_ _01145_ clknet_leaf_310_clock u2.mem\[147\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10478_ _04998_ u2.mem\[55\]\[3\] _05051_ _05055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12217_ _00096_ clknet_leaf_44_clock u2.mem\[5\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10244__S _04905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13197_ _01076_ clknet_leaf_294_clock u2.mem\[136\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12148_ _00027_ clknet_leaf_74_clock u2.mem\[1\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06521__I _02005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12079_ net13 clknet_2_0__leaf_clock_a data_in_trans\[15\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_328_clock_I clknet_5_17_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12303__CLK clknet_leaf_179_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06640_ _02027_ _02032_ _02125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07352__I _02543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06571_ _02005_ _02056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10297__I0 _04920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08310_ _03683_ _03684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09290_ _04256_ u2.mem\[27\]\[2\] _04313_ _04316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08384__S _03737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12453__CLK clknet_leaf_90_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06114__A1 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08241_ _03548_ u2.mem\[4\]\[1\] _03634_ _03636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06665__A2 _02077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08172_ _03593_ _00040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07123_ u2.mem\[52\]\[0\] _02599_ _02601_ u2.mem\[21\]\[0\] _02602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07054_ u2.mem\[49\]\[0\] _02528_ _02532_ u2.mem\[46\]\[0\] _02533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11549__I0 _05713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06005_ _01504_ _01509_ _01513_ _01514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_115_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10154__S _04851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09943__S _04724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10221__I0 _04893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07956_ _03416_ _03417_ _03418_ _03419_ _03420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_112_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06907_ _02364_ _02371_ _02353_ _02386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA_input28_I mem_address_a[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10888__I _05004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07887_ u2.mem\[61\]\[13\] _02553_ _02555_ u2.mem\[63\]\[13\] _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09626_ _04524_ _00563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06838_ _02315_ _02316_ _02317_ _02318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06353__A1 u2.mem\[193\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07550__B1 _03020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06353__B2 u2.mem\[177\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09557_ _04481_ _00537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06769_ u2.mem\[164\]\[3\] _02051_ _02054_ u2.mem\[178\]\[3\] _02251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08508_ _03691_ _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10288__I0 _04911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_52_clock_I clknet_5_13_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09488_ _04437_ _00512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07302__B1 _02690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08439_ _03722_ u2.mem\[7\]\[15\] _03768_ _03772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_168_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12946__CLK clknet_leaf_151_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09189__I _04248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11450_ _05633_ u2.mem\[165\]\[4\] _05654_ _05660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11788__I0 _05872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10401_ _03682_ _05007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06408__A2 _01887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11381_ _05587_ u2.mem\[161\]\[1\] _05616_ _05618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09917__I _04604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13120_ _00999_ clknet_leaf_258_clock u2.mem\[62\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10332_ _04918_ u2.mem\[51\]\[14\] _04959_ _04962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_277_clock_I clknet_5_23_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13051_ _00930_ clknet_leaf_264_clock u2.mem\[58\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10263_ _04922_ _04923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10212__I0 _04885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12002_ _00014_ clknet_leaf_41_clock u2.mem\[0\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06341__I _01843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10194_ _04804_ u2.mem\[48\]\[9\] _04875_ _04877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_79_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12326__CLK clknet_leaf_93_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11960__I0 _05911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_163_clock clknet_5_26_0_clock clknet_leaf_163_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_93_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12904_ _00783_ clknet_leaf_52_clock u2.mem\[48\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06344__A1 u2.mem\[172\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07172__I _02498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06344__B2 u2.mem\[150\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12835_ _00714_ clknet_leaf_113_clock u2.mem\[44\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10279__I0 _04902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_178_clock clknet_5_27_0_clock clknet_leaf_178_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12766_ _00645_ clknet_leaf_219_clock u2.mem\[40\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06647__A2 _02129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11717_ _05828_ _01350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12697_ _00576_ clknet_leaf_143_clock u2.mem\[35\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07121__B _02474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11648_ _05758_ u2.mem\[177\]\[5\] _05778_ _05785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08932__S _04079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_101_clock clknet_5_10_0_clock clknet_leaf_101_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xinput12 data_in_a[14] net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__11779__I0 _05864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput23 inverter_select_a net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput34 mem_write_n_a net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_11579_ _05742_ _01298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13318_ _01197_ clknet_leaf_318_clock u2.mem\[156\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07072__A2 _02548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13101__CLK clknet_leaf_281_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_116_clock clknet_5_14_0_clock clknet_leaf_116_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_171_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13249_ _01128_ clknet_leaf_302_clock u2.mem\[145\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10203__I0 _04813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09763__S _04606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06251__I _01592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08021__A1 mem_address_trans\[2\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07810_ _02486_ _03277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13251__CLK clknet_leaf_307_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08790_ _03992_ _00259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09562__I _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12819__CLK clknet_leaf_113_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07741_ u2.mem\[40\]\[11\] _03022_ _03023_ u2.mem\[30\]\[11\] _03209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11703__I0 _05790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07672_ _02568_ _03142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_168_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07082__I _02448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09411_ _04391_ u2.mem\[29\]\[15\] _04385_ _04392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_19_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06623_ _02107_ _02104_ _02108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12969__CLK clknet_leaf_127_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09342_ _04335_ _04346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_146_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06554_ _02038_ _02039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08906__I _04050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07810__I _02486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09273_ _04289_ _04305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_166_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10149__S _04846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06485_ u2.mem\[0\]\[13\] _01973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11332__I _05504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09938__S _04719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08224_ _03572_ u2.mem\[3\]\[12\] _03623_ _03624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10690__I0 _05110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11993__CLK clknet_leaf_334_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08155_ _03582_ _03583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_146_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07599__B1 _03069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07106_ _02447_ _02449_ _02454_ _02575_ _02585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_88_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08086_ _03532_ _03528_ _03533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_162_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12349__CLK clknet_leaf_208_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07037_ _02480_ _02516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__06271__B1 _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06810__A2 _02156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08012__A1 _01613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10745__I1 u2.mem\[61\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11942__I0 _05222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_80_clock clknet_5_8_0_clock clknet_leaf_80_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_103_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12499__CLK clknet_leaf_119_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08988_ _04114_ _00335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07771__B1 _03149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07939_ _03400_ _03401_ _03402_ _03403_ _03404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_28_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10411__I _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10950_ _05346_ u2.mem\[134\]\[3\] _05337_ _05347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08088__I data_in_trans\[15\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06326__B2 u2.mem\[194\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_95_clock clknet_5_10_0_clock clknet_leaf_95_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09609_ _04514_ _00556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06877__A2 _02353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10881_ _05302_ _01040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12620_ _00499_ clknet_leaf_201_clock u2.mem\[31\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12551_ _00430_ clknet_leaf_123_clock u2.mem\[26\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06629__A2 _02001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11502_ _05695_ _01268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09848__S _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10681__I0 _05101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12482_ _00361_ clknet_leaf_172_clock u2.mem\[22\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08752__S _03967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13124__CLK clknet_leaf_20_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11433_ _05650_ _01244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_33_clock clknet_5_3_0_clock clknet_leaf_33_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_153_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07054__A2 _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11364_ _05607_ _05608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_152_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10315_ _04952_ _00824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13103_ _00982_ clknet_leaf_259_clock u2.mem\[61\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06801__A2 _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13274__CLK clknet_leaf_7_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11295_ _05564_ _01192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13034_ _00913_ clknet_leaf_51_clock u2.mem\[56\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10246_ _04601_ _04911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08003__A1 u2.active_mem\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08003__B2 u2.active_mem\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_48_clock clknet_5_7_0_clock clknet_leaf_48_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_26_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11933__I0 _05213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11618__S _05760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08199__S _03608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10177_ _04867_ _00771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06565__A1 _02031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07762__B1 _03060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07116__B _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06317__A1 u2.mem\[158\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07514__B1 _02884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06317__B2 u2.mem\[151\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12818_ _00697_ clknet_leaf_166_clock u2.mem\[43\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07630__I _02435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12749_ _00628_ clknet_leaf_223_clock u2.mem\[39\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06270_ u2.mem\[171\]\[2\] _01611_ _01774_ u2.mem\[157\]\[2\] _01775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07293__A2 _02559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07832__A4 _03298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10991__I _05372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11377__A1 _05285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09290__I0 _04256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09960_ _04735_ _00686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08911_ _04046_ u2.mem\[18\]\[14\] _04066_ _04069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12641__CLK clknet_leaf_157_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09891_ _04578_ _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11924__I0 _05913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08842_ _04025_ _00278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07753__B1 _03045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08773_ _03979_ _00255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11327__I _05499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07724_ u2.mem\[9\]\[10\] _03071_ _03072_ u2.mem\[25\]\[10\] _03193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_2_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12791__CLK clknet_leaf_339_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08837__S _04015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06308__A1 u2.mem\[171\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07505__B1 _02872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06308__B2 u2.mem\[157\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_225_clock_I clknet_5_29_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07655_ _02520_ _03125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06859__A2 row_select_trans\[4\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06606_ _02080_ _01999_ _02091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07586_ _03026_ _03038_ _03047_ _03056_ _03057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__12021__CLK clknet_2_3__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09325_ _04246_ u2.mem\[28\]\[0\] _04336_ _04337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06537_ _02004_ _01997_ _02022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09256_ _04260_ u2.mem\[26\]\[4\] _04295_ _04296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07284__A2 _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06468_ _01927_ _01960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07823__A4 _03289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08207_ _03614_ _00054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13297__CLK clknet_leaf_382_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09187_ _03748_ _03774_ _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_06399_ u2.mem\[154\]\[5\] _01699_ _01701_ u2.mem\[162\]\[5\] _01900_ _01901_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_135_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05995__I _01503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10415__I0 _05016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08138_ _03570_ u2.mem\[1\]\[11\] _03564_ _03571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08069_ _03520_ _03518_ _03521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_150_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06795__A1 u2.mem\[149\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10100_ _04822_ _00739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06795__B2 u2.mem\[175\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11080_ _05428_ u2.mem\[142\]\[3\] _05422_ _05429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11915__I0 _05903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10031_ _04707_ u2.mem\[44\]\[11\] _04772_ _04776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07339__A3 _02810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07744__B1 _03028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11237__I _05528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09336__I1 u2.mem\[28\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08747__S _03962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11982_ _05225_ u2.mem\[194\]\[13\] _05985_ _05989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10933_ _05333_ _01061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11173__S _05484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10864_ _05202_ u2.mem\[129\]\[3\] _05287_ _05291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12603_ _00482_ clknet_leaf_214_clock u2.mem\[30\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08847__I0 _04028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10795_ _05249_ _01007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12514__CLK clknet_leaf_174_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11901__S _05942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12534_ _00413_ clknet_leaf_101_clock u2.mem\[25\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06066__I col_select_trans\[0\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06483__B1 _01943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12465_ _00344_ clknet_leaf_173_clock u2.mem\[21\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_173_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11700__I _05817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11416_ _05640_ _01237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12396_ _00275_ clknet_leaf_193_clock u2.mem\[17\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_165_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12664__CLK clknet_leaf_141_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11347_ _04417_ _05566_ _05597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_154_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06786__A1 u2.mem\[185\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07983__B1 _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06786__B2 u2.mem\[182\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_174_clock_I clknet_5_27_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11278_ _05513_ _05554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10229_ _04899_ _00791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13017_ _00896_ clknet_leaf_50_clock u2.mem\[55\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07735__B1 _03161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold1 output_active_hold\[0\] net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_66_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08657__S _03905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12044__CLK clknet_leaf_315_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11083__S _05421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07440_ _02910_ _02911_ _02912_ _02913_ _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__10893__I0 _05294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07360__I _02558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07371_ _02585_ _02846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_99_clock_I clknet_5_10_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09110_ _03751_ _04122_ _04202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06322_ _01823_ _01824_ _01825_ _01826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_148_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07266__A2 _02385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06069__A3 _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09041_ _04156_ _00346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06474__B1 _01948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06253_ u2.mem\[166\]\[1\] _01757_ _01758_ u2.mem\[161\]\[1\] _01759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07018__A2 _02391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06184_ _01566_ _01616_ _01691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06777__A1 u2.mem\[145\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06777__B2 u2.mem\[177\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09943_ _04694_ u2.mem\[42\]\[5\] _04724_ _04726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11258__S _05537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09874_ _04679_ _00656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08825_ _04012_ _04013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08567__S _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08756_ _03918_ u2.mem\[15\]\[6\] _03967_ _03970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_85_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input10_I data_in_a[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09750__I _04566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_376_clock_I clknet_5_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07707_ u2.mem\[54\]\[10\] _03116_ _03117_ u2.mem\[55\]\[10\] _03176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08687_ _03928_ _00220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07638_ u2.mem\[15\]\[9\] _03027_ _03028_ u2.mem\[13\]\[9\] _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07569_ u2.mem\[54\]\[8\] _02883_ _02884_ u2.mem\[55\]\[8\] _03040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_107_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09398__S _04376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09308_ _04274_ u2.mem\[27\]\[10\] _04323_ _04326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_16_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10580_ _05117_ u2.mem\[57\]\[10\] _05113_ _05118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12687__CLK clknet_leaf_157_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_7_0_clock clknet_3_3_0_clock clknet_4_7_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_10_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09239_ _04284_ _00416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12250_ _00129_ clknet_leaf_56_clock u2.mem\[7\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07009__A2 _02381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06614__I _02098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11201_ _03495_ _05504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12181_ _00060_ clknet_leaf_78_clock u2.mem\[3\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06768__A1 u2.mem\[169\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06768__B2 u2.mem\[147\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11132_ _05334_ _05460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09006__I0 _04128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11063_ _05417_ _01107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12067__CLK clknet_2_1__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07717__B1 _03133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10014_ _04766_ _00709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13312__CLK clknet_leaf_363_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06940__A1 _02412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09660__I _04543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11116__I1 u2.mem\[144\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11965_ _05979_ _01447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13462__CLK clknet_leaf_360_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08276__I _03655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10916_ _05305_ u2.mem\[132\]\[4\] _05318_ _05324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11896_ u2.mem\[192\]\[8\] _03517_ _05937_ _05940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10847_ _05200_ u2.mem\[128\]\[2\] _05278_ _05281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10627__I0 _05121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07248__A2 _02675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13566_ _01445_ clknet_leaf_13_clock u2.mem\[194\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10778_ _05209_ u2.mem\[62\]\[6\] _05237_ _05240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06456__B1 _01947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12517_ _00396_ clknet_leaf_107_clock u2.mem\[24\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10247__S _04905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13497_ _01376_ clknet_leaf_329_clock u2.mem\[186\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06524__I row_select_trans\[3\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12448_ _00327_ clknet_leaf_168_clock u2.mem\[20\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12379_ _00258_ clknet_leaf_233_clock u2.mem\[16\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06759__A1 u2.mem\[187\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06759__B2 u2.mem\[192\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07420__A2 _02892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06940_ _02412_ _02413_ _02417_ _02418_ _02419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_84_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07708__B1 _03042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input2_I col_select_a[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07355__I _02538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09771__S _04618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11355__I1 u2.mem\[159\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06871_ col_select_trans\[5\].data_sync _01986_ _02350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_94_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07184__A1 u2.mem\[49\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11806__S _05878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08610_ _03629_ _03541_ _03877_ _03878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_132_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09590_ _04469_ u2.mem\[34\]\[2\] _04501_ _04504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08541_ _03838_ _00164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_29_0_clock_I clknet_4_14_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08472_ _03776_ _03792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_35_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10866__I0 _05204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07090__I _02568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07423_ _02891_ _02894_ _02895_ _02896_ _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_126_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11541__S _05708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10618__I0 _05112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07354_ _02536_ _02829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07239__A2 _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09011__S _04124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06305_ _01808_ _01809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_149_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07285_ _02757_ _02758_ _02759_ _02760_ _02761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_149_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09024_ data_in_trans\[5\].data_sync _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_164_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06236_ u2.mem\[146\]\[1\] _01692_ _01694_ u2.mem\[186\]\[1\] _01742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06434__I _01923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11043__I0 _05384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06167_ u2.mem\[144\]\[0\] _01671_ _01673_ u2.mem\[182\]\[0\] _01674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_144_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09745__I _04601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06214__A3 _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13335__CLK clknet_leaf_14_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07411__A2 _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06098_ u2.mem\[175\]\[0\] _01602_ _01604_ u2.mem\[159\]\[0\] _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_172_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09926_ _04715_ _00672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09681__S _04554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09857_ _04589_ u2.mem\[40\]\[7\] _04666_ _04670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11716__S _05827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08808_ _04002_ _00267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10620__S _05141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06922__A1 _02390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09788_ _04630_ _00619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08739_ _03938_ u2.mem\[14\]\[15\] _03956_ _03960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_122_clock_I clknet_5_14_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11750_ _05825_ u2.mem\[184\]\[0\] _05849_ _05850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06609__I _02093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10701_ _05173_ _05189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_144_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11681_ _05806_ _01336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13420_ _01299_ clknet_leaf_313_clock u2.mem\[173\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10609__I0 _05103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10632_ _05149_ _00944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11282__I0 _05556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13351_ _01230_ clknet_leaf_377_clock u2.mem\[162\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10563_ _05004_ _05106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06989__B2 u2.mem\[33\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12302_ _00181_ clknet_leaf_200_clock u2.mem\[11\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07650__A2 _03044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10494_ _05016_ u2.mem\[55\]\[10\] _05061_ _05064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13282_ _01161_ clknet_leaf_383_clock u2.mem\[150\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11034__I0 _05390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12233_ _00112_ clknet_leaf_54_clock u2.mem\[6\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12164_ _00043_ clknet_leaf_78_clock u2.mem\[2\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_47_clock_I clknet_5_7_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11115_ _05450_ _01126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06756__A4 _02238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12702__CLK clknet_leaf_224_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12095_ _01493_ clknet_leaf_338_clock u2.active_mem\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11046_ _05407_ _01100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07166__B2 u2.mem\[33\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11626__S _05771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10530__S _05083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06913__A1 _02348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12997_ _00876_ clknet_leaf_66_clock u2.mem\[54\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11425__I _05605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07124__B _02393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07469__A2 _02880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06519__I row_select_trans\[5\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11948_ _05229_ u2.mem\[193\]\[15\] _05965_ _05969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13208__CLK clknet_leaf_297_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06141__A2 _01629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11879_ _05930_ _01410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11273__I0 _05550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13549_ _01428_ clknet_leaf_9_clock u2.mem\[193\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_146_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_324_clock_I clknet_5_16_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07070_ _02395_ _02529_ _02530_ _02546_ _02549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__12232__CLK clknet_leaf_55_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13358__CLK clknet_leaf_372_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07641__A2 _03036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06021_ u2.driver_mem\[10\] _01512_ _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09769__I1 u2.mem\[38\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09565__I _04160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12382__CLK clknet_leaf_232_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07944__A3 _03407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07972_ _03420_ _03425_ _03430_ _03435_ _03436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_102_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07085__I _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09711_ _04575_ _04576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06923_ _02363_ _02370_ _02374_ _02401_ _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__07157__B2 u2.mem\[34\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09642_ _04533_ _00570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06854_ _02331_ _02332_ _02333_ _02334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06904__A1 _02377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09006__S _04124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09573_ _04491_ u2.mem\[33\]\[12\] _04492_ _04493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06785_ u2.mem\[179\]\[3\] _02151_ _02153_ u2.mem\[191\]\[3\] _02267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_97_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11335__I _05507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06380__A2 _01880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08524_ _03827_ _00158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08455_ _03675_ u2.mem\[8\]\[4\] _03782_ _03783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06132__A2 _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07406_ _02492_ _02880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08386_ _03701_ u2.mem\[6\]\[10\] _03737_ _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07880__A2 _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07337_ _02489_ _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11070__I _05421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09209__I0 _04263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07268_ u2.mem\[27\]\[3\] _02638_ _02639_ u2.mem\[35\]\[3\] _02744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_87_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06164__I _01670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07632__A2 _03019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09007_ _04129_ _00339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11016__I0 _05388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06219_ _01545_ _01555_ _01725_ _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06840__B1 _02078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07199_ u2.mem\[26\]\[1\] _02675_ _02676_ u2.mem\[10\]\[1\] _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12725__CLK clknet_leaf_24_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10615__S _05136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07396__A1 u2.mem\[40\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07396__B2 u2.mem\[30\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10414__I _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11319__I1 u2.mem\[157\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12875__CLK clknet_leaf_228_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09909_ _04703_ u2.mem\[41\]\[9\] _04701_ _04704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_24_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11446__S _05655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12920_ _00799_ clknet_leaf_133_clock u2.mem\[49\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07699__A2 _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12851_ _00730_ clknet_leaf_86_clock u2.mem\[45\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12105__CLK clknet_leaf_25_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06371__A2 _01675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_273_clock_I clknet_5_23_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11802_ _05870_ u2.mem\[187\]\[2\] _05879_ _05882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12782_ _00661_ clknet_leaf_268_clock u2.mem\[41\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11733_ _05354_ _05808_ _05839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12255__CLK clknet_leaf_241_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09448__I0 _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11664_ _05676_ _05796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10058__I1 u2.mem\[45\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13403_ _01282_ clknet_leaf_326_clock u2.mem\[170\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10615_ _05110_ u2.mem\[58\]\[7\] _05136_ _05140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09073__A1 _04180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11595_ _05752_ u2.mem\[174\]\[2\] _05748_ _05753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09586__S _04501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06074__I _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13334_ _01213_ clknet_leaf_3_clock u2.mem\[159\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08490__S _03799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_4_0_clock clknet_0_clock clknet_3_4_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_10546_ _04249_ _05071_ _05094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11007__I0 _05380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06831__B1 _02034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10525__S _05078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06831__C2 _02038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13265_ _01144_ clknet_leaf_311_clock u2.mem\[147\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10477_ _05054_ _00884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12216_ _00095_ clknet_leaf_54_clock u2.mem\[5\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13196_ _01075_ clknet_leaf_293_clock u2.mem\[136\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12147_ _00026_ clknet_leaf_75_clock u2.mem\[1\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_173_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07139__A1 _02506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12078_ data_in_trans\[14\].A clknet_leaf_349_clock data_in_trans\[14\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08187__I0 _03575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10260__S _04914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11029_ _05397_ _01093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_331_clock clknet_5_18_0_clock clknet_leaf_331_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_20_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06570_ u2.mem\[164\]\[0\] _02051_ _02054_ u2.mem\[178\]\[0\] _02055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_3490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_346_clock clknet_5_5_0_clock clknet_leaf_346_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06114__A2 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08240_ _03635_ _00066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09439__I0 _04380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07862__A2 _03160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13180__CLK clknet_leaf_279_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08171_ _03559_ u2.mem\[2\]\[6\] _03590_ _03593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12748__CLK clknet_leaf_223_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07122_ _02600_ _02601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09496__S _04443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07053_ _02531_ _02532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10435__S _05030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07808__I _02482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11549__I1 u2.mem\[171\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06004_ u2.driver_mem\[2\] _01512_ _01513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06712__I _02136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10221__I1 u2.mem\[49\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_6_0_clock clknet_4_3_0_clock clknet_5_6_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_07955_ u2.mem\[27\]\[15\] _02420_ _02426_ u2.mem\[35\]\[15\] _03419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08178__I0 _03566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12128__CLK clknet_leaf_37_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06906_ _02384_ _02385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08878__A1 _03583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07886_ _03336_ _03341_ _03346_ _03351_ _03352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_29_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09625_ _04467_ u2.mem\[35\]\[1\] _04522_ _04524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_16_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06837_ u2.mem\[159\]\[5\] _02108_ _02109_ u2.mem\[149\]\[5\] _02317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_83_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07550__A1 u2.mem\[32\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12278__CLK clknet_leaf_99_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09556_ _04480_ u2.mem\[33\]\[7\] _04474_ _04481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08575__S _03856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06768_ u2.mem\[169\]\[3\] _02142_ _02144_ u2.mem\[147\]\[3\] _02158_ u2.mem\[186\]\[3\]
+ _02250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_70_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13523__CLK clknet_leaf_13_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08507_ _03815_ _00153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09487_ _04389_ u2.mem\[31\]\[14\] _04434_ _04437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06699_ _02180_ _02181_ _02182_ _02183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07302__B2 u2.mem\[38\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08438_ _03771_ _00128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08369_ _03730_ _00100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11788__I1 u2.mem\[186\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07066__B1 _02544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10400_ _05006_ _00855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11380_ _05617_ _01224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07605__A2 _03074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06408__A3 _01896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10331_ _04961_ _00831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10345__S _04966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10262_ _03583_ _04863_ _04922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06622__I _02022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13050_ _00929_ clknet_leaf_337_clock u2.mem\[57\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12001_ _00013_ clknet_leaf_41_clock u2.mem\[0\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10193_ _04876_ _00778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06041__A1 col_select_trans\[2\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11960__I1 u2.mem\[194\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08169__I0 _03557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13053__CLK clknet_leaf_274_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10080__S _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07453__I _02621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06497__C _01911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12903_ _00782_ clknet_leaf_147_clock u2.mem\[48\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12834_ _00713_ clknet_leaf_164_clock u2.mem\[44\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12765_ _00644_ clknet_leaf_219_clock u2.mem\[40\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08284__I _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11716_ _05825_ u2.mem\[182\]\[0\] _05827_ _05828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07844__A2 _03148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12696_ _00575_ clknet_leaf_140_clock u2.mem\[35\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11647_ _05784_ _01324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput13 data_in_a[15] net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_30_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput24 mem_address_a[0] net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_122_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput35 output_active_a net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_11578_ _05713_ u2.mem\[173\]\[2\] _05739_ _05742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13317_ _01196_ clknet_leaf_317_clock u2.mem\[156\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10529_ _05084_ _00906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06280__A1 u2.mem\[187\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13248_ _01127_ clknet_leaf_308_clock u2.mem\[144\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06280__B2 u2.mem\[192\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11400__I0 _05629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13179_ _01058_ clknet_leaf_279_clock u2.mem\[133\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08021__A2 mem_address_trans\[3\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_270_clock clknet_5_23_0_clock clknet_leaf_270_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11086__S _05421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07740_ u2.mem\[32\]\[11\] _03019_ _03020_ u2.mem\[2\]\[11\] _03208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07363__I _02571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12420__CLK clknet_leaf_102_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11703__I1 u2.mem\[181\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13546__CLK clknet_leaf_38_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07671_ _02566_ _03141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07532__A1 u2.mem\[28\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09410_ _04176_ _04391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06622_ _02022_ _02107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08395__S _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_285_clock clknet_5_20_0_clock clknet_leaf_285_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_80_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09341_ _04345_ _00457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06553_ _01999_ _02037_ _02038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_169_clock_I clknet_5_26_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12570__CLK clknet_leaf_128_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08332__I0 _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06099__A1 _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09272_ _04304_ _00429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06484_ _01969_ _01970_ _01971_ _01972_ _01461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_21_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08223_ _03607_ _03623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__11219__I0 _05517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08154_ _03484_ _03581_ _03582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07105_ _02565_ _02570_ _02578_ _02583_ _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_119_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_221_clock_I clknet_5_29_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08085_ data_in_trans\[14\].data_sync _03532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_223_clock clknet_5_23_0_clock clknet_leaf_223_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_66_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09954__S _04729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07036_ _02478_ _02515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__06271__B2 u2.mem\[164\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13076__CLK clknet_leaf_26_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_29_0_clock clknet_4_14_0_clock clknet_5_29_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08012__A2 _03471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09753__I data_in_trans\[13\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input40_I row_select_a[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06023__A1 u2.driver_mem\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08987_ _04044_ u2.mem\[20\]\[13\] _04112_ _04114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_238_clock clknet_5_25_0_clock clknet_leaf_238_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_87_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07938_ u2.mem\[28\]\[14\] _03307_ _03308_ u2.mem\[31\]\[14\] _03403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_5_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09899__I0 _04696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07273__I _02358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07869_ u2.mem\[27\]\[13\] _02420_ _02426_ u2.mem\[35\]\[13\] _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_95_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06326__A2 _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09608_ _04487_ u2.mem\[34\]\[10\] _04511_ _04514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10880_ _05301_ u2.mem\[130\]\[2\] _05297_ _05302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11458__I0 _05663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09539_ _04131_ _04469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12550_ _00429_ clknet_leaf_100_clock u2.mem\[26\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07287__B1 _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10130__I0 _04817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11501_ _05671_ u2.mem\[168\]\[2\] _05692_ _05695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12481_ _00360_ clknet_leaf_172_clock u2.mem\[22\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11432_ _05629_ u2.mem\[164\]\[2\] _05647_ _05650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11630__I0 _05754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13419__CLK clknet_leaf_318_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11363_ _03486_ _05606_ _05607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__07448__I _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09864__S _04671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06262__A1 u2.mem\[189\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13102_ _00981_ clknet_leaf_282_clock u2.mem\[61\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10314_ _04900_ u2.mem\[51\]\[6\] _04949_ _04952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06262__B2 u2.mem\[176\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11294_ _05554_ u2.mem\[155\]\[4\] _05558_ _05564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13033_ _00912_ clknet_leaf_51_clock u2.mem\[56\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12006__D mem_address_trans\[0\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10245_ _04910_ _00796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08003__A2 _03458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06014__A1 u2.driver_mem\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12443__CLK clknet_leaf_185_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11933__I1 u2.mem\[193\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10176_ _04786_ u2.mem\[48\]\[1\] _04865_ _04867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13569__CLK clknet_leaf_12_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06565__A2 _02041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07762__B2 u2.mem\[62\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08279__I _03658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11697__I0 _05798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12593__CLK clknet_leaf_161_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11634__S _05770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09104__S _04197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12817_ _00696_ clknet_leaf_167_clock u2.mem\[43\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_170_clock_I clknet_5_26_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07132__B _02488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07278__B1 _02483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10121__I0 _04808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12748_ _00627_ clknet_leaf_223_clock u2.mem\[39\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08943__S _04084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12679_ _00558_ clknet_leaf_142_clock u2.mem\[34\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08742__I _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_156_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13099__CLK clknet_leaf_260_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09290__I1 u2.mem\[27\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06253__A1 u2.mem\[166\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07450__B1 _02923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06253__B2 u2.mem\[161\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08910_ _04068_ _00303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_30_0_clock clknet_4_15_0_clock clknet_5_30_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_98_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10713__S _05196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09890_ _04690_ _00661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07202__B1 _02582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_95_clock_I clknet_5_10_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11924__I1 u2.mem\[193\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08841_ _04023_ u2.mem\[17\]\[4\] _04024_ _04025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07348__A4 _02822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07753__A1 u2.mem\[58\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12936__CLK clknet_leaf_147_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08772_ _03934_ u2.mem\[15\]\[13\] _03977_ _03979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07093__I _02571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07723_ u2.mem\[29\]\[10\] _03068_ _03069_ u2.mem\[11\]\[10\] _03192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07505__A1 u2.mem\[27\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06308__A2 _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07654_ u2.mem\[44\]\[9\] _03122_ _03123_ u2.mem\[42\]\[9\] _03124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_168_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06605_ u2.mem\[151\]\[0\] _02085_ _02087_ u2.mem\[158\]\[0\] u2.mem\[193\]\[0\]
+ _02089_ _02090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07585_ _03048_ _03049_ _03052_ _03055_ _03056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_94_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09324_ _04335_ _04336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06536_ u2.mem\[176\]\[0\] _02003_ _02013_ u2.mem\[172\]\[0\] _02020_ u2.mem\[189\]\[0\]
+ _02021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__10112__I0 _04799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09255_ _04289_ _04295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__12316__CLK clknet_leaf_185_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06467_ u2.mem\[192\]\[9\] _01929_ _01959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09748__I data_in_trans\[12\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08206_ _03554_ u2.mem\[3\]\[4\] _03613_ _03614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06492__A1 _01976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09186_ _04118_ _04246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06398_ _01897_ _01898_ _01899_ _01900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xclkbuf_leaf_162_clock clknet_5_26_0_clock clknet_leaf_162_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_120_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_372_clock_I clknet_5_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11612__I0 _05752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08137_ _03524_ _03570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12466__CLK clknet_leaf_174_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08068_ data_in_trans\[9\].data_sync _03520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11719__S _05827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07019_ _02473_ _02422_ _02423_ _02497_ _02498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_103_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_177_clock clknet_5_27_0_clock clknet_leaf_177_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_153_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10030_ _04775_ _00716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11915__I1 u2.mem\[193\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08099__I mem_address_trans\[0\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_3_0_clock clknet_3_1_0_clock clknet_4_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xclkbuf_leaf_100_clock clknet_5_10_0_clock clknet_leaf_100_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_75_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11981_ _05988_ _01454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10932_ _05307_ u2.mem\[133\]\[5\] _05326_ _05333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08827__I _04014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10863_ _05290_ _01034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_115_clock clknet_5_14_0_clock clknet_leaf_115_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12602_ _00481_ clknet_leaf_116_clock u2.mem\[29\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10103__I0 _04790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08763__S _03972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10794_ _05225_ u2.mem\[62\]\[13\] _05247_ _05249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_169_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12533_ _00412_ clknet_leaf_104_clock u2.mem\[25\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11851__I0 _05911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13241__CLK clknet_leaf_288_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09658__I _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08562__I _03834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07680__B1 _03149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12464_ _00343_ clknet_leaf_174_clock u2.mem\[21\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12809__CLK clknet_leaf_129_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11415_ _05627_ u2.mem\[163\]\[1\] _05638_ _05640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12395_ _00274_ clknet_leaf_190_clock u2.mem\[17\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07178__I _02513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06235__B2 u2.mem\[179\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07432__B1 _02905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11346_ _05596_ _01211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13391__CLK clknet_leaf_367_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_117_clock_I clknet_5_14_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06786__A2 _02120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12959__CLK clknet_leaf_168_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11277_ _05553_ _01185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13016_ _00895_ clknet_leaf_339_clock u2.mem\[55\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10228_ _04898_ u2.mem\[49\]\[5\] _04896_ _04899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07735__A1 u2.mem\[6\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10159_ _04855_ _00765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold2 output_active_trans.data_sync net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XANTENNA__10590__I0 _05124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_169_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12339__CLK clknet_leaf_93_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09769__S _04618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07370_ u2.mem\[23\]\[4\] _02682_ _02683_ u2.mem\[22\]\[4\] _02845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06321_ u2.mem\[159\]\[3\] _01604_ _01595_ u2.mem\[149\]\[3\] _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11842__I0 _05903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09568__I _04163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09040_ _04154_ u2.mem\[21\]\[8\] _04155_ _04156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06252_ _01598_ _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06474__A1 u2.mem\[193\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12489__CLK clknet_leaf_125_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08472__I _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06183_ u2.mem\[170\]\[0\] _01687_ _01689_ u2.mem\[156\]\[0\] _01690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10507__I _04862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07018__A3 _02392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07088__I _02566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_94_clock clknet_5_10_0_clock clknet_leaf_94_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_102_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06777__A2 _02081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07974__A1 u2.mem\[60\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09942_ _04725_ _00678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07816__I _02527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09873_ _04612_ u2.mem\[40\]\[14\] _04676_ _04679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11338__I _05510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08774__I0 _03936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08824_ _03482_ _03539_ _03544_ _04012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_161_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13114__CLK clknet_leaf_45_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08755_ _03969_ _00247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_319_clock_I clknet_5_16_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08526__I0 _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07706_ u2.mem\[50\]\[10\] _03113_ _03114_ u2.mem\[51\]\[10\] _03175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08647__I _03655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08686_ _03927_ u2.mem\[13\]\[10\] _03923_ _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_32_clock clknet_5_3_0_clock clknet_leaf_32_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07551__I _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07637_ _03101_ _03102_ _03103_ _03106_ _03107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11073__I _05339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13264__CLK clknet_leaf_287_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09679__S _04554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07568_ u2.mem\[50\]\[8\] _02880_ _02881_ u2.mem\[51\]\[8\] _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_80_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09307_ _04325_ _00443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_47_clock clknet_5_7_0_clock clknet_leaf_47_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_10_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06519_ row_select_trans\[5\].data_sync _02004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11833__I0 _05872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10618__S _05141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07499_ _02968_ _02969_ _02970_ _02971_ _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_139_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06465__A1 _01954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09238_ _04283_ u2.mem\[25\]\[14\] _04279_ _04284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09169_ _04154_ u2.mem\[24\]\[8\] _04236_ _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07009__A3 _02382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10417__I _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11200_ _05503_ _01158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12180_ _00059_ clknet_leaf_78_clock u2.mem\[3\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07965__A1 u2.mem\[58\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_3_0_clock_I clknet_4_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07965__B2 u2.mem\[36\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11131_ _05459_ _01133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06630__I _02114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11062_ _05388_ u2.mem\[141\]\[3\] _05413_ _05417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07717__A1 u2.mem\[61\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08765__I0 _03927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10013_ _04689_ u2.mem\[44\]\[3\] _04762_ _04766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08758__S _03967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06940__A2 _02413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11964_ _05915_ u2.mem\[194\]\[5\] _05975_ _05979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10915_ _05323_ _01053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11895_ _05939_ _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_43_clock_I clknet_5_6_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06077__I col_select_trans\[2\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08493__S _03799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10846_ _05280_ _01027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12631__CLK clknet_leaf_113_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13565_ _01444_ clknet_leaf_13_clock u2.mem\[194\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10627__I1 u2.mem\[58\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10528__S _05083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10777_ _05239_ _00999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09388__I _04357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06456__A1 _01945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12516_ _00395_ clknet_leaf_107_clock u2.mem\[24\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08292__I _03501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13496_ _01375_ clknet_leaf_259_clock u2.mem\[186\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12447_ _00326_ clknet_leaf_168_clock u2.mem\[20\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10327__I _04943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12781__CLK clknet_leaf_268_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12378_ _00257_ clknet_leaf_60_clock u2.mem\[15\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_268_clock_I clknet_5_22_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11359__S _05597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11329_ _05584_ _05585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_4_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12011__CLK clknet_2_1__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13137__CLK clknet_leaf_335_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08756__I0 _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06870_ _02348_ _02349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_95_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07184__A2 _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_320_clock_I clknet_5_16_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13287__CLK clknet_leaf_382_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11094__S _05435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08540_ _03803_ u2.mem\[10\]\[2\] _03835_ _03838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_48_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07371__I _02585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08471_ _03791_ _00141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07422_ u2.mem\[43\]\[5\] _02820_ _02821_ u2.mem\[20\]\[5\] _02896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_165_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07892__B1 _02569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11815__I0 _05868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07353_ u2.mem\[60\]\[4\] _02826_ _02827_ u2.mem\[62\]\[4\] _02828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10618__I1 u2.mem\[58\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11621__I _05768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06304_ u2.mem\[0\]\[3\] _01808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11440__A1 _04120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06715__I _02134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07284_ u2.mem\[43\]\[3\] _02505_ _02508_ u2.mem\[20\]\[3\] _02760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09023_ _04142_ _00342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10237__I _04886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06235_ u2.mem\[191\]\[1\] _01682_ _01684_ u2.mem\[179\]\[1\] _01741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_156_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06166_ _01672_ _01673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07947__B2 u2.mem\[4\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06097_ _01603_ _01604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07546__I _02360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09925_ _04714_ u2.mem\[41\]\[14\] _04710_ _04715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11068__I _05334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08747__I0 _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09856_ _04669_ _00648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10901__S _05309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10554__I0 _05099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09761__I data_in_trans\[15\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07175__A2 _02476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08807_ _03925_ u2.mem\[16\]\[9\] _04000_ _04002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_150_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09787_ _04596_ u2.mem\[38\]\[9\] _04628_ _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06383__B1 _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06999_ _02368_ _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06922__A2 _02400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08738_ _03959_ _00240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08669_ _03679_ _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10700_ _05188_ _00973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06686__A1 u2.mem\[146\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11680_ _05796_ u2.mem\[179\]\[4\] _05800_ _05806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06686__B2 u2.mem\[186\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09202__S _04252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11806__I0 _05874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10609__I1 u2.mem\[58\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10631_ _05126_ u2.mem\[58\]\[14\] _05146_ _05149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11531__I _05670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06438__A1 u2.mem\[192\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07230__B _02359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13350_ _01229_ clknet_leaf_7_clock u2.mem\[161\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10562_ _05105_ _00918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12301_ _00180_ clknet_leaf_205_clock u2.mem\[11\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06989__A2 _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13281_ _01160_ clknet_leaf_384_clock u2.mem\[150\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10493_ _05063_ _00891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12034__CLK clknet_leaf_301_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12232_ _00111_ clknet_leaf_55_clock u2.mem\[6\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08840__I _04014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11179__S _05483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12163_ _00042_ clknet_leaf_79_clock u2.mem\[2\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06071__C1 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06610__A1 u2.mem\[177\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11114_ _05430_ u2.mem\[144\]\[4\] _05444_ _05450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06610__B2 u2.mem\[168\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12094_ _01486_ clknet_leaf_337_clock u2.active_mem\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12184__CLK clknet_leaf_62_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11907__S _05942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11045_ _05386_ u2.mem\[140\]\[2\] _05404_ _05407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12014__D mem_address_trans\[4\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07166__A2 _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06913__A2 _02350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_0_0_clock clknet_0_clock clknet_3_0_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_76_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08287__I _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12996_ _00875_ clknet_leaf_65_clock u2.mem\[54\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11947_ _05968_ _01440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07124__C _02506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11642__S _05779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11670__A1 _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11878_ u2.mem\[192\]\[0\] _03491_ _05929_ _05930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09112__S _04203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06141__A3 _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_158_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10829_ u2.mem\[63\]\[12\] _03527_ _05268_ _05269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11273__I1 u2.mem\[154\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06535__I _02019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13548_ _01427_ clknet_leaf_37_clock u2.mem\[193\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10057__I _04783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13479_ _01358_ clknet_leaf_304_clock u2.mem\[183\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_173_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06020_ u2.driver_mem\[11\] _01508_ _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12527__CLK clknet_leaf_189_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07366__I _02579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09782__S _04623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07944__A4 _03408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07971_ _03431_ _03432_ _03433_ _03434_ _03435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_113_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09710_ _04134_ _04575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11817__S _05888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06922_ _02390_ _02400_ _02382_ _02401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_45_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07157__A2 _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09581__I _04176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09641_ _04482_ u2.mem\[35\]\[8\] _04532_ _04533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06853_ u2.mem\[146\]\[5\] _02155_ _02157_ u2.mem\[186\]\[5\] _02333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_7_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06365__B1 _01672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06904__A2 _02381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09572_ _04464_ _04492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06784_ u2.mem\[170\]\[3\] _02146_ _02148_ u2.mem\[156\]\[3\] _02266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_83_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08523_ _03825_ u2.mem\[9\]\[12\] _03826_ _03827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_24_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08454_ _03776_ _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07865__B1 _03290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09022__S _04141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07405_ _02875_ _02876_ _02877_ _02878_ _02879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_23_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08385_ _03739_ _00107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_5_2_0_clock clknet_4_1_0_clock clknet_5_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_143_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12057__CLK clknet_2_0__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07336_ _02486_ _02811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13302__CLK clknet_leaf_5_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07267_ u2.mem\[40\]\[3\] _02403_ _02410_ u2.mem\[30\]\[3\] _02743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09209__I1 u2.mem\[25\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09006_ _04128_ u2.mem\[21\]\[1\] _04124_ _04129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06218_ _01648_ _01669_ _01724_ _01725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__06840__A1 u2.mem\[165\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06840__B2 u2.mem\[163\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07198_ _02568_ _02676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_145_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06149_ _01561_ _01564_ _01596_ _01656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_117_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06180__I _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09908_ _04595_ _04703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10631__S _05146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09839_ _04440_ _04659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06356__B1 _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10430__I _03720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12850_ _00729_ clknet_leaf_154_clock u2.mem\[45\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09145__I0 _04177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_216_clock_I clknet_5_29_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11801_ _05881_ _01381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12781_ _00660_ clknet_leaf_268_clock u2.mem\[41\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11732_ _05838_ _01355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_159_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_5_11_0_clock_I clknet_4_5_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11663_ _05795_ _01329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09448__I1 u2.mem\[30\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13402_ _01281_ clknet_leaf_312_clock u2.mem\[170\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10614_ _05139_ _00936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11594_ _05670_ _05752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07084__A1 _02560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13333_ _01212_ clknet_leaf_3_clock u2.mem\[159\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10545_ _04986_ _05093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10806__S _05253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06831__A1 u2.mem\[155\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13264_ _01143_ clknet_leaf_287_clock u2.mem\[147\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10476_ _04995_ u2.mem\[55\]\[2\] _05051_ _05054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12215_ _00094_ clknet_leaf_43_clock u2.mem\[5\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13195_ _01074_ clknet_leaf_294_clock u2.mem\[136\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06090__I _01596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12146_ _00025_ clknet_leaf_238_clock u2.mem\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_150_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12077_ net12 clknet_2_1__leaf_clock_a data_in_trans\[14\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07139__A2 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11028_ _05384_ u2.mem\[139\]\[1\] _05395_ _05397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11191__I0 _05470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09136__I0 _04164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12979_ _00858_ clknet_leaf_30_clock u2.mem\[53\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13325__CLK clknet_leaf_323_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09439__I1 u2.mem\[30\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08170_ _03592_ _00039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07121_ _02560_ _02561_ _02474_ _02589_ _02600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__07075__A1 _02463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_146_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10716__S _05196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13475__CLK clknet_leaf_311_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07052_ _02395_ _02529_ _02530_ _02406_ _02531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_106_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06003_ _01511_ _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07096__I _02347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07954_ u2.mem\[40\]\[15\] _03255_ _03256_ u2.mem\[30\]\[15\] _03418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_64_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06905_ _02363_ _02370_ _02374_ _02383_ _02384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_101_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07885_ _03347_ _03348_ _03349_ _03350_ _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_56_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10250__I _04886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09624_ _04523_ _00562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07045__B _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06836_ u2.mem\[188\]\[5\] _02103_ _02105_ u2.mem\[175\]\[5\] _02316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09127__I0 _04151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07550__A2 _03019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09555_ _04150_ _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06767_ u2.mem\[148\]\[3\] _02129_ _02131_ u2.mem\[152\]\[3\] _02248_ _02249_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_102_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11282__S _05545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08506_ _03814_ u2.mem\[9\]\[7\] _03808_ _03815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_19_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09486_ _04436_ _00511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06698_ u2.mem\[184\]\[1\] _02071_ _01993_ _02182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07302__A2 _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_5_25_0_clock clknet_4_12_0_clock clknet_5_25_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08437_ _03718_ u2.mem\[7\]\[14\] _03768_ _03771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_93_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06175__I _01681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08591__S _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08368_ _03667_ u2.mem\[6\]\[2\] _03727_ _03730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_109_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07319_ _02444_ _02794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08299_ _03674_ _03675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06408__A4 _01909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10996__I0 _05343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10330_ _04916_ u2.mem\[51\]\[13\] _04959_ _04961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08390__I _03726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10261_ _04921_ _00801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10748__I0 _05220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07369__A2 _02837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12000_ _00012_ clknet_leaf_19_clock u2.mem\[0\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10192_ _04801_ u2.mem\[48\]\[8\] _04875_ _04876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06041__A2 col_select_trans\[3\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10361__S _04976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12992__CLK clknet_leaf_256_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09366__I0 _04360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11173__I0 _05466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10160__I _04840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12902_ _00781_ clknet_leaf_71_clock u2.mem\[48\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09118__I0 _04136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12222__CLK clknet_leaf_225_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_367_clock_I clknet_5_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13348__CLK clknet_leaf_14_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12833_ _00712_ clknet_5_26_0_clock u2.mem\[44\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12764_ _00643_ clknet_leaf_220_clock u2.mem\[40\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11715_ _05826_ _05827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_72_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12372__CLK clknet_leaf_79_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12695_ _00574_ clknet_leaf_140_clock u2.mem\[35\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13498__CLK clknet_leaf_329_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11646_ _05756_ u2.mem\[177\]\[4\] _05778_ _05784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07057__A1 _02455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput14 data_in_a[1] net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_174_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput25 mem_address_a[1] net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_35_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11577_ _05741_ _01297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput36 row_col_select_a net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_168_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13316_ _01195_ clknet_leaf_316_clock u2.mem\[156\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06804__A1 _02277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10528_ _05011_ u2.mem\[56\]\[8\] _05083_ _05084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08006__B1 _03459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13247_ _01126_ clknet_leaf_288_clock u2.mem\[144\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10459_ _05018_ u2.mem\[54\]\[11\] _05040_ _05044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10739__I0 _05213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11400__I1 u2.mem\[162\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13178_ _01057_ clknet_leaf_293_clock u2.mem\[133\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11367__S _05608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12129_ _01470_ clknet_leaf_36_clock u2.driver_mem\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11164__I0 _05472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11166__I _05442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10070__I _04783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07670_ _03134_ _03135_ _03136_ _03139_ _03140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_42_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06621_ u2.mem\[188\]\[0\] _02103_ _02105_ u2.mem\[175\]\[0\] _02106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12715__CLK clknet_leaf_268_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09340_ _04267_ u2.mem\[28\]\[7\] _04341_ _04345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06552_ _02017_ _02036_ _02037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08332__I1 u2.mem\[5\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09271_ _04276_ u2.mem\[26\]\[11\] _04300_ _04304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_91_clock_I clknet_5_10_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06483_ u2.mem\[193\]\[12\] _01960_ _01943_ u2.mem\[194\]\[12\] _01964_ _01972_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_142_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08222_ _03622_ _00061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11219__I1 u2.mem\[150\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12865__CLK clknet_leaf_154_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07048__A1 _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08153_ _03542_ _03543_ _03581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_53_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10446__S _05035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10978__I0 _05335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07599__A2 _03068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07104_ u2.mem\[28\]\[0\] _02580_ _02582_ u2.mem\[31\]\[0\] _02583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07819__I _02504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08084_ _01973_ _03526_ _03531_ _00014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_49_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07035_ _02513_ _02514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06271__A2 _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07220__A1 _02674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06023__A2 _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08986_ _04113_ _00334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12245__CLK clknet_leaf_74_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input33_I mem_address_a[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07771__A2 _03148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07937_ u2.mem\[9\]\[14\] _03304_ _03305_ u2.mem\[25\]\[14\] _03402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_151_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11076__I _05342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12112__D _01475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07868_ u2.mem\[40\]\[13\] _03255_ _03256_ u2.mem\[30\]\[13\] _03334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_17_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07523__A2 _02984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09607_ _04513_ _00555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06819_ u2.mem\[154\]\[4\] _02225_ _02226_ u2.mem\[162\]\[4\] _02299_ _02300_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_56_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12395__CLK clknet_leaf_190_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07799_ _02464_ _03266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09538_ _04468_ _00531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_169_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09520__I0 _04382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09469_ _04371_ u2.mem\[31\]\[6\] _04424_ _04427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07287__B2 u2.mem\[63\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11500_ _05694_ _01267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12480_ _00359_ clknet_leaf_176_clock u2.mem\[22\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11431_ _05649_ _01243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_330_clock clknet_5_18_0_clock clknet_leaf_330_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_165_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11362_ _05605_ _05606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_164_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11630__I1 u2.mem\[176\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06798__B1 _02061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13101_ _00980_ clknet_leaf_281_clock u2.mem\[61\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10313_ _04951_ _00823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13020__CLK clknet_leaf_272_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06262__A2 _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11293_ _05563_ _01191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13032_ _00911_ clknet_leaf_48_clock u2.mem\[56\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10244_ _04909_ u2.mem\[49\]\[10\] _04905_ _04910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11394__I0 _05623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11187__S _05492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_345_clock clknet_5_7_0_clock clknet_leaf_345_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06014__A2 _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10175_ _04866_ _00770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13170__CLK clknet_leaf_283_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07762__A2 _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09880__S _04683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12738__CLK clknet_leaf_248_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11915__S _05950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11697__I1 u2.mem\[180\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07514__A2 _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_113_clock_I clknet_5_11_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12816_ _00695_ clknet_leaf_167_clock u2.mem\[43\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09511__I0 _04373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12888__CLK clknet_leaf_57_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07132__C _02562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12747_ _00626_ clknet_leaf_271_clock u2.mem\[39\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12678_ _00557_ clknet_leaf_63_clock u2.mem\[34\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12118__CLK clknet_leaf_349_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11629_ _05774_ _01316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10266__S _04923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12268__CLK clknet_leaf_194_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_171_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10337__A1 _04095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13513__CLK clknet_leaf_354_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11385__I0 _05591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_38_clock_I clknet_5_6_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08840_ _04014_ _04024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_112_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08250__I0 _03557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07374__I _02598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07753__A2 _03044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08771_ _03978_ _00254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07722_ u2.mem\[26\]\[10\] _03141_ _03142_ u2.mem\[10\]\[10\] _03191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07505__A2 _02871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07653_ _02517_ _03123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06604_ _02088_ _02089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07584_ u2.mem\[43\]\[8\] _03053_ _03054_ u2.mem\[20\]\[8\] _03055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_168_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09323_ _04011_ _04334_ _04335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09502__I0 _04364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06535_ _02019_ _02020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11560__S _05731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09254_ _04294_ _00421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06466_ net49 _01958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_107_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08205_ _03607_ _03613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_21_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09185_ _04245_ _00401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13043__CLK clknet_leaf_31_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06397_ u2.mem\[152\]\[5\] _01712_ _01714_ u2.mem\[148\]\[5\] _01899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_120_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07549__I _02396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_315_clock_I clknet_5_17_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09965__S _04734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08136_ _03569_ _00028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11612__I1 u2.mem\[175\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_4_3_0_clock_I clknet_3_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08067_ _01954_ _03516_ _03519_ _00009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_162_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09569__I0 _04489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07018_ _02405_ _02391_ _02392_ _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA__13193__CLK clknet_leaf_292_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08241__I0 _03548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07744__A2 _03027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08969_ _04026_ u2.mem\[20\]\[5\] _04102_ _04104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_124_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11735__S _05840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11980_ _05222_ u2.mem\[194\]\[12\] _05985_ _05988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_17_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10931_ _05332_ _01060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11534__I _05673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06704__C2 u2.mem\[192\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10862_ _05200_ u2.mem\[129\]\[2\] _05287_ _05290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09004__I _04126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12601_ _00480_ clknet_leaf_135_clock u2.mem\[29\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10793_ _05248_ _01006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12532_ _00411_ clknet_leaf_101_clock u2.mem\[25\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08843__I _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12463_ _00342_ clknet_leaf_174_clock u2.mem\[21\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06483__A2 _01960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11414_ _05639_ _01236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12410__CLK clknet_leaf_124_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12394_ _00273_ clknet_leaf_140_clock u2.mem\[16\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11345_ _05595_ u2.mem\[158\]\[5\] _05584_ _05596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07983__A2 _02594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_284_clock clknet_5_20_0_clock clknet_leaf_284_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_49_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11276_ _05552_ u2.mem\[154\]\[3\] _05546_ _05553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11367__I0 _05587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13015_ _00894_ clknet_leaf_149_clock u2.mem\[55\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12560__CLK clknet_leaf_159_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10227_ _04582_ _04898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07194__I _02549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07735__A2 _03160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09980__I0 _04694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10158_ _04808_ u2.mem\[47\]\[11\] _04851_ _04855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold3 output_active_hold\[1\] net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_48_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_299_clock clknet_5_21_0_clock clknet_leaf_299_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_82_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10089_ _04611_ _04815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_264_clock_I clknet_5_22_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_222_clock clknet_5_29_0_clock clknet_leaf_222_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_1_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06538__I _02022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13066__CLK clknet_leaf_339_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08999__A1 _04121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06320_ u2.mem\[187\]\[3\] _01633_ _01636_ u2.mem\[192\]\[3\] _01824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_237_clock clknet_5_25_0_clock clknet_leaf_237_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06251_ _01592_ _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06474__A2 _01960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09785__S _04628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06273__I _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06182_ _01688_ _01689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07423__A1 _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12903__CLK clknet_leaf_147_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09941_ _04691_ u2.mem\[42\]\[4\] _04724_ _04725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09872_ _04678_ _00655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09971__I0 _04685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08823_ _03987_ _04011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11555__S _05721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08754_ _03916_ u2.mem\[15\]\[5\] _03967_ _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07705_ _03170_ _03171_ _03172_ _03173_ _03174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08685_ _03700_ _03927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13409__CLK clknet_leaf_319_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07636_ u2.mem\[27\]\[9\] _03104_ _03105_ u2.mem\[35\]\[9\] _03106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07567_ _03029_ _03032_ _03035_ _03037_ _03038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_53_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11290__S _05559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09306_ _04272_ u2.mem\[27\]\[9\] _04323_ _04325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10097__I0 _04782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06518_ _02002_ _02003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12433__CLK clknet_leaf_171_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07498_ u2.mem\[6\]\[6\] _02927_ _02928_ u2.mem\[47\]\[6\] _02971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11833__I1 u2.mem\[189\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07257__A4 _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13559__CLK clknet_leaf_33_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09237_ _04173_ _04283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06449_ _01878_ _01938_ _01941_ _01944_ _01469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06465__A2 _01955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09168_ _04225_ _04236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_119_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08119_ _03557_ u2.mem\[1\]\[5\] _03555_ _03558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07414__A1 _02882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12583__CLK clknet_leaf_112_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09099_ _04164_ u2.mem\[22\]\[11\] _04192_ _04196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11130_ _05432_ u2.mem\[145\]\[5\] _05452_ _05459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06911__I _02376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11349__I0 _05583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11061_ _05416_ _01106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10012_ _04765_ _00708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_7_0_clock_I clknet_4_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07717__A2 _03132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08765__I1 u2.mem\[15\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11963_ _05978_ _01446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13089__CLK clknet_leaf_257_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11264__I _05499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11521__I0 _05680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10914_ _05303_ u2.mem\[132\]\[3\] _05319_ _05323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_75_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08774__S _03977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11894_ u2.mem\[192\]\[7\] _03514_ _05937_ _05939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07350__B1 _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10845_ _05198_ u2.mem\[128\]\[1\] _05278_ _05280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09669__I _04543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13564_ _01443_ clknet_leaf_10_clock u2.mem\[194\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10776_ _05207_ u2.mem\[62\]\[5\] _05237_ _05239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12515_ _00394_ clknet_leaf_109_clock u2.mem\[24\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06456__A2 _01938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13495_ _01374_ clknet_leaf_328_clock u2.mem\[186\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10608__I _05130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12926__CLK clknet_leaf_221_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07189__I _02554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12446_ _00325_ clknet_leaf_188_clock u2.mem\[20\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07405__A1 _02875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12377_ _00256_ clknet_leaf_114_clock u2.mem\[15\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10260__I0 _04920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07956__A2 _03417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11328_ _04393_ _05566_ _05584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_125_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11259_ _05541_ _01179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07708__A2 _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12306__CLK clknet_leaf_173_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06977__B _02454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11760__I0 _05837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11375__S _05607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07652__I _02513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_161_clock clknet_5_27_0_clock clknet_leaf_161_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08470_ _03705_ u2.mem\[8\]\[11\] _03787_ _03791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06268__I _01772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06144__A1 _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12456__CLK clknet_leaf_128_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07341__B1 _02660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07421_ u2.mem\[49\]\[5\] _02817_ _02818_ u2.mem\[46\]\[5\] _02895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_39_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10719__S _05196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_176_clock clknet_5_27_0_clock clknet_leaf_176_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08483__I _03798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07352_ _02543_ _02827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11815__I1 u2.mem\[188\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06303_ _01773_ _01555_ _01807_ _01482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_31_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07283_ u2.mem\[49\]\[3\] _02528_ _02532_ u2.mem\[46\]\[3\] _02759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11440__A2 _05645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10518__I _05072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09022_ _04140_ u2.mem\[21\]\[4\] _04141_ _04142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06234_ u2.mem\[170\]\[1\] _01687_ _01689_ u2.mem\[156\]\[1\] _01740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_163_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06165_ _01665_ _01591_ _01623_ _01672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_85_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10251__I0 _04913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06096_ _01566_ _01600_ _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_46_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09149__A1 _04224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_114_clock clknet_5_14_0_clock clknet_leaf_114_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09924_ _04611_ _04714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10253__I _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09855_ _04586_ u2.mem\[40\]\[6\] _04666_ _04669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08806_ _04001_ _00266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13231__CLK clknet_leaf_302_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06998_ _02407_ _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_09786_ _04629_ _00618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06383__A1 u2.mem\[171\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07562__I _02464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_129_clock clknet_5_15_0_clock clknet_leaf_129_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06922__A3 _02382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08737_ _03936_ u2.mem\[14\]\[14\] _03956_ _03959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11503__I0 _05674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09321__A1 _03629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08668_ _03915_ _00214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06135__A1 _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07332__B1 _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13381__CLK clknet_leaf_319_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_7_clock_I clknet_5_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07619_ _02616_ _03090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06686__A2 _02156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08599_ _03855_ _03871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10629__S _05146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11812__I _05887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12949__CLK clknet_leaf_63_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10630_ _05148_ _00943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06906__I _02384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07511__B _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11806__I1 u2.mem\[187\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06438__A2 _01931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10561_ _05103_ u2.mem\[57\]\[4\] _05104_ _05105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_167_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08683__I0 _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12300_ _00179_ clknet_leaf_200_clock u2.mem\[11\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10490__I0 _05011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13280_ _01159_ clknet_leaf_380_clock u2.mem\[150\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10492_ _05014_ u2.mem\[55\]\[9\] _05061_ _05063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12231_ _00110_ clknet_leaf_54_clock u2.mem\[6\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08435__I0 _03714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07399__B1 _02872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12162_ _00041_ clknet_leaf_236_clock u2.mem\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12329__CLK clknet_leaf_135_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06071__B1 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11113_ _05449_ _01125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06071__C2 u2.mem\[193\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12093_ _00017_ clknet_leaf_380_clock u3.enable vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06610__A2 _02092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11044_ _05406_ _01099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06374__A1 _01844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12479__CLK clknet_leaf_176_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12995_ _00874_ clknet_leaf_31_clock u2.mem\[54\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06088__I _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06126__A1 _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11946_ _05227_ u2.mem\[193\]\[14\] _05965_ _05968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_93_clock clknet_5_10_0_clock clknet_leaf_93_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11877_ _05928_ _05929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06141__A4 _01647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10828_ _05252_ _05268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_38_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10338__I _04965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13547_ _01426_ clknet_leaf_36_clock u2.mem\[193\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10759_ _05228_ _00992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10481__I0 _05001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13478_ _01357_ clknet_leaf_307_clock u2.mem\[183\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12429_ _00308_ clknet_leaf_192_clock u2.mem\[19\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_161_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08426__I0 _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07929__A2 _03383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07647__I _02500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_31_clock clknet_5_3_0_clock clknet_leaf_31_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_154_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08051__A1 _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07970_ u2.mem\[43\]\[15\] _03286_ _03287_ u2.mem\[20\]\[15\] _03434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06601__A2 _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13254__CLK clknet_leaf_308_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06921_ _02399_ _02400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_45_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09640_ _04521_ _04532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06852_ u2.mem\[179\]\[5\] _02150_ _02152_ u2.mem\[191\]\[5\] _02332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10801__I _05252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06365__A1 u2.mem\[144\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07382__I _02616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06904__A3 _02382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09571_ _04166_ _04491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06783_ _02261_ _02262_ _02263_ _02264_ _02265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_08522_ _03798_ _03826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__11833__S _05896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06117__A1 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08453_ _03781_ _00133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07865__A1 _01969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_161_clock_I clknet_5_27_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07404_ u2.mem\[3\]\[5\] _02803_ _02749_ _02878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08384_ _03697_ u2.mem\[6\]\[9\] _03737_ _03739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11996__CLK clknet_leaf_334_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07617__A1 _03078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07335_ u2.mem\[53\]\[4\] _02808_ _02809_ u2.mem\[56\]\[4\] _02810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_104_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10472__I0 _04987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07266_ u2.mem\[32\]\[3\] _02385_ _02397_ u2.mem\[2\]\[3\] _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_104_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09005_ _04127_ _04128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06217_ _01674_ _01697_ _01718_ _01723_ _01724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_118_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08417__I0 _03680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07197_ _02566_ _02675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06840__A2 _02075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07557__I _02451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09973__S _04740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06148_ u2.mem\[189\]\[0\] _01650_ _01652_ u2.mem\[176\]\[0\] u2.mem\[172\]\[0\]
+ _01654_ _01655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__08042__A1 _01773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09090__I0 _04151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11079__I _05345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_21_0_clock clknet_4_10_0_clock clknet_5_21_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_06079_ _01584_ _01559_ _01585_ _01586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10912__S _05319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12621__CLK clknet_leaf_201_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_86_clock_I clknet_5_9_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09907_ _04702_ _00666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09838_ _04658_ _00641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06356__A1 u2.mem\[159\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06356__B2 u2.mem\[149\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09769_ _04570_ u2.mem\[38\]\[1\] _04618_ _04620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12771__CLK clknet_leaf_83_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11800_ _05868_ u2.mem\[187\]\[1\] _05879_ _05881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06108__A1 _01612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12780_ _00659_ clknet_leaf_268_clock u2.mem\[41\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07305__B1 _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11731_ _05837_ u2.mem\[182\]\[5\] _05826_ _05838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10359__S _04976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06636__I _02120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12001__CLK clknet_leaf_41_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11662_ _05794_ u2.mem\[178\]\[3\] _05788_ _05795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13127__CLK clknet_leaf_39_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13401_ _01280_ clknet_leaf_318_clock u2.mem\[170\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10613_ _05108_ u2.mem\[58\]\[6\] _05136_ _05139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11593_ _05751_ _01303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_5_15_0_clock_I clknet_4_7_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10544_ _05092_ _00913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13332_ _01211_ clknet_leaf_6_clock u2.mem\[158\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07084__A2 _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12151__CLK clknet_leaf_56_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08408__I0 _03663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_363_clock_I clknet_5_4_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06831__A2 _02029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13263_ _01142_ clknet_leaf_286_clock u2.mem\[147\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13277__CLK clknet_leaf_8_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10475_ _05053_ _00883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10215__I0 _04889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09883__S _04683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12214_ _00093_ clknet_leaf_72_clock u2.mem\[5\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08033__A1 _03491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09081__I0 _04136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13194_ _01073_ clknet_leaf_287_clock u2.mem\[135\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12145_ _00024_ clknet_leaf_230_clock u2.mem\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10822__S _05263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12076_ data_in_trans\[13\].A clknet_leaf_39_clock data_in_trans\[13\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07139__A3 _02615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11027_ _05396_ _01092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08298__I _03673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06347__B2 u2.mem\[183\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11191__I1 u2.mem\[149\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11653__S _05788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12978_ _00857_ clknet_leaf_265_clock u2.mem\[53\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09123__S _04208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08895__I0 _04030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11929_ _05958_ _01432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08962__S _04097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06546__I _02005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06990__B _02424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07120_ _02598_ _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07051_ _02480_ _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_173_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06822__A2 _02300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07377__I _02603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06002_ u2.select_mem_row\[0\] _01502_ _01510_ _01511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12644__CLK clknet_leaf_94_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08024__A1 _03480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10906__A1 _04095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_108_clock_I clknet_5_11_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10732__S _05205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06586__A1 _02060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07953_ u2.mem\[32\]\[15\] _03252_ _03253_ u2.mem\[2\]\[15\] _03417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_87_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06904_ _02377_ _02381_ _02382_ _02383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA__12794__CLK clknet_leaf_338_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07884_ u2.mem\[43\]\[13\] _03286_ _03287_ u2.mem\[20\]\[13\] _03350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06338__A1 _01814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09623_ _04463_ u2.mem\[35\]\[0\] _04522_ _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07045__C _02450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06835_ u2.mem\[187\]\[5\] _02100_ _02101_ u2.mem\[192\]\[5\] _02315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_55_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08936__I _04073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09554_ _04479_ _00536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06766_ _02246_ _02247_ _02248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12024__CLK clknet_leaf_321_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07840__I _02579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08505_ _03687_ _03814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08886__I0 _04021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09485_ _04387_ u2.mem\[31\]\[13\] _04434_ _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06697_ u2.mem\[167\]\[1\] _02058_ _02061_ u2.mem\[183\]\[1\] _02181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11362__I _05605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10693__I0 _05112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08436_ _03770_ _00127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12174__CLK clknet_leaf_232_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08367_ _03729_ _00099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07318_ _02785_ _02788_ _02791_ _02792_ _02793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07066__A2 _02542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08298_ _03673_ _03674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07249_ u2.mem\[29\]\[2\] _02559_ _02564_ u2.mem\[11\]\[2\] _02726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10260_ _04920_ u2.mem\[49\]\[15\] _04914_ _04921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10748__I1 u2.mem\[61\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07369__A3 _02840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10191_ _04864_ _04875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08112__S _03546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12901_ _00780_ clknet_leaf_70_clock u2.mem\[48\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12832_ _00711_ clknet_leaf_164_clock u2.mem\[44\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08846__I _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12763_ _00642_ clknet_leaf_219_clock u2.mem\[40\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12517__CLK clknet_leaf_107_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11272__I _05507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11714_ _04179_ _05808_ _05826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10684__I0 _05103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12694_ _00573_ clknet_leaf_82_clock u2.mem\[35\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11645_ _05783_ _01323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_161_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08581__I _03855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12667__CLK clknet_leaf_211_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput15 data_in_a[2] net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_167_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11576_ _05711_ u2.mem\[173\]\[1\] _05739_ _05741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinput26 mem_address_a[2] net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_156_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput37 row_select_a[0] net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13315_ _01194_ clknet_leaf_316_clock u2.mem\[156\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10527_ _05072_ _05083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06804__A2 _02282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07197__I _02566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10458_ _05043_ _00876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13246_ _01125_ clknet_leaf_289_clock u2.mem\[144\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10739__I1 u2.mem\[61\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11648__S _05778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06568__A1 _02052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13177_ _01056_ clknet_leaf_292_clock u2.mem\[133\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10389_ _04997_ _04998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09118__S _04203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12128_ _01469_ clknet_leaf_37_clock u2.driver_mem\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07780__A3 _03246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12059_ net18 clknet_2_1__leaf_clock_a data_in_trans\[5\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12047__CLK clknet_2_2__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11313__A1 _05411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11164__I1 u2.mem\[147\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06985__B _02383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06620_ _02056_ _02104_ _02105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06740__A1 _02219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06551_ _02008_ _01989_ _02036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_59_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12197__CLK clknet_leaf_23_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13442__CLK clknet_leaf_364_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09270_ _04303_ _00428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06099__A3 _01599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_34_clock_I clknet_5_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06482_ u2.mem\[192\]\[12\] _01929_ _01971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08221_ _03570_ u2.mem\[3\]\[11\] _03618_ _03622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08152_ _03580_ _00033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07048__A2 _02433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07103_ _02581_ _02582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08083_ _03530_ _03528_ _03531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_3_3_0_clock_I clknet_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07034_ _02455_ _02510_ _02511_ _02512_ _02513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_173_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_259_clock_I clknet_5_19_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10462__S _05045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07835__I _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07756__B1 _03126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07220__A2 _02681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08985_ _04041_ u2.mem\[20\]\[12\] _04112_ _04113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07936_ u2.mem\[29\]\[14\] _03301_ _03302_ u2.mem\[11\]\[14\] _03401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_102_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input26_I mem_address_a[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07867_ u2.mem\[32\]\[13\] _03252_ _03253_ u2.mem\[2\]\[13\] _03333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_leaf_311_clock_I clknet_5_17_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09606_ _04485_ u2.mem\[34\]\[9\] _04511_ _04513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07523__A3 _02989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08666__I _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06818_ _02296_ _02297_ _02298_ _02299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07798_ u2.mem\[1\]\[12\] _03263_ _03264_ u2.mem\[7\]\[12\] _03265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07570__I _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09537_ _04467_ u2.mem\[33\]\[1\] _04465_ _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06749_ u2.mem\[185\]\[2\] _02121_ _02123_ u2.mem\[173\]\[2\] _02232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_19_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10666__I0 _05124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09520__I1 u2.mem\[32\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09468_ _04426_ _00503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07287__A2 _02666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08419_ _03684_ u2.mem\[7\]\[6\] _03758_ _03761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10637__S _05152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09399_ _04383_ _00477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11430_ _05627_ u2.mem\[164\]\[1\] _05647_ _05649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10043__A1 _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11361_ _04439_ _05274_ _05605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_165_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10312_ _04898_ u2.mem\[51\]\[5\] _04949_ _04951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06798__B2 u2.mem\[183\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13100_ _00979_ clknet_leaf_281_clock u2.mem\[61\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11292_ _05552_ u2.mem\[155\]\[3\] _05559_ _05563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10243_ _04598_ _04909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13031_ _00910_ clknet_leaf_51_clock u2.mem\[56\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11543__A1 _04310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11394__I1 u2.mem\[162\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10174_ _04782_ u2.mem\[48\]\[0\] _04865_ _04866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13315__CLK clknet_leaf_316_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10171__I _04862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13465__CLK clknet_leaf_362_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06722__A1 u2.mem\[164\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12815_ _00694_ clknet_leaf_167_clock u2.mem\[43\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10657__I0 _05115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09511__I1 u2.mem\[32\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07278__A2 _02476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12746_ _00625_ clknet_leaf_44_clock u2.mem\[38\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12677_ _00556_ clknet_leaf_84_clock u2.mem\[34\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11730__I _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10409__I0 _05011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11628_ _05752_ u2.mem\[176\]\[2\] _05771_ _05774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11559_ _05730_ _05731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06789__A1 _02255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09027__I0 _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07450__A2 _02922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_260_clock_I clknet_5_22_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10282__S _04933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13229_ _01108_ clknet_leaf_301_clock u2.mem\[141\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07655__I _02520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07738__B1 _03185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11385__I1 u2.mem\[161\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07202__A2 _02580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08770_ _03931_ u2.mem\[15\]\[12\] _03977_ _03978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07721_ _03186_ _03187_ _03188_ _03189_ _03190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_113_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_4_10_0_clock_I clknet_3_5_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08486__I _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07652_ _02513_ _03122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06713__A1 u2.mem\[153\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06713__B2 u2.mem\[152\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06603_ _01992_ _02080_ _02088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07583_ _02507_ _03054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09502__I1 u2.mem\[32\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06534_ _02015_ _02018_ _02019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09322_ _04333_ _04334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10648__I0 _05106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_167_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09253_ _04258_ u2.mem\[26\]\[3\] _04290_ _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_146_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06465_ _01954_ _01955_ _01956_ _01957_ _01472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10457__S _05040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12982__CLK clknet_leaf_55_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08204_ _03612_ _00053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09184_ _04177_ u2.mem\[24\]\[15\] _04241_ _04245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06396_ u2.mem\[153\]\[5\] _01707_ _01709_ u2.mem\[160\]\[5\] _01898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_147_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08135_ _03568_ u2.mem\[1\]\[10\] _03564_ _03569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06229__B1 _01734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10256__I _04611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12212__CLK clknet_leaf_72_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08066_ _03517_ _03518_ _03519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13338__CLK clknet_leaf_6_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07017_ u2.mem\[50\]\[0\] _02493_ _02495_ u2.mem\[51\]\[0\] _02496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11288__S _05559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07992__A3 _03454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07729__B1 _03083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07565__I _02469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_7_0_clock_I clknet_3_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12362__CLK clknet_leaf_137_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13488__CLK clknet_leaf_314_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06401__B1 _01721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08968_ _04103_ _00326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08597__S _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06952__A1 _02363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11128__I1 u2.mem\[145\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07919_ u2.mem\[50\]\[14\] _02493_ _02495_ u2.mem\[51\]\[14\] _03384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08899_ _04062_ _00298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10930_ _05305_ u2.mem\[133\]\[4\] _05326_ _05332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06704__A1 u2.mem\[188\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06704__B2 u2.mem\[187\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10861_ _05289_ _01033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12600_ _00479_ clknet_leaf_115_clock u2.mem\[29\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10639__I0 _05097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10792_ _05222_ u2.mem\[62\]\[12\] _05247_ _05248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12531_ _00410_ clknet_leaf_111_clock u2.mem\[25\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12462_ _00341_ clknet_leaf_193_clock u2.mem\[21\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06644__I _02128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07680__A2 _03148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09020__I _04139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11413_ _05623_ u2.mem\[163\]\[0\] _05638_ _05639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11064__I0 _05390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12393_ _00272_ clknet_leaf_140_clock u2.mem\[16\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07968__B1 _02525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11344_ _05516_ _05595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07432__A2 _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12705__CLK clknet_leaf_242_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11275_ _05510_ _05552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11367__I1 u2.mem\[160\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13014_ _00893_ clknet_leaf_66_clock u2.mem\[55\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10226_ _04897_ _00790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11926__S _05955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10157_ _04854_ _00764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold4 output_active_hold\[2\] net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XANTENNA__12855__CLK clknet_leaf_143_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10088_ _04814_ _00735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_207_clock_I clknet_5_30_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_169_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09496__I0 _04356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06459__B1 _01948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10277__S _04928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12729_ _00608_ clknet_leaf_45_clock u2.mem\[37\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11460__I _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06250_ u2.mem\[159\]\[1\] _01604_ _01595_ u2.mem\[149\]\[1\] _01756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12235__CLK clknet_leaf_230_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06554__I _02038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10076__I _04598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06181_ _01557_ _01630_ _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12385__CLK clknet_leaf_235_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09940_ _04718_ _04724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_171_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07385__I _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09871_ _04609_ u2.mem\[40\]\[13\] _04676_ _04678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07187__A1 _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08822_ _03655_ _04010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09306__S _04323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08753_ _03968_ _00246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07704_ u2.mem\[3\]\[10\] _03036_ _02982_ _03173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08684_ _03926_ _00219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07635_ _02425_ _03105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06162__A2 _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09487__I0 _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07566_ u2.mem\[3\]\[8\] _03036_ _02982_ _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_41_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09305_ _04324_ _00442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11294__I0 _05554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06517_ _01999_ _02001_ _02002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_344_clock clknet_5_7_0_clock clknet_leaf_344_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07497_ u2.mem\[8\]\[6\] _02860_ _02861_ u2.mem\[4\]\[6\] _02970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09236_ _04282_ _00415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08880__S _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06448_ u2.mem\[193\]\[5\] _01942_ _01943_ u2.mem\[194\]\[5\] _01934_ _01944_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__13160__CLK clknet_leaf_293_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12118__D _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09167_ _04235_ _00393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06379_ u2.mem\[180\]\[5\] _01664_ _01667_ u2.mem\[150\]\[5\] _01881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_108_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12728__CLK clknet_leaf_44_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09775__I _04617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_359_clock clknet_5_5_0_clock clknet_leaf_359_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08118_ _03510_ _03557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07414__A2 _02885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06217__A3 _01718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09098_ _04195_ _00364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08049_ _03505_ _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_3_clock_I clknet_5_0_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11349__I1 u2.mem\[159\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_156_clock_I clknet_5_24_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11060_ _05386_ u2.mem\[141\]\[2\] _05413_ _05416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12878__CLK clknet_leaf_225_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09411__I0 _04391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10011_ _04687_ u2.mem\[44\]\[2\] _04762_ _04765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06925__A1 _02352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06386__C1 u2.mem\[163\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11962_ _05913_ u2.mem\[194\]\[4\] _05975_ _05978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09015__I _04135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10913_ _05322_ _01052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06153__A2 _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11893_ _05938_ _01416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07350__A1 u2.mem\[61\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09478__I0 _04380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12258__CLK clknet_leaf_241_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10844_ _05279_ _01026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_16_0_clock clknet_4_8_0_clock clknet_5_16_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_129_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10097__S _04820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13563_ _01442_ clknet_leaf_10_clock u2.mem\[194\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10775_ _05238_ _00998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_160_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12514_ _00393_ clknet_leaf_174_clock u2.mem\[24\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09886__S _04683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13494_ _01373_ clknet_leaf_309_clock u2.mem\[185\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12445_ _00324_ clknet_leaf_187_clock u2.mem\[20\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07405__A2 _02876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12376_ _00255_ clknet_leaf_61_clock u2.mem\[15\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09650__I0 _04491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11327_ _05499_ _05583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09402__I0 _04384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11258_ _05511_ u2.mem\[153\]\[3\] _05537_ _05541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11656__S _05788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10209_ _04564_ _04885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06377__C1 u2.mem\[172\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11189_ _05468_ u2.mem\[149\]\[3\] _05492_ _05496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_171_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06977__C _02455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11760__I1 u2.mem\[184\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13033__CLK clknet_leaf_51_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_358_clock_I clknet_5_5_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06144__A2 _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07341__B2 u2.mem\[12\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07420_ u2.mem\[14\]\[5\] _02892_ _02893_ u2.mem\[12\]\[5\] _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_78_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07892__A2 _02567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09469__I0 _04371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06695__A3 _02175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13183__CLK clknet_leaf_294_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11276__I0 _05552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07351_ _02541_ _02826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09796__S _04633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06302_ _01780_ _01784_ _01793_ _01806_ _01807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_52_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07282_ u2.mem\[14\]\[3\] _02659_ _02660_ u2.mem\[12\]\[3\] _02758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09021_ _04123_ _04141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_136_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11028__I0 _05384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06233_ u2.mem\[173\]\[1\] _01720_ _01722_ u2.mem\[185\]\[1\] _01739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06852__B1 _02152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10735__S _05205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06164_ _01670_ _01671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09641__I0 _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07329__B _02749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06095_ _01601_ _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09923_ _04713_ _00671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_160_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11566__S _05731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09854_ _04668_ _00647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06907__A1 _02364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08805_ _03922_ u2.mem\[16\]\[8\] _04000_ _04001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09785_ _04592_ u2.mem\[38\]\[8\] _04628_ _04629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06997_ _02475_ _02476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06383__A2 _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08736_ _03958_ _00239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12400__CLK clknet_leaf_172_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11503__I1 u2.mem\[168\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13526__CLK clknet_leaf_327_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08667_ _03913_ u2.mem\[13\]\[4\] _03914_ _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06135__A2 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07618_ u2.mem\[5\]\[8\] _02922_ _02923_ u2.mem\[38\]\[8\] _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_26_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08598_ _03870_ _00189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_283_clock clknet_5_22_0_clock clknet_leaf_283_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_126_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11267__I0 _05544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07549_ _02396_ _03020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_82_clock_I clknet_5_8_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12550__CLK clknet_leaf_100_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08132__I0 _03566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06194__I _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10560_ _05094_ _05104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09880__I0 _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11019__I0 _05390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09219_ _04269_ u2.mem\[25\]\[8\] _04270_ _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_298_clock clknet_5_21_0_clock clknet_leaf_298_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_154_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10491_ _05062_ _00890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12230_ _00109_ clknet_leaf_73_clock u2.mem\[6\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_163_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09632__I0 _04473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07399__A1 u2.mem\[27\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12161_ _00040_ clknet_leaf_237_clock u2.mem\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_221_clock clknet_5_29_0_clock clknet_leaf_221_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06071__A1 u2.mem\[158\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11112_ _05428_ u2.mem\[144\]\[3\] _05445_ _05449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06071__B2 u2.mem\[151\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12092_ inverter_select_trans.A clknet_leaf_304_clock inverter_select_trans.data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08199__I0 _03548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13056__CLK clknet_leaf_256_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11043_ _05384_ u2.mem\[140\]\[1\] _05404_ _05406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_46_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08849__I _03687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_236_clock clknet_5_25_0_clock clknet_leaf_236_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_65_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11275__I _05510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12080__CLK clknet_leaf_348_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12994_ _00873_ clknet_leaf_251_clock u2.mem\[54\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11945_ _05967_ _01439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06126__A2 _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06677__A3 _02140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11876_ _05927_ _05928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10827_ _05267_ _01021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13546_ _01425_ clknet_leaf_38_clock u2.mem\[192\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10758_ _05227_ u2.mem\[61\]\[14\] _05223_ _05228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09871__I0 _04609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13477_ _01356_ clknet_leaf_305_clock u2.mem\[183\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10689_ _05182_ _00968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12428_ _00307_ clknet_leaf_192_clock u2.mem\[19\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09623__I0 _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07929__A3 _03388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11430__I0 _05627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12359_ _00238_ clknet_leaf_138_clock u2.mem\[14\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06598__C1 u2.mem\[145\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06920_ _02355_ _02379_ _02399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07663__I _02554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06851_ u2.mem\[170\]\[5\] _02145_ _02147_ u2.mem\[156\]\[5\] _02331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06365__A2 _01670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09570_ _04490_ _00541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06782_ u2.mem\[176\]\[3\] _02002_ _02019_ u2.mem\[189\]\[3\] _02264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_82_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08521_ _03708_ _03825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11497__I0 _05663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06117__A2 _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12573__CLK clknet_leaf_201_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_104_clock_I clknet_5_10_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08452_ _03671_ u2.mem\[8\]\[3\] _03777_ _03781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07403_ u2.mem\[16\]\[5\] _02800_ _02801_ u2.mem\[33\]\[5\] _02877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08383_ _03738_ _00106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07334_ _02482_ _02809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09862__I0 _04596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06825__B1 _02068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07265_ u2.mem\[45\]\[3\] _02633_ _02634_ u2.mem\[34\]\[3\] _02741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07838__I _02576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09004_ _04126_ _04127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06216_ u2.mem\[173\]\[0\] _01720_ _01722_ u2.mem\[185\]\[0\] _01723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06742__I _02126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08417__I1 u2.mem\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07196_ _02668_ _02669_ _02670_ _02673_ _02674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_118_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13079__CLK clknet_leaf_47_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11421__I0 _05633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06147_ _01653_ _01654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07250__B1 _02577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06078_ _01573_ _01574_ _01585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_29_clock_I clknet_5_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11296__S _05558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09906_ _04700_ u2.mem\[41\]\[8\] _04701_ _04702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08669__I _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07573__I _02486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09837_ _04615_ u2.mem\[39\]\[15\] _04654_ _04658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06356__A2 _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07553__B2 u2.mem\[30\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12916__CLK clknet_leaf_87_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09768_ _04619_ _00610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08719_ _03918_ u2.mem\[14\]\[6\] _03946_ _03949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11488__I0 _05674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06108__A2 _01613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09699_ _04566_ _04567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_162_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08353__I0 _03718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11730_ _03678_ _05837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11661_ _05673_ _05794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13400_ _01279_ clknet_leaf_313_clock u2.mem\[170\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10612_ _05138_ _00935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09853__I0 _04583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11592_ _05750_ u2.mem\[174\]\[1\] _05748_ _05751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13331_ _01210_ clknet_leaf_2_clock u2.mem\[158\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06816__B1 _02200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10543_ _05027_ u2.mem\[56\]\[15\] _05088_ _05092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_306_clock_I clknet_5_20_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13262_ _01141_ clknet_leaf_310_clock u2.mem\[147\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10474_ _04992_ u2.mem\[55\]\[1\] _05051_ _05053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_170_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_160_clock clknet_5_27_0_clock clknet_leaf_160_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10215__I1 u2.mem\[49\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12213_ _00092_ clknet_leaf_23_clock u2.mem\[5\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_5_19_0_clock_I clknet_4_9_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13193_ _01072_ clknet_leaf_292_clock u2.mem\[135\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12446__CLK clknet_leaf_188_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12144_ _00023_ clknet_leaf_230_clock u2.mem\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12075_ net11 clknet_2_0__leaf_clock_a data_in_trans\[13\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_175_clock clknet_5_27_0_clock clknet_leaf_175_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_42_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07139__A4 _02383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11026_ _05380_ u2.mem\[139\]\[0\] _05395_ _05396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07544__A1 _03000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12596__CLK clknet_leaf_95_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12977_ _00856_ clknet_leaf_253_clock u2.mem\[53\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11928_ _05209_ u2.mem\[193\]\[6\] _05955_ _05958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11859_ _04416_ _05886_ _05917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_113_clock clknet_5_11_0_clock clknet_leaf_113_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_92_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09844__I0 _04570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06990__C _02459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13529_ _01408_ clknet_leaf_332_clock u2.mem\[191\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13221__CLK clknet_leaf_300_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07050_ _02478_ _02529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07480__B1 _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_128_clock clknet_5_15_0_clock clknet_leaf_128_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_103_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06822__A3 _02301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06001_ _01505_ _01502_ _01510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11403__I0 _05631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07232__B1 _02648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13371__CLK clknet_leaf_375_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_30_clock_I clknet_5_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06586__A2 _02070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08489__I _03666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07952_ u2.mem\[45\]\[15\] _02432_ _02436_ u2.mem\[34\]\[15\] _03416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12939__CLK clknet_leaf_225_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07393__I _02435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06903_ _02351_ _02382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_96_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07883_ u2.mem\[49\]\[13\] _03283_ _03284_ u2.mem\[46\]\[13\] _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07535__A1 u2.mem\[17\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06338__A2 _01819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09622_ _04521_ _04522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_68_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06834_ _02310_ _02311_ _02312_ _02313_ _02314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_28_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09553_ _04478_ u2.mem\[33\]\[6\] _04474_ _04479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06765_ u2.mem\[153\]\[3\] _02196_ _02200_ u2.mem\[160\]\[3\] _02247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_71_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08504_ _03813_ _00152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07299__B1 _02601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09484_ _04435_ _00510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06696_ u2.mem\[164\]\[1\] _02050_ _02053_ u2.mem\[178\]\[1\] _02180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_36_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10259__I _04614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08435_ _03714_ u2.mem\[7\]\[13\] _03768_ _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12319__CLK clknet_leaf_161_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08366_ _03663_ u2.mem\[6\]\[1\] _03727_ _03729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09835__I0 _04612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07317_ u2.mem\[27\]\[4\] _02638_ _02639_ u2.mem\[35\]\[4\] _02792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11642__I0 _05752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08297_ _03505_ _03673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09984__S _04745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06274__A1 u2.mem\[184\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12469__CLK clknet_leaf_104_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07248_ u2.mem\[26\]\[2\] _02675_ _02676_ u2.mem\[10\]\[2\] _02725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_125_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07471__B1 _02809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07179_ _02517_ _02657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07223__B1 _02397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_92_clock clknet_5_10_0_clock clknet_leaf_92_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10190_ _04874_ _00777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12900_ _00779_ clknet_leaf_70_clock u2.mem\[48\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11754__S _05849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12831_ _00710_ clknet_leaf_163_clock u2.mem\[44\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12762_ _00641_ clknet_leaf_51_clock u2.mem\[39\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_30_clock clknet_5_3_0_clock clknet_leaf_30_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_14_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11713_ _03654_ _05825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12693_ _00572_ clknet_leaf_82_clock u2.mem\[35\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13244__CLK clknet_leaf_295_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09958__I _04718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08862__I _03704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11644_ _05754_ u2.mem\[177\]\[3\] _05779_ _05783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09826__I0 _04599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_45_clock clknet_5_6_0_clock clknet_leaf_45_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11575_ _05740_ _01296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput16 data_in_a[3] net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput27 mem_address_a[3] net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_35_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_5_30_0_clock_I clknet_4_15_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput38 row_select_a[1] net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_13314_ _01193_ clknet_5_5_0_clock u2.mem\[155\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06265__A1 _01745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07462__B1 _02872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10526_ _05082_ _00905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06804__A3 _02283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13245_ _01124_ clknet_leaf_307_clock u2.mem\[144\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10457_ _05016_ u2.mem\[54\]\[10\] _05040_ _05043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08006__A2 _03458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10833__S _05268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13176_ _01055_ clknet_leaf_284_clock u2.mem\[132\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10388_ _04134_ _04997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06568__A2 _01999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12127_ _01468_ clknet_leaf_36_clock u2.driver_mem\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08102__I _03545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12058_ data_in_trans\[4\].A clknet_leaf_375_clock data_in_trans\[4\].data_sync vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07517__A1 _02985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08565__I0 _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11009_ _05339_ _05384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10372__I0 _04920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09134__S _04213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06985__C _02463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06550_ _02034_ _02035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10124__I0 _04810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10079__I _04601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06481_ _01920_ _01970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06099__A4 _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08220_ _03621_ _00060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09868__I _04660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09817__I0 _04586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08151_ _03579_ u2.mem\[1\]\[15\] _03573_ _03580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11624__I0 _05746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07102_ _02573_ _02574_ _02442_ _02575_ _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_174_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08082_ data_in_trans\[13\].data_sync _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07033_ _02441_ _02429_ _02382_ _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_146_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12761__CLK clknet_leaf_51_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_7_0_clock_I clknet_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08984_ _04096_ _04112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_142_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07220__A3 _02688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13117__CLK clknet_leaf_276_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07935_ u2.mem\[26\]\[14\] _02567_ _02569_ u2.mem\[10\]\[14\] _03400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_87_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08556__I0 _03819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11574__S _05739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07866_ u2.mem\[45\]\[13\] _02432_ _02436_ u2.mem\[34\]\[13\] _03332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_29_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10363__I0 _04911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07851__I _02603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09044__S _04155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09605_ _04512_ _00554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input19_I data_in_a[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06817_ u2.mem\[148\]\[4\] _02129_ _02131_ u2.mem\[152\]\[4\] _02298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07523__A4 _02994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07797_ _02460_ _03264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12141__CLK clknet_leaf_231_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06731__A2 _02211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13267__CLK clknet_leaf_384_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09536_ _04127_ _04467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10115__I0 _04801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06748_ u2.mem\[154\]\[2\] _02225_ _02226_ u2.mem\[162\]\[2\] _02230_ _02231_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09467_ _04369_ u2.mem\[31\]\[5\] _04424_ _04426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11863__I0 _05907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10918__S _05318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06679_ _01545_ _01996_ _02163_ _01474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_24_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08418_ _03760_ _00119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12291__CLK clknet_leaf_110_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08682__I _03696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07692__B1 _03161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09398_ _04382_ u2.mem\[29\]\[11\] _04376_ _04383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09808__I0 _04573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08349_ _03715_ _00095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10043__A2 _04760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11360_ _05604_ _01217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06798__A2 _02058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10311_ _04950_ _00822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11291_ _05562_ _01190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09219__S _04270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13030_ _00909_ clknet_leaf_66_clock u2.mem\[56\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10242_ _04908_ _00795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11543__A2 _05690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10452__I _05029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10173_ _04864_ _04865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_78_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09018__I data_in_trans\[4\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08547__I0 _03810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11484__S _05683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10354__I0 _04902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06707__C1 u2.mem\[181\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12814_ _00693_ clknet_leaf_186_clock u2.mem\[43\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09889__S _04683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10106__I0 _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08793__S _03990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12634__CLK clknet_leaf_115_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12745_ _00624_ clknet_leaf_44_clock u2.mem\[38\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11854__I0 _05913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12676_ _00555_ clknet_leaf_83_clock u2.mem\[34\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11627_ _05773_ _01315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12784__CLK clknet_leaf_336_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06238__A1 u2.mem\[147\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06238__B2 u2.mem\[169\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11558_ _04333_ _05729_ _05730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_128_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07001__I _02372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06789__A2 _02260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11659__S _05788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10509_ _05072_ _05073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_144_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_203_clock_I clknet_5_31_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11489_ _05687_ _01263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12014__CLK clknet_leaf_315_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11909__I1 _03532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13228_ _01107_ clknet_leaf_298_clock u2.mem\[141\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07738__A1 _01962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13159_ _01038_ clknet_leaf_280_clock u2.mem\[130\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10593__I0 _05126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08538__I0 _03801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11394__S _05625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07720_ u2.mem\[57\]\[10\] _03137_ _03138_ u2.mem\[41\]\[10\] _03189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10345__I0 _04893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07671__I _02566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07651_ _03115_ _03118_ _03119_ _03120_ _03121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_81_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07910__A1 u2.mem\[32\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06602_ _02086_ _02087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07582_ _02504_ _03053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09321_ _03629_ _03539_ _03877_ _04333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA_clkbuf_4_14_0_clock_I clknet_3_7_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06533_ _02017_ _02010_ _02018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11845__I0 _05907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08710__I0 _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06477__A1 u2.mem\[194\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09252_ _04293_ _00420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07674__B1 _03069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06464_ u2.mem\[193\]\[8\] _01942_ _01943_ u2.mem\[194\]\[8\] _01949_ _01957_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08203_ _03552_ u2.mem\[3\]\[3\] _03608_ _03612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_2_1__f_clock_a_I clknet_0_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09183_ _04244_ _00400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09415__A1 _04394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06395_ u2.mem\[190\]\[5\] _01702_ _01704_ u2.mem\[194\]\[5\] _01897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06229__A1 u2.mem\[145\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06229__B2 u2.mem\[177\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08134_ _03522_ _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10820__I1 _03517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08065_ _03492_ _03518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07846__I _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07016_ _02494_ _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_150_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12507__CLK clknet_leaf_191_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10272__I _04922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06401__B2 u2.mem\[185\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08967_ _04023_ u2.mem\[20\]\[4\] _04102_ _04103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08529__I0 _03830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07918_ _03379_ _03380_ _03381_ _03382_ _03383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_5_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08898_ _04032_ u2.mem\[18\]\[8\] _04061_ _04062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_5_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12657__CLK clknet_leaf_235_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07849_ _02600_ _03316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07901__A1 _03363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06704__A2 _02185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10860_ _05198_ u2.mem\[129\]\[1\] _05287_ _05289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09502__S _04443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09519_ _04456_ _00524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_152_clock_I clknet_5_24_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10791_ _05231_ _05247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_73_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12530_ _00409_ clknet_leaf_178_clock u2.mem\[25\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07665__B1 _03060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12461_ _00340_ clknet_leaf_194_clock u2.mem\[21\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11412_ _05637_ _05638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__12037__CLK clknet_2_2__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07417__B1 _02890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12392_ _00271_ clknet_leaf_140_clock u2.mem\[16\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07968__A1 u2.mem\[14\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11343_ _05594_ _01210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10811__I1 _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11274_ _05551_ _01184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12187__CLK clknet_leaf_266_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11278__I _05513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13013_ _00892_ clknet_leaf_67_clock u2.mem\[55\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10225_ _04895_ u2.mem\[49\]\[4\] _04896_ _04897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10182__I _04864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_12_0_clock clknet_4_6_0_clock clknet_5_12_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__07196__A2 _02669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_77_clock_I clknet_5_8_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10156_ _04806_ u2.mem\[47\]\[10\] _04851_ _04854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold5 u2.mem\[0\]\[9\] net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_10087_ _04813_ u2.mem\[45\]\[13\] _04811_ _04814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09193__I0 _04246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07499__A3 _02970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11942__S _05965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11827__I0 _05864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10989_ _05371_ _01079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12728_ _00607_ clknet_leaf_44_clock u2.mem\[37\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09211__I _04147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12659_ _00538_ clknet_leaf_77_clock u2.mem\[33\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07408__B1 _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06180_ _01686_ _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11389__S _05615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10293__S _04938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_354_clock_I clknet_5_5_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10802__I1 _03491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06092__C1 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10092__I _04614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09870_ _04677_ _00654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08821_ _04009_ _00273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07726__A4 _03194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06395__B1 _01704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08752_ _03913_ u2.mem\[15\]\[4\] _03967_ _03968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09184__I0 _04177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07703_ u2.mem\[16\]\[10\] _03033_ _03034_ u2.mem\[33\]\[10\] _03172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08683_ _03925_ u2.mem\[13\]\[9\] _03923_ _03926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07634_ _02419_ _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06698__A1 u2.mem\[184\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07565_ _02469_ _03036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10468__S _05045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09304_ _04269_ u2.mem\[27\]\[8\] _04323_ _04324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06516_ _01991_ _02000_ _02001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11294__I1 u2.mem\[155\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07496_ u2.mem\[39\]\[6\] _02857_ _02858_ u2.mem\[48\]\[6\] _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__13305__CLK clknet_leaf_376_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09235_ _04281_ u2.mem\[25\]\[13\] _04279_ _04282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06447_ _01923_ _01943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09166_ _04151_ u2.mem\[24\]\[7\] _04231_ _04235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06378_ u2.mem\[174\]\[5\] _01656_ _01658_ u2.mem\[155\]\[5\] _01660_ u2.mem\[181\]\[5\]
+ _01880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_159_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08117_ _03556_ _00022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09097_ _04161_ u2.mem\[22\]\[10\] _04192_ _04195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13455__CLK clknet_leaf_321_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07414__A3 _02886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08048_ data_in_trans\[4\].data_sync _03505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10557__I0 _05101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10010_ _04764_ _00707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09999_ _04757_ _00703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06386__B1 _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06386__C2 _01643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11826__I _05895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06925__A2 _02375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09175__I0 _04164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11961_ _05977_ _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06689__A1 u2.mem\[145\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10912_ _05301_ u2.mem\[132\]\[2\] _05319_ _05322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06689__B2 u2.mem\[168\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11892_ u2.mem\[192\]\[6\] _03512_ _05937_ _05938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07350__A2 _02666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10843_ _05194_ u2.mem\[128\]\[0\] _05278_ _05279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10378__S _04989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07638__B1 _03028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13562_ _01441_ clknet_leaf_32_clock u2.mem\[193\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10774_ _05204_ u2.mem\[62\]\[4\] _05237_ _05238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12513_ _00392_ clknet_leaf_175_clock u2.mem\[24\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13493_ _01372_ clknet_leaf_309_clock u2.mem\[185\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12444_ _00323_ clknet_leaf_187_clock u2.mem\[20\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06861__A1 row_select_trans\[0\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08989__I0 _04046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12375_ _00254_ clknet_leaf_138_clock u2.mem\[15\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10905__I _05275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11002__S _05372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10796__I0 _05227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11326_ _05582_ _01205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06613__A1 _02006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06323__C _01826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11257_ _05540_ _01178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10208_ _04884_ _00785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11188_ _05495_ _01154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10139_ _04844_ _00756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12972__CLK clknet_leaf_223_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09166__I0 _04151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08913__I0 _04048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11672__S _05801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07877__B1 _02501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12202__CLK clknet_leaf_43_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07341__A2 _02659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13328__CLK clknet_leaf_1_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10288__S _04933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06695__A4 _02178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07350_ u2.mem\[61\]\[4\] _02666_ _02667_ u2.mem\[63\]\[4\] _02825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11276__I1 u2.mem\[154\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06301_ _01798_ _01799_ _01800_ _01805_ _01806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_31_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12352__CLK clknet_leaf_161_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07281_ u2.mem\[44\]\[3\] _02656_ _02657_ u2.mem\[42\]\[3\] _02757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__13478__CLK clknet_leaf_307_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09020_ _04139_ _04140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06232_ u2.mem\[144\]\[1\] _01671_ _01673_ u2.mem\[182\]\[1\] _01738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06852__B2 u2.mem\[191\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08780__I mem_address_trans\[5\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06163_ _01612_ _01635_ _01670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10787__I0 _05218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06094_ _01600_ _01587_ _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_100_clock_I clknet_5_10_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09922_ _04712_ u2.mem\[41\]\[13\] _04710_ _04713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10539__I0 _05023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09853_ _04583_ u2.mem\[40\]\[5\] _04666_ _04668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_8_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08221__S _03618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06368__B1 _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08804_ _03989_ _04000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09784_ _04617_ _04628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_22_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06996_ _02473_ _02422_ _02423_ _02474_ _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09157__I0 _04136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08735_ _03934_ u2.mem\[14\]\[13\] _03956_ _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08020__I mem_address_trans\[0\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11582__S _05738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08904__I0 _04039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08666_ _03904_ _03914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08955__I _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09321__A3 _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09052__S _04155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07332__A2 _02650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07617_ _03078_ _03081_ _03084_ _03087_ _03088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08597_ _03823_ u2.mem\[11\]\[11\] _03866_ _03870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09987__S _04750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07548_ _02384_ _03019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_25_clock_I clknet_5_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11267__I1 u2.mem\[154\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08891__S _04056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07479_ _02936_ _02941_ _02946_ _02951_ _02952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_14_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10926__S _05327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09218_ _04251_ _04270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_33_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10490_ _05011_ u2.mem\[55\]\[8\] _05061_ _05062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12845__CLK clknet_leaf_214_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09149_ _04224_ _04122_ _04225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10725__I _05195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10778__I0 _05209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07399__A2 _02871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12160_ _00039_ clknet_leaf_236_clock u2.mem\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11111_ _05448_ _01124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06071__A2 _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12995__CLK clknet_leaf_31_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12091_ net23 clknet_2_2__leaf_clock_a inverter_select_trans.A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10661__S _05162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11042_ _05405_ _01098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12225__CLK clknet_leaf_242_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09026__I _04144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_302_clock_I clknet_5_21_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12993_ _00872_ clknet_leaf_253_clock u2.mem\[54\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11492__S _05682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08865__I _03708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11944_ _05225_ u2.mem\[193\]\[13\] _05965_ _05967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10702__I0 _05121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11875_ _03485_ _05926_ _05927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_2974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10826_ u2.mem\[63\]\[11\] _03524_ _05263_ _05267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11258__I1 u2.mem\[153\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07087__A1 _02522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10757_ _03716_ _05227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13545_ _01424_ clknet_leaf_40_clock u2.mem\[192\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07626__A3 _03095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09871__I1 u2.mem\[40\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09696__I _04117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13476_ _01355_ clknet_leaf_309_clock u2.mem\[182\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_173_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10688_ _05108_ u2.mem\[60\]\[6\] _05179_ _05182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_173_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12427_ _00306_ clknet_leaf_190_clock u2.mem\[19\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10769__I0 _05200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12358_ _00237_ clknet_leaf_92_clock u2.mem\[14\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11430__I1 u2.mem\[164\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08105__I _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07929__A4 _03393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11309_ _05554_ u2.mem\[156\]\[4\] _05567_ _05573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13000__CLK clknet_leaf_338_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12289_ _00168_ clknet_leaf_179_clock u2.mem\[10\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_343_clock clknet_5_7_0_clock clknet_leaf_343_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_122_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06850_ u2.mem\[185\]\[5\] _02120_ _02122_ u2.mem\[173\]\[5\] _02330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08976__S _04107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09139__I0 _04167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13150__CLK clknet_leaf_281_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06781_ u2.mem\[150\]\[3\] _02047_ _02034_ u2.mem\[174\]\[3\] u2.mem\[181\]\[3\]
+ _02038_ _02263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_23_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08520_ _03824_ _00157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11497__I1 u2.mem\[168\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_358_clock clknet_5_5_0_clock clknet_leaf_358_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_24_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08451_ _03780_ _00132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07402_ u2.mem\[1\]\[5\] _02797_ _02798_ u2.mem\[7\]\[5\] _02876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_91_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08382_ _03692_ u2.mem\[6\]\[8\] _03737_ _03738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_199_clock_I clknet_5_31_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07333_ _02475_ _02808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09862__I1 u2.mem\[40\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06825__A1 u2.mem\[171\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06286__C1 _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07264_ _01772_ _02361_ _02719_ _02740_ _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09003_ data_in_trans\[1\].data_sync _04126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06215_ _01721_ _01722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10545__I _04986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07195_ u2.mem\[57\]\[1\] _02671_ _02672_ u2.mem\[41\]\[1\] _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06146_ _01607_ _01630_ _01653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11421__I1 u2.mem\[163\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_251_clock_I clknet_5_19_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10481__S _05056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07250__B2 u2.mem\[25\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06077_ col_select_trans\[2\].data_sync _01584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12248__CLK clknet_leaf_56_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09905_ _04682_ _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_119_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11185__I0 _05464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09836_ _04657_ _00640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08886__S _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10932__I0 _05307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06979_ _02405_ _02391_ _02416_ _02458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_86_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09767_ _04565_ u2.mem\[38\]\[0\] _04618_ _04619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12398__CLK clknet_leaf_191_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08718_ _03948_ _00231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08685__I _03700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07803__B _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09698_ _04121_ _04542_ _04566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11488__I1 u2.mem\[167\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07305__A2 _02694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06108__A3 _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09550__I0 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08649_ _03748_ _03876_ _03901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11660_ _05793_ _01328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10611_ _05106_ u2.mem\[58\]\[5\] _05136_ _05138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_74_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11591_ _05667_ _05750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09853__I1 u2.mem\[40\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13330_ _01209_ clknet_leaf_1_clock u2.mem\[158\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06933__I _02386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10542_ _05091_ _00912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13261_ _01140_ clknet_leaf_286_clock u2.mem\[147\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10473_ _05052_ _00882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12212_ _00091_ clknet_leaf_72_clock u2.mem\[5\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13192_ _01071_ clknet_leaf_293_clock u2.mem\[135\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_163_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10376__A1 _04121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12143_ _00022_ clknet_leaf_239_clock u2.mem\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09369__I0 _04362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07792__A2 _03254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13173__CLK clknet_leaf_278_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12074_ data_in_trans\[12\].A clknet_leaf_362_clock data_in_trans\[12\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11025_ _05394_ _05395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_46_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07544__A2 _03005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08741__A1 _03480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06752__B1 _02157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12976_ _00855_ clknet_leaf_264_clock u2.mem\[53\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11927_ _05957_ _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11858_ _05916_ _01403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07004__I _02482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10809_ _05257_ _01013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11100__I0 _05432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11789_ _05873_ _01377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13528_ _01407_ clknet_leaf_332_clock u2.mem\[191\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_146_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07075__A4 _02442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08009__B1 _03462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10365__I _04965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07480__A1 u2.mem\[61\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13459_ _01338_ clknet_leaf_362_clock u2.mem\[180\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_173_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06000_ u2.driver_mem\[3\] _01508_ _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11403__I1 u2.mem\[162\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13516__CLK clknet_leaf_347_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11397__S _05625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08280__I0 _03656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_282_clock clknet_5_22_0_clock clknet_leaf_282_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_99_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07951_ _01976_ _03250_ _03394_ _03415_ _01491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_101_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11196__I _05499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06902_ _02380_ _02381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_64_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12540__CLK clknet_leaf_198_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07882_ u2.mem\[14\]\[13\] _02521_ _02525_ u2.mem\[12\]\[13\] _03348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_64_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10914__I0 _05303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06338__A3 _01828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09621_ _04072_ _04441_ _04521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09780__I0 _04586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06833_ u2.mem\[180\]\[5\] _02042_ _02013_ u2.mem\[172\]\[5\] _02313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_297_clock clknet_5_21_0_clock clknet_leaf_297_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_37_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09552_ _04147_ _04478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06764_ u2.mem\[194\]\[3\] _02198_ _02199_ u2.mem\[190\]\[3\] _02246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08503_ _03812_ u2.mem\[9\]\[6\] _03808_ _03813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12690__CLK clknet_leaf_157_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07299__A1 u2.mem\[52\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09483_ _04384_ u2.mem\[31\]\[12\] _04434_ _04435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06695_ _02172_ _02173_ _02175_ _02178_ _02179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_24_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_220_clock clknet_5_29_0_clock clknet_leaf_220_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08434_ _03769_ _00126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08365_ _03728_ _00098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10476__S _05051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13046__CLK clknet_leaf_33_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07849__I _02600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07316_ u2.mem\[40\]\[4\] _02789_ _02790_ u2.mem\[30\]\[4\] _02791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08296_ _03672_ _00085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11642__I1 u2.mem\[177\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_235_clock clknet_5_25_0_clock clknet_leaf_235_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06274__A2 _01778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07247_ _02720_ _02721_ _02722_ _02723_ _02724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_118_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09599__I0 _04478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12070__CLK clknet_leaf_379_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13196__CLK clknet_leaf_293_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07178_ _02513_ _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_145_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06129_ _01552_ _01635_ _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06026__A2 _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11100__S _05434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11158__I0 _05466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09771__I0 _04573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09819_ _04589_ u2.mem\[39\]\[7\] _04644_ _04648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12830_ _00709_ clknet_leaf_208_clock u2.mem\[44\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06928__I _02346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09523__I0 _04384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12761_ _00640_ clknet_leaf_51_clock u2.mem\[39\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11330__I0 _05583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11770__S _05857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11712_ _05824_ _01349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12692_ _00571_ clknet_leaf_84_clock u2.mem\[35\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11643_ _05782_ _01322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10386__S _04989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06663__I _02147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11574_ _05707_ u2.mem\[173\]\[0\] _05739_ _05740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12413__CLK clknet_leaf_193_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07057__A4 _02474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput17 data_in_a[4] net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput28 mem_address_a[4] net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_122_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07462__A1 u2.mem\[27\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10525_ _05009_ u2.mem\[56\]\[7\] _05078_ _05082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13313_ _01192_ clknet_leaf_365_clock u2.mem\[155\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput39 row_select_a[2] net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__06265__A2 _01755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06804__A4 _02284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13244_ _01123_ clknet_leaf_295_clock u2.mem\[144\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10456_ _05042_ _00875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11397__I0 _05627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12563__CLK clknet_leaf_112_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13175_ _01054_ clknet_leaf_280_clock u2.mem\[132\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10387_ _04996_ _00852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11010__S _05382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12126_ _01467_ clknet_leaf_349_clock u2.driver_mem\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_147_clock_I clknet_5_13_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12057_ net17 clknet_2_0__leaf_clock_a data_in_trans\[4\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07517__A2 _02986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11008_ _05383_ _01086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09214__I _04150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09514__I0 _04375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12959_ _00838_ clknet_leaf_168_clock u2.mem\[52\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11321__I0 _05552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13069__CLK clknet_leaf_274_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11680__S _05800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06480_ u2.mem\[0\]\[12\] _01969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12093__CLK clknet_leaf_380_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08150_ _03534_ _03579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11624__I1 u2.mem\[176\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07048__A4 _02454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07101_ _02579_ _02580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06256__A2 _01759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08081_ _01969_ _03526_ _03529_ _00013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_31_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12906__CLK clknet_leaf_52_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07032_ _02373_ _02511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_162_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07756__A2 _03125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08983_ _04111_ _00333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07934_ _03395_ _03396_ _03397_ _03398_ _03399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_29_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09325__S _04336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07865_ _01969_ _03250_ _03290_ _03331_ _01489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11560__I0 _05707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09604_ _04482_ u2.mem\[34\]\[8\] _04511_ _04512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06816_ u2.mem\[153\]\[4\] _02196_ _02200_ u2.mem\[160\]\[4\] _02297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07796_ _02456_ _03263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09505__I0 _04366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_349_clock_I clknet_5_6_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09535_ _04466_ _00530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06747_ _02227_ _02228_ _02229_ _02230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_52_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09466_ _04425_ _00502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_169_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06678_ _02049_ _02074_ _02113_ _02162_ _02163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__12436__CLK clknet_leaf_102_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07692__A1 u2.mem\[6\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08417_ _03680_ u2.mem\[7\]\[5\] _03758_ _03760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09397_ _04163_ _04382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07579__I _02527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_174_clock clknet_5_27_0_clock clknet_leaf_174_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_127_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08348_ _03714_ u2.mem\[5\]\[13\] _03710_ _03715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07444__B2 u2.mem\[24\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12586__CLK clknet_leaf_117_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08279_ _03658_ _03659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_165_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10310_ _04895_ u2.mem\[51\]\[4\] _04949_ _04950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11290_ _05550_ u2.mem\[155\]\[2\] _05559_ _05562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11379__I0 _05583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_189_clock clknet_5_30_0_clock clknet_leaf_189_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_152_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10241_ _04907_ u2.mem\[49\]\[9\] _04905_ _04908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_65_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10051__I0 _04788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10172_ _03982_ _04863_ _04864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_112_clock clknet_5_11_0_clock clknet_leaf_112_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10354__I1 u2.mem\[52\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11551__I0 _05715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13211__CLK clknet_leaf_301_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06183__A1 u2.mem\[170\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09034__I _04150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06183__B2 u2.mem\[156\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_127_clock clknet_5_15_0_clock clknet_leaf_127_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12813_ _00692_ clknet_leaf_206_clock u2.mem\[43\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11303__I0 _05548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12744_ _00623_ clknet_leaf_43_clock u2.mem\[38\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_163_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13361__CLK clknet_leaf_369_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06486__A2 _01933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12675_ _00554_ clknet_leaf_62_clock u2.mem\[34\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12929__CLK clknet_leaf_151_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_73_clock_I clknet_5_8_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11626_ _05750_ u2.mem\[176\]\[1\] _05771_ _05773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06238__A2 _01676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11557_ _05605_ _05729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_141_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10508_ _04224_ _05071_ _05072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11488_ _05674_ u2.mem\[167\]\[3\] _05683_ _05687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10990__A1 _04249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13227_ _01106_ clknet_leaf_300_clock u2.mem\[141\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10439_ _04995_ u2.mem\[54\]\[2\] _05030_ _05033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07199__B1 _02676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07738__A2 _03017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_298_clock_I clknet_5_21_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13158_ _01037_ clknet_leaf_260_clock u2.mem\[129\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10593__I1 u2.mem\[57\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12109_ _01492_ clknet_leaf_48_clock u2.active_mem\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13089_ _00968_ clknet_leaf_257_clock u2.mem\[60\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09145__S _04218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10345__I1 u2.mem\[52\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07650_ u2.mem\[58\]\[9\] _03044_ _03045_ u2.mem\[36\]\[9\] _03120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_93_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06174__A1 _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12459__CLK clknet_leaf_188_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06601_ _02023_ _02033_ _02086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_350_clock_I clknet_5_4_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07581_ u2.mem\[49\]\[8\] _03050_ _03051_ u2.mem\[46\]\[8\] _03052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_168_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09320_ _04332_ _00449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09879__I _04682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06532_ _02016_ _01986_ _02017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_146_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07123__B1 _02601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07269__A4 _02744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_91_clock clknet_5_10_0_clock clknet_leaf_91_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09251_ _04256_ u2.mem\[26\]\[2\] _04290_ _04293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_167_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06477__A2 _01946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06463_ u2.mem\[192\]\[8\] _01931_ _01956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08202_ _03611_ _00052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09182_ _04174_ u2.mem\[24\]\[14\] _04241_ _04244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06394_ _01888_ _01889_ _01890_ _01895_ _01896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_147_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08133_ _03567_ _00027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06229__A2 _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08064_ data_in_trans\[8\].data_sync _03517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08224__S _03623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07015_ _02477_ _02479_ _02481_ _02424_ _02494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__08226__I0 _03575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07729__A2 _03082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13234__CLK clknet_leaf_289_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06401__A2 _01719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08966_ _04096_ _04102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input31_I mem_address_a[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07917_ u2.mem\[3\]\[14\] _03269_ _03215_ _03382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_25_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08897_ _04050_ _04061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_leaf_44_clock clknet_5_6_0_clock clknet_leaf_44_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07848_ _02598_ _03315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06165__A1 _01665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13384__CLK clknet_leaf_318_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07779_ u2.mem\[6\]\[11\] _03160_ _03161_ u2.mem\[47\]\[11\] _03247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_71_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09518_ _04380_ u2.mem\[32\]\[10\] _04453_ _04456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_59_clock clknet_5_12_0_clock clknet_leaf_59_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10790_ _05246_ _01005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09449_ _04414_ _00496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10728__I _05004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07665__B2 u2.mem\[62\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12460_ _00339_ clknet_leaf_195_clock u2.mem\[21\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11411_ _04071_ _05606_ _05637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_137_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12391_ _00270_ clknet_leaf_140_clock u2.mem\[16\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07968__A2 _02521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11342_ _05593_ u2.mem\[158\]\[4\] _05584_ _05594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06941__I _02419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08090__A1 _01980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11559__I _05730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08217__I0 _03566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11273_ _05550_ u2.mem\[154\]\[2\] _05546_ _05551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08917__A1 _04072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09029__I data_in_trans\[6\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09965__I0 _04716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10224_ _04886_ _04896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_13012_ _00891_ clknet_leaf_69_clock u2.mem\[55\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11772__I0 _05835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10155_ _04853_ _00763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09717__I0 _04579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12601__CLK clknet_leaf_135_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10086_ _04608_ _04813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_169_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06156__A1 _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12751__CLK clknet_leaf_247_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09699__I _04566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11827__I1 u2.mem\[189\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10988_ _05352_ u2.mem\[136\]\[5\] _05364_ _05371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06459__A2 _01942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12727_ _00606_ clknet_leaf_45_clock u2.mem\[37\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08108__I _03499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12658_ _00537_ clknet_leaf_235_clock u2.mem\[33\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11609_ _05762_ _01308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10574__S _05113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12589_ _00468_ clknet_leaf_205_clock u2.mem\[29\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08081__A1 _01969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07423__A4 _02896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11469__I _05673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08208__I0 _03557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06092__C2 u2.mem\[161\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13257__CLK clknet_leaf_286_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06631__A2 _02046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09956__I0 _04707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06919__B1 _02397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07187__A3 _02655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08820_ _03938_ u2.mem\[16\]\[15\] _04005_ _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06395__B2 u2.mem\[194\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09708__I0 _04573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08751_ _03961_ _03967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_6_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11515__I0 _05671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07702_ u2.mem\[1\]\[10\] _03030_ _03031_ u2.mem\[7\]\[10\] _03171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08682_ _03696_ _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07633_ u2.mem\[40\]\[9\] _03022_ _03023_ u2.mem\[30\]\[9\] _03103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06698__A2 _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11932__I _05949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07564_ u2.mem\[16\]\[8\] _03033_ _03034_ u2.mem\[33\]\[8\] _03035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_41_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08219__S _03618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11999__CLK clknet_leaf_18_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09303_ _04312_ _04323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_94_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06515_ _01985_ _01986_ _02000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07495_ u2.mem\[5\]\[6\] _02922_ _02923_ u2.mem\[38\]\[6\] _02968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_55_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09234_ _04170_ _04281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06446_ _01927_ _01942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08018__I _03478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09165_ _04234_ _00392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06377_ u2.mem\[189\]\[5\] _01649_ _01652_ u2.mem\[176\]\[5\] u2.mem\[172\]\[5\]
+ _01653_ _01879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_147_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10254__I0 _04916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08116_ _03554_ u2.mem\[1\]\[4\] _03555_ _03556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07857__I _02618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09096_ _04194_ _00363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08072__A1 _03522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06083__B1 _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08047_ _03488_ _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08889__S _04056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09947__I0 _04698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11754__I0 _05831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_21_clock_I clknet_5_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08688__I _03704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09998_ _04712_ u2.mem\[43\]\[13\] _04755_ _04757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07592__I _02538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06386__B2 u2.mem\[165\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08949_ _04091_ _00319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12774__CLK clknet_leaf_76_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11960_ _05911_ u2.mem\[194\]\[3\] _05975_ _05977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07335__B1 _02809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10911_ _05321_ _01051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10659__S _05162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11891_ _05928_ _05937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_clkbuf_leaf_246_clock_I clknet_5_18_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10842_ _05277_ _05278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__12004__CLK clknet_leaf_41_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08129__S _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09312__I _04312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08686__I0 _03927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13561_ _01440_ clknet_leaf_32_clock u2.mem\[193\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10773_ _05231_ _05237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_12512_ _00391_ clknet_leaf_176_clock u2.mem\[24\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13492_ _01371_ clknet_leaf_307_clock u2.mem\[185\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12154__CLK clknet_leaf_57_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12443_ _00322_ clknet_leaf_185_clock u2.mem\[20\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06861__A2 row_select_trans\[2\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06671__I _02155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12374_ _00253_ clknet_leaf_81_clock u2.mem\[15\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11325_ _05556_ u2.mem\[157\]\[5\] _05575_ _05582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06613__A2 _02080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09938__I0 _04689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11256_ _05508_ u2.mem\[153\]\[2\] _05537_ _05540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_4_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11745__I0 _05837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10207_ _04817_ u2.mem\[48\]\[15\] _04880_ _04884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10921__I _05326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11187_ _05466_ u2.mem\[149\]\[2\] _05492_ _05495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06377__A1 u2.mem\[189\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06377__B2 u2.mem\[176\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10138_ _04788_ u2.mem\[47\]\[2\] _04841_ _04844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11953__S _05972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10069_ _04591_ _04801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06129__A1 _01552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09423__S _04396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06300_ u2.mem\[147\]\[2\] _01676_ _01680_ u2.mem\[169\]\[2\] _01804_ _01805_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_91_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07280_ _02752_ _02753_ _02754_ _02755_ _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_31_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06301__A1 _01798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06231_ u2.mem\[158\]\[1\] _01728_ _01729_ u2.mem\[151\]\[1\] _01736_ _01737_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06852__A2 _02150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06162_ _01655_ _01662_ _01668_ _01669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06581__I _02065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10936__A1 _04180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11984__I0 _05227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10787__I1 u2.mem\[62\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07801__A1 u2.mem\[16\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06093_ _01546_ _01560_ _01600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09892__I _04682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09921_ _04608_ _04712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09852_ _04667_ _00646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_195_clock_I clknet_5_31_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06368__A1 u2.mem\[191\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06368__B2 u2.mem\[179\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08803_ _03999_ _00265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06907__A3 _02353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09783_ _04627_ _00617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06995_ _02428_ _02441_ _02381_ _02474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11863__S _05918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08734_ _03957_ _00238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12027__CLK clknet_2_2__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07317__B1 _02639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07868__A1 u2.mem\[40\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08665_ _03674_ _03913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07868__B2 u2.mem\[30\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07616_ u2.mem\[18\]\[8\] _03085_ _03086_ u2.mem\[19\]\[8\] _03087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_121_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08596_ _03869_ _00188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07547_ u2.mem\[45\]\[8\] _02866_ _02867_ u2.mem\[34\]\[8\] _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07478_ _02947_ _02948_ _02949_ _02950_ _02951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_14_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09217_ _04153_ _04269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06429_ _01918_ _01929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08045__A1 _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09093__I0 _04154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09148_ _04223_ _04224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09079_ _04132_ u2.mem\[22\]\[2\] _04182_ _04185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_159_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10942__S _05337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11110_ _05426_ u2.mem\[144\]\[2\] _05445_ _05448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12090_ output_active_trans.A clknet_leaf_305_clock output_active_trans.data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_162_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08412__S _03753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11041_ _05380_ u2.mem\[140\]\[0\] _05404_ _05405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_2_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10741__I _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07308__B1 _02762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11104__A1 _03486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12992_ _00871_ clknet_leaf_256_clock u2.mem\[54\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11943_ _05966_ _01438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06666__I _02150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11874_ _03477_ _03984_ _05925_ _05926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09042__I data_in_trans\[9\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10825_ _05266_ _01020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09977__I _04739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10466__I0 _05025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13544_ _01423_ clknet_leaf_31_clock u2.mem\[192\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10756_ _05226_ _00991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13475_ _01354_ clknet_leaf_311_clock u2.mem\[182\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10687_ _05181_ _00967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10218__I0 _04891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11013__S _05382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12426_ _00305_ clknet_leaf_121_clock u2.mem\[18\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09084__I0 _04140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11948__S _05965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08831__I0 _04017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12357_ _00236_ clknet_leaf_95_clock u2.mem\[14\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06598__A1 u2.mem\[165\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06598__B2 u2.mem\[163\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11308_ _05572_ _01197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08322__S _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12288_ _00167_ clknet_leaf_179_clock u2.mem\[10\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11747__I _05768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11239_ _05530_ _01170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07547__B1 _02867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09217__I _04153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_171_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08121__I _03512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06780_ u2.mem\[155\]\[3\] _02029_ _02262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06770__A1 u2.mem\[167\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09153__S _04226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06770__B2 u2.mem\[183\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08898__I0 _04032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13445__CLK clknet_leaf_352_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08450_ _03667_ u2.mem\[8\]\[2\] _03777_ _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07401_ u2.mem\[15\]\[5\] _02794_ _02795_ u2.mem\[13\]\[5\] _02875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08381_ _03726_ _03737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_56_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10457__I0 _05016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07332_ u2.mem\[54\]\[4\] _02650_ _02651_ u2.mem\[55\]\[4\] _02807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07617__A4 _03087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06286__B1 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07263_ _02724_ _02729_ _02734_ _02739_ _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__06286__C2 u2.mem\[168\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06825__A2 _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09002_ _04125_ _00338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06214_ _01678_ _01582_ _01614_ _01721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__09075__I0 _04119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07194_ _02549_ _02672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06145_ _01651_ _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07250__A2 _02572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06076_ _01582_ _01576_ _01583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11709__I0 _05796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09904_ _04591_ _04700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11185__I1 u2.mem\[149\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09835_ _04612_ u2.mem\[39\]\[14\] _04654_ _04657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08031__I _03487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08966__I _04096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09766_ _04617_ _04618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06978_ _02456_ _02457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08717_ _03916_ u2.mem\[14\]\[5\] _03946_ _03948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08889__I0 _04023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09697_ _04564_ _04565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09998__S _04755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10002__S _04755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08648_ _03724_ _03481_ _03900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06513__A1 row_select_trans\[5\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12812__CLK clknet_leaf_207_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08579_ _03805_ u2.mem\[11\]\[3\] _03856_ _03860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10448__I0 _05007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10610_ _05137_ _00934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11590_ _05749_ _01302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10541_ _05025_ u2.mem\[56\]\[14\] _05088_ _05091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06277__C2 u2.mem\[181\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12962__CLK clknet_leaf_168_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13260_ _01139_ clknet_leaf_311_clock u2.mem\[146\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10472_ _04987_ u2.mem\[55\]\[0\] _05051_ _05052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07110__I _02347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11948__I0 _05229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12211_ _00090_ clknet_leaf_68_clock u2.mem\[5\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11768__S _05857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13191_ _01070_ clknet_leaf_296_clock u2.mem\[135\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07777__B1 _03091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10620__I0 _05115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12142_ _00021_ clknet_leaf_230_clock u2.mem\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13318__CLK clknet_leaf_318_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07241__A2 _02715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08142__S _03573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_0_clock_a clock_a clknet_0_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_155_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10471__I _05050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12073_ net10 clknet_2_0__leaf_clock_a data_in_trans\[12\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07529__B1 _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09037__I data_in_trans\[8\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11024_ _04311_ _05363_ _05394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_46_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12342__CLK clknet_leaf_92_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07544__A3 _03010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13468__CLK clknet_leaf_360_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06752__A1 u2.mem\[146\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06752__B2 u2.mem\[186\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12975_ _00854_ clknet_leaf_254_clock u2.mem\[53\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11926_ _05915_ u2.mem\[193\]\[5\] _05955_ _05957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12492__CLK clknet_leaf_197_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07701__B1 _03028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11857_ _05915_ u2.mem\[190\]\[5\] _05904_ _05916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10847__S _05278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_143_clock_I clknet_5_13_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10439__I0 _04995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10808_ u2.mem\[63\]\[3\] _03502_ _05253_ _05257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11788_ _05872_ u2.mem\[186\]\[3\] _05866_ _05873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13527_ _01406_ clknet_leaf_325_clock u2.mem\[191\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10739_ _05213_ u2.mem\[61\]\[8\] _05214_ _05215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09057__I0 _04167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13458_ _01337_ clknet_leaf_325_clock u2.mem\[179\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07480__A2 _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07020__I _02498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11939__I0 _05220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11678__S _05801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12409_ _00288_ clknet_leaf_124_clock u2.mem\[17\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13389_ _01268_ clknet_leaf_372_clock u2.mem\[168\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07768__B1 _03072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10611__I0 _05106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07232__A2 _02647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07950_ _03399_ _03404_ _03409_ _03414_ _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_155_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06901_ _02355_ _02379_ _02380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_68_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_68_clock_I clknet_5_9_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07881_ u2.mem\[44\]\[13\] _02514_ _02518_ u2.mem\[42\]\[13\] _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_25_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09620_ _04520_ _00561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06338__A4 _01841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08786__I _03989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06832_ u2.mem\[176\]\[5\] _02003_ _02020_ u2.mem\[189\]\[5\] _02312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07690__I _02621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07940__B1 _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12835__CLK clknet_leaf_113_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09551_ _04477_ _00535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06763_ u2.mem\[154\]\[3\] _02225_ _02226_ u2.mem\[162\]\[3\] _02245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_71_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08502_ _03683_ _03812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07299__A2 _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09482_ _04418_ _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06694_ u2.mem\[149\]\[1\] _02176_ _02177_ u2.mem\[175\]\[1\] _02178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_97_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08433_ _03709_ u2.mem\[7\]\[12\] _03768_ _03769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12985__CLK clknet_leaf_50_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08364_ _03656_ u2.mem\[6\]\[0\] _03727_ _03728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_123_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09410__I _04176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06259__B1 _01708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07315_ _02409_ _02790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10556__I _04997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08295_ _03671_ u2.mem\[5\]\[3\] _03659_ _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09048__I0 _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12215__CLK clknet_leaf_43_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07246_ u2.mem\[57\]\[2\] _02671_ _02672_ u2.mem\[41\]\[2\] _02723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_165_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10492__S _05061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07177_ _02649_ _02652_ _02653_ _02654_ _02655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA_clkbuf_leaf_345_clock_I clknet_5_7_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06128_ _01548_ _01585_ _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10602__I0 _05097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07223__A2 _02385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06059_ _01556_ _01566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11158__I1 u2.mem\[147\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09818_ _04647_ _00632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06734__A1 u2.mem\[159\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06734__B2 u2.mem\[149\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09749_ _04604_ _04605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09523__I1 u2.mem\[32\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12760_ _00639_ clknet_leaf_52_clock u2.mem\[39\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11330__I1 u2.mem\[158\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11711_ _05798_ u2.mem\[181\]\[5\] _05817_ _05824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12691_ _00570_ clknet_leaf_61_clock u2.mem\[35\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11850__I _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06944__I _02373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11642_ _05752_ u2.mem\[177\]\[2\] _05779_ _05782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11573_ _05738_ _05739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_leaf_342_clock clknet_5_7_0_clock clknet_leaf_342_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_161_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput18 data_in_a[5] net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_11_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13312_ _01191_ clknet_leaf_363_clock u2.mem\[155\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10524_ _05081_ _00904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput29 mem_address_a[5] net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_168_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07462__A2 _02871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06265__A3 _01762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13243_ _01122_ clknet_leaf_289_clock u2.mem\[144\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10455_ _05014_ u2.mem\[54\]\[9\] _05040_ _05042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11397__I1 u2.mem\[162\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_357_clock clknet_5_5_0_clock clknet_leaf_357_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_139_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13174_ _01053_ clknet_leaf_279_clock u2.mem\[132\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10386_ _04995_ u2.mem\[53\]\[2\] _04989_ _04996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12125_ _01466_ clknet_leaf_349_clock u2.driver_mem\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12858__CLK clknet_leaf_143_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08600__S _03871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12056_ data_in_trans\[3\].A clknet_leaf_376_clock data_in_trans\[3\].data_sync vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07517__A3 _02987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11007_ _05380_ u2.mem\[138\]\[0\] _05382_ _05383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06725__A1 u2.mem\[184\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09514__I1 u2.mem\[32\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12958_ _00837_ clknet_leaf_197_clock u2.mem\[52\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11321__I1 u2.mem\[157\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11909_ u2.mem\[192\]\[14\] _03532_ _05928_ _05947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10577__S _05113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12889_ _00768_ clknet_leaf_52_clock u2.mem\[47\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_294_clock_I clknet_5_21_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09278__I0 _04283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12238__CLK clknet_leaf_230_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09230__I _04166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07100_ _02439_ _02440_ _02512_ _02408_ _02579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_9_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08080_ _03527_ _03528_ _03529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_173_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07031_ _02369_ _02510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__12388__CLK clknet_leaf_79_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07685__I _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09450__I0 _04391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08982_ _04039_ u2.mem\[20\]\[11\] _04107_ _04111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09606__S _04511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09202__I0 _04258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07933_ u2.mem\[57\]\[14\] _02548_ _02550_ u2.mem\[41\]\[14\] _03398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08510__S _03817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10899__I0 _05303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07864_ _03299_ _03310_ _03321_ _03330_ _03331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_29_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09603_ _04500_ _04511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__11560__I1 u2.mem\[172\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06815_ u2.mem\[194\]\[4\] _02198_ _02199_ u2.mem\[190\]\[4\] _02296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07795_ u2.mem\[15\]\[12\] _03260_ _03261_ u2.mem\[13\]\[12\] _03262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09505__I1 u2.mem\[32\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09534_ _04463_ u2.mem\[33\]\[0\] _04465_ _04466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06746_ u2.mem\[148\]\[2\] _02128_ _02130_ u2.mem\[152\]\[2\] _02229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09465_ _04366_ u2.mem\[31\]\[4\] _04424_ _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10487__S _05056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06677_ _02118_ _02124_ _02140_ _02161_ _02162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_145_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08416_ _03759_ _00118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09269__I0 _04274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09396_ _04381_ _00476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07692__A2 _03160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08347_ _03713_ _03714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08278_ _03657_ _03544_ _03632_ _03658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_165_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07229_ u2.mem\[16\]\[2\] _02465_ _02467_ u2.mem\[33\]\[2\] _02706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11379__I1 u2.mem\[161\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10240_ _04595_ _04907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09441__I0 _04382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06404__B1 _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10171_ _04862_ _04863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10950__S _05337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09516__S _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06939__I _02407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06707__A1 u2.mem\[155\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11551__I1 u2.mem\[171\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07380__A1 _02845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12812_ _00691_ clknet_leaf_207_clock u2.mem\[43\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09251__S _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11303__I1 u2.mem\[156\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13506__CLK clknet_leaf_333_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12743_ _00622_ clknet_leaf_43_clock u2.mem\[38\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08180__I0 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12674_ _00553_ clknet_leaf_153_clock u2.mem\[34\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_281_clock clknet_5_23_0_clock clknet_leaf_281_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_16_clock_I clknet_5_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09050__I data_in_trans\[11\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11625_ _05772_ _01314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12530__CLK clknet_leaf_178_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11556_ _05728_ _01289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10507_ _04862_ _05071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_296_clock clknet_5_21_0_clock clknet_leaf_296_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06789__A4 _02270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11487_ _05686_ _01262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05997__A2 row_col_select_trans.data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13226_ _01105_ clknet_leaf_299_clock u2.mem\[141\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09432__I0 _04373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10438_ _05032_ _00867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07199__A1 u2.mem\[26\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13157_ _01036_ clknet_leaf_285_clock u2.mem\[129\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10860__S _05287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10369_ _04983_ _00847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06946__A1 _02421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12108_ _01491_ clknet_leaf_48_clock u2.active_mem\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13088_ _00967_ clknet_leaf_258_clock u2.mem\[60\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13036__CLK clknet_leaf_276_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12039_ net2 clknet_2_2__leaf_clock_a col_select_trans\[1\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_152_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_234_clock clknet_5_28_0_clock clknet_leaf_234_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_20_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11691__S _05810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06600_ _02084_ _02085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07580_ _02531_ _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12060__CLK clknet_leaf_375_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13186__CLK clknet_leaf_293_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06531_ _01984_ _02016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_94_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08171__I0 _03559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09250_ _04292_ _00419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_249_clock clknet_5_18_0_clock clknet_leaf_249_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_33_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06462_ _01914_ _01955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07674__A2 _03068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08201_ _03550_ u2.mem\[3\]\[2\] _03608_ _03611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11058__I0 _05384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09181_ _04243_ _00399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06393_ u2.mem\[166\]\[5\] _01592_ _01598_ u2.mem\[161\]\[5\] _01894_ _01895_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_30_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08132_ _03566_ u2.mem\[1\]\[9\] _03564_ _03567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08063_ _03488_ _03516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07014_ _02492_ _02493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08304__I _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09423__I0 _04364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08965_ _04101_ _00325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07916_ u2.mem\[16\]\[14\] _03266_ _03267_ u2.mem\[33\]\[14\] _03381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_25_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06952__A4 _02430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08896_ _04060_ _00297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12403__CLK clknet_leaf_109_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input24_I mem_address_a[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13529__CLK clknet_leaf_332_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07847_ u2.mem\[17\]\[12\] _03312_ _03313_ u2.mem\[24\]\[12\] _03314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_17_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06165__A2 _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07901__A3 _03365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07778_ u2.mem\[8\]\[11\] _03093_ _03094_ u2.mem\[4\]\[11\] _03246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09517_ _04455_ _00523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06729_ u2.mem\[176\]\[2\] _02003_ _02020_ u2.mem\[189\]\[2\] _02212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12553__CLK clknet_leaf_123_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08162__I0 _03550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11106__S _05445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09448_ _04389_ u2.mem\[30\]\[14\] _04411_ _04414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07665__A2 _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11049__I0 _05390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09379_ _04369_ u2.mem\[29\]\[5\] _04367_ _04370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11410_ _05636_ _01235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07417__A2 _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12390_ _00269_ clknet_leaf_81_clock u2.mem\[16\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11341_ _05513_ _05593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10744__I _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08214__I _03607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11272_ _05507_ _05550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_152_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_242_clock_I clknet_5_25_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13011_ _00890_ clknet_leaf_30_clock u2.mem\[55\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13059__CLK clknet_leaf_31_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10223_ _04578_ _04895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_152_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11772__I1 u2.mem\[185\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10154_ _04804_ u2.mem\[47\]\[9\] _04851_ _04853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07274__B _02749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10085_ _04812_ _00734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12083__CLK clknet_leaf_381_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06156__A2 _01618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11288__I0 _05548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10987_ _05370_ _01078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11016__S _05382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12726_ _00605_ clknet_leaf_24_clock u2.mem\[37\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12657_ _00536_ clknet_leaf_235_clock u2.mem\[33\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11608_ _05746_ u2.mem\[175\]\[0\] _05761_ _05762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07408__A2 _02880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12588_ _00467_ clknet_leaf_205_clock u2.mem\[29\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11539_ _05718_ _01282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10654__I _05151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09405__I0 _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06092__B2 u2.mem\[149\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08124__I _03514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13209_ _01088_ clknet_leaf_300_clock u2.mem\[138\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11912__A1 _01981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12426__CLK clknet_leaf_121_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07187__A4 _02664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06395__A2 _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08750_ _03966_ _00245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06579__I _02056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_173_clock clknet_5_26_0_clock clknet_leaf_173_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11515__I1 u2.mem\[169\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07701_ u2.mem\[15\]\[10\] _03027_ _03028_ u2.mem\[13\]\[10\] _03170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_6_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08681_ _03924_ _00218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12576__CLK clknet_leaf_184_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07632_ u2.mem\[32\]\[9\] _03019_ _03020_ u2.mem\[2\]\[9\] _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_65_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11279__I0 _05554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_188_clock clknet_5_30_0_clock clknet_leaf_188_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07563_ _02466_ _03034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09302_ _04322_ _00441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06514_ _01998_ _01999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07494_ _02963_ _02964_ _02965_ _02966_ _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA_clkbuf_leaf_191_clock_I clknet_5_30_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09233_ _04280_ _00414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06855__B1 _02143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06445_ u2.mem\[192\]\[5\] _01931_ _01941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10765__S _05232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_111_clock clknet_5_11_0_clock clknet_leaf_111_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_124_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09164_ _04148_ u2.mem\[24\]\[6\] _04231_ _04234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06376_ _01877_ _01878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08115_ _03545_ _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09095_ _04158_ u2.mem\[22\]\[9\] _04192_ _04194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13201__CLK clknet_leaf_295_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08072__A2 _03518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06083__A1 u2.mem\[177\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06083__B2 u2.mem\[168\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08046_ _01809_ _03489_ _03503_ _00004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_126_clock clknet_5_15_0_clock clknet_leaf_126_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_163_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11203__I0 _05505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11754__I1 u2.mem\[184\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13351__CLK clknet_leaf_377_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09997_ _04756_ _00702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06386__A2 _01583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08948_ _04044_ u2.mem\[19\]\[13\] _04089_ _04091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12919__CLK clknet_leaf_134_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08879_ _04050_ _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_3825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10910_ _05299_ u2.mem\[132\]\[1\] _05319_ _05321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07886__A2 _03341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11890_ _05936_ _01415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10841_ _03982_ _05276_ _05277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08135__I0 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07099__B1 _02577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13560_ _01439_ clknet_leaf_32_clock u2.mem\[193\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07638__A2 _03027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10772_ _05236_ _00997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09883__I0 _04685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12511_ _00390_ clknet_leaf_176_clock u2.mem\[24\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06846__B1 _02137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13491_ _01370_ clknet_leaf_307_clock u2.mem\[185\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10675__S _05174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12442_ _00321_ clknet_leaf_120_clock u2.mem\[19\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08145__S _03573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11442__I0 _05623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12373_ _00252_ clknet_leaf_80_clock u2.mem\[15\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12449__CLK clknet_leaf_169_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07271__B1 _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11324_ _05581_ _01204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11255_ _05539_ _01177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08879__I _04050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07783__I _02360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11745__I1 u2.mem\[183\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10206_ _04883_ _00784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07023__B1 _02501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_90_clock clknet_5_10_0_clock clknet_leaf_90_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_80_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11186_ _05494_ _01153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06377__A2 _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12599__CLK clknet_leaf_115_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10137_ _04843_ _00755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09704__S _04567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10068_ _04800_ _00729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06129__A2 _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07877__A2 _02499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12709_ _00588_ clknet_leaf_64_clock u2.mem\[36\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06301__A2 _01799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06230_ _01730_ _01733_ _01735_ _01736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_43_clock clknet_5_6_0_clock clknet_leaf_43_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10384__I _04130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06161_ u2.mem\[180\]\[0\] _01664_ _01667_ u2.mem\[150\]\[0\] _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_157_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06065__A1 _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06092_ u2.mem\[166\]\[0\] _01592_ _01595_ u2.mem\[149\]\[0\] _01598_ u2.mem\[161\]\[0\]
+ _01599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__13374__CLK clknet_leaf_369_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09920_ _04711_ _00670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_58_clock clknet_5_12_0_clock clknet_leaf_58_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_138_clock_I clknet_5_14_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09851_ _04579_ u2.mem\[40\]\[4\] _04666_ _04667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06368__A2 _01681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08802_ _03920_ u2.mem\[16\]\[7\] _03995_ _03999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09782_ _04589_ u2.mem\[38\]\[7\] _04623_ _04627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06994_ _02346_ _02473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_26_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08733_ _03931_ u2.mem\[14\]\[12\] _03956_ _03957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07317__A1 u2.mem\[27\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08664_ _03912_ _00213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07615_ _02605_ _03086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10872__A1 _05295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10559__I _05000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08595_ _03821_ u2.mem\[11\]\[10\] _03866_ _03869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07546_ _02360_ _03017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08029__I data_in_trans\[0\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11672__I0 _05786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07477_ u2.mem\[43\]\[6\] _02820_ _02821_ u2.mem\[20\]\[6\] _02950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_10_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09216_ _04268_ _00409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06428_ _01927_ _01928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09617__I0 _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09147_ _03628_ _03748_ _03774_ _04223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__07089__B _02485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06359_ _01854_ _01855_ _01856_ _01861_ _01862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_135_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07253__B1 _02683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09078_ _04184_ _00355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08029_ data_in_trans\[0\].data_sync _03490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12741__CLK clknet_leaf_24_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07005__B1 _02483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11040_ _05403_ _05404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_46_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07108__I _02412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12891__CLK clknet_leaf_224_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12991_ _00870_ clknet_leaf_254_clock u2.mem\[54\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07308__A1 _01808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11853__I _03673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07308__B2 _02783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11942_ _05222_ u2.mem\[193\]\[12\] _05965_ _05966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06947__I _02425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10163__I0 _04813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11873_ _03985_ _03986_ _05925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13247__CLK clknet_leaf_288_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12121__CLK clknet_leaf_348_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10824_ u2.mem\[63\]\[10\] _03522_ _05263_ _05266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13543_ _01422_ clknet_leaf_40_clock u2.mem\[192\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10755_ _05225_ u2.mem\[61\]\[13\] _05223_ _05226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_40_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06295__A1 u2.mem\[173\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09608__I0 _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06295__B2 u2.mem\[185\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13474_ _01353_ clknet_leaf_308_clock u2.mem\[182\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13397__CLK clknet_leaf_327_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10686_ _05106_ u2.mem\[60\]\[5\] _05179_ _05181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12425_ _00304_ clknet_leaf_120_clock u2.mem\[18\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10218__I1 u2.mem\[49\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11415__I0 _05627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07244__B1 _02544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12356_ _00235_ clknet_leaf_93_clock u2.mem\[14\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11307_ _05552_ u2.mem\[156\]\[3\] _05568_ _05572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_5_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12287_ _00166_ clknet_leaf_178_clock u2.mem\[10\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11989__CLK clknet_leaf_335_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11238_ _05500_ u2.mem\[152\]\[0\] _05529_ _05530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_150_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08595__I0 _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11964__S _05975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11169_ _05460_ u2.mem\[148\]\[0\] _05484_ _05485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10154__I0 _04804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07400_ _02868_ _02869_ _02870_ _02873_ _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_91_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08380_ _03736_ _00105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12614__CLK clknet_leaf_92_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07331_ u2.mem\[50\]\[4\] _02647_ _02648_ u2.mem\[51\]\[4\] _02806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_91_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_64_clock_I clknet_5_9_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06286__A1 u2.mem\[158\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07262_ _02735_ _02736_ _02737_ _02738_ _02739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06286__B2 u2.mem\[151\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07483__B1 _02905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09001_ _04119_ u2.mem\[21\]\[0\] _04124_ _04125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11406__I0 _05633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06213_ _01719_ _01720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07193_ _02547_ _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12764__CLK clknet_leaf_220_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07235__B1 _02490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06144_ _01582_ _01635_ _01651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08513__S _03817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06589__A2 _02063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06075_ _01581_ _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_289_clock_I clknet_5_21_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09903_ _04699_ _00665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06033__S _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08586__I0 _03812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09834_ _04656_ _00639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06210__A1 _01706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09765_ _04180_ _04542_ _04617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06977_ _02412_ _02413_ _02454_ _02455_ _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__12144__CLK clknet_leaf_230_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06761__A2 _02241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08716_ _03947_ _00230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09696_ _04117_ _04564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10145__I0 _04795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_341_clock_I clknet_5_7_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08647_ _03655_ _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06513__A2 _01997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12294__CLK clknet_leaf_99_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08578_ _03859_ _00180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_168_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07529_ u2.mem\[26\]\[7\] _02908_ _02909_ u2.mem\[10\]\[7\] _03001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_25_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08510__I0 _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07598__I _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11114__S _05444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06277__A1 u2.mem\[174\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07474__B1 _02890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10540_ _05090_ _00911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06277__B2 u2.mem\[155\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10471_ _05050_ _05051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_109_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12210_ _00089_ clknet_leaf_252_clock u2.mem\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13190_ _01069_ clknet_leaf_297_clock u2.mem\[135\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12141_ _00020_ clknet_leaf_231_clock u2.mem\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10620__I1 u2.mem\[58\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12072_ data_in_trans\[11\].A clknet_leaf_379_clock data_in_trans\[11\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08577__I0 _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11023_ _05393_ _01091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06737__C1 u2.mem\[145\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06752__A2 _02155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10136__I0 _04786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12974_ _00853_ clknet_leaf_271_clock u2.mem\[53\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12637__CLK clknet_leaf_214_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11925_ _05956_ _01430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07701__A1 u2.mem\[15\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11856_ _03678_ _05915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10807_ _05256_ _01012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09454__A1 _04417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11787_ _03669_ _05872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12787__CLK clknet_leaf_31_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13526_ _01405_ clknet_leaf_327_clock u2.mem\[191\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10738_ _05195_ _05214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_9_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08009__A2 _03461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13457_ _01336_ clknet_leaf_325_clock u2.mem\[179\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10669_ _05170_ _00960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12017__CLK clknet_2_3__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12408_ _00287_ clknet_leaf_124_clock u2.mem\[17\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11939__I1 u2.mem\[193\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13388_ _01267_ clknet_leaf_372_clock u2.mem\[168\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12339_ _00218_ clknet_leaf_93_clock u2.mem\[13\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10611__I1 u2.mem\[58\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_290_clock_I clknet_5_21_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06440__A1 _01809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06440__B2 _01937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12167__CLK clknet_leaf_62_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06900_ _02352_ _02341_ _02342_ _02378_ _02379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_151_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07880_ _03342_ _03343_ _03344_ _03345_ _03346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06728__C1 u2.mem\[181\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06831_ u2.mem\[155\]\[5\] _02029_ _02034_ u2.mem\[174\]\[5\] u2.mem\[181\]\[5\]
+ _02038_ _02311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_68_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09550_ _04476_ u2.mem\[33\]\[5\] _04474_ _04477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10103__S _04820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06587__I _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06762_ u2.mem\[166\]\[3\] _02097_ _02099_ u2.mem\[161\]\[3\] _02243_ _02244_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08501_ _03811_ _00151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13562__CLK clknet_leaf_32_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09481_ _04433_ _00509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06693_ _02105_ _02177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08432_ _03752_ _03768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_91_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08363_ _03726_ _03727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10837__I mem_address_trans\[6\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07314_ _02402_ _02789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06259__A1 u2.mem\[152\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06259__B2 u2.mem\[153\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08294_ _03670_ _03671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07211__I _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07245_ u2.mem\[37\]\[2\] _02537_ _02539_ u2.mem\[59\]\[2\] _02722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07208__B1 _02601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07176_ u2.mem\[58\]\[1\] _02487_ _02490_ u2.mem\[36\]\[1\] _02654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08243__S _03634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06127_ _01633_ _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10572__I _03690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10602__I1 u2.mem\[58\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09138__I _04202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06431__A1 _01727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06058_ _01557_ _01561_ _01564_ _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13092__CLK clknet_leaf_26_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10366__I0 _04913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09817_ _04586_ u2.mem\[39\]\[6\] _04644_ _04647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06734__A2 _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07931__A1 u2.mem\[60\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10013__S _04762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09748_ data_in_trans\[12\].data_sync _04604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09679_ _04482_ u2.mem\[36\]\[8\] _04554_ _04555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11710_ _05823_ _01348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12690_ _00569_ clknet_leaf_157_clock u2.mem\[35\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07695__B1 _03131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06498__B2 _01980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11641_ _05781_ _01321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11618__I0 _05758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10747__I _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11572_ _05411_ _05729_ _05738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_161_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13311_ _01190_ clknet_leaf_363_clock u2.mem\[155\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11779__S _05866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10523_ _05007_ u2.mem\[56\]\[6\] _05078_ _05081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput19 data_in_a[6] net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_17_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09249__S _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06670__A1 _02022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13242_ _01121_ clknet_leaf_287_clock u2.mem\[143\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06960__I _02386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10454_ _05041_ _00874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08798__I0 _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13173_ _01052_ clknet_leaf_278_clock u2.mem\[132\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10385_ _04994_ _04995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12124_ _01465_ clknet_leaf_37_clock u2.driver_mem\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_174_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07765__A4 _03232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_12_clock_I clknet_5_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12055_ net16 clknet_2_0__leaf_clock_a data_in_trans\[3\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10357__I0 _04904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11006_ _05381_ _05382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_38_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07922__A1 u2.mem\[58\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07922__B2 u2.mem\[36\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11019__S _05381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09712__S _04567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11857__I0 _05915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12957_ _00836_ clknet_leaf_197_clock u2.mem\[52\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10858__S _05287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_237_clock_I clknet_5_25_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11908_ _05946_ _01423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12888_ _00767_ clknet_leaf_57_clock u2.mem\[47\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11839_ _03654_ _05903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08127__I _03517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11689__S _05810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13509_ _01388_ clknet_leaf_347_clock u2.mem\[188\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_174_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07030_ u2.mem\[43\]\[0\] _02505_ _02508_ u2.mem\[20\]\[0\] _02509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_173_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06870__I _02348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08789__I0 _03907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10392__I _04138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09450__I1 u2.mem\[30\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10596__I0 _05128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07610__B1 _03080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08981_ _04110_ _00332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07932_ u2.mem\[37\]\[14\] _03295_ _03296_ u2.mem\[59\]\[14\] _03397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_138_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10348__I0 _04895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07863_ _03322_ _03325_ _03328_ _03329_ _03330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_96_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07913__A1 _03374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09602_ _04510_ _00553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06814_ u2.mem\[169\]\[4\] _02142_ _02144_ u2.mem\[147\]\[4\] _02294_ _02295_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__12952__CLK clknet_leaf_148_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07794_ _02451_ _03261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09533_ _04464_ _04465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06745_ u2.mem\[153\]\[2\] _02196_ _02200_ u2.mem\[160\]\[2\] _02228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11848__I0 _05909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11951__I _05970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09464_ _04418_ _04424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_24_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06676_ u2.mem\[169\]\[0\] _02142_ _02144_ u2.mem\[147\]\[0\] _02160_ _02161_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_51_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13308__CLK clknet_leaf_369_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08415_ _03675_ u2.mem\[7\]\[4\] _03758_ _03759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09395_ _04380_ u2.mem\[29\]\[10\] _04376_ _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09269__I1 u2.mem\[26\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08346_ _03712_ _03713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12332__CLK clknet_5_28_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08277_ _03540_ _03657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_165_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13458__CLK clknet_leaf_325_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09069__S _04168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07228_ u2.mem\[1\]\[2\] _02457_ _02461_ u2.mem\[7\]\[2\] _02705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06652__A1 _02056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07097__B _02546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07159_ u2.mem\[40\]\[1\] _02403_ _02410_ u2.mem\[30\]\[1\] _02637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10587__I0 _05121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09441__I1 u2.mem\[30\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06404__A1 u2.mem\[146\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12482__CLK clknet_leaf_172_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06404__B2 u2.mem\[186\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10170_ _03985_ _03986_ _04861_ _04862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_160_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10339__I0 _04885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_186_clock_I clknet_5_30_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08952__I0 _04048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12811_ _00690_ clknet_leaf_184_clock u2.mem\[43\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06955__I _02373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12742_ _00621_ clknet_leaf_24_clock u2.mem\[38\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08148__S _03573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12673_ _00552_ clknet_leaf_153_clock u2.mem\[34\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11624_ _05746_ u2.mem\[176\]\[0\] _05771_ _05772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11555_ _05719_ u2.mem\[171\]\[5\] _05721_ _05728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07786__I _02396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10506_ _05070_ _00897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11486_ _05671_ u2.mem\[167\]\[2\] _05683_ _05686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12825__CLK clknet_leaf_129_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13225_ _01104_ clknet_leaf_301_clock u2.mem\[141\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10437_ _04992_ u2.mem\[54\]\[1\] _05030_ _05032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_48_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09432__I1 u2.mem\[30\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07199__A2 _02675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13156_ _01035_ clknet_leaf_283_clock u2.mem\[129\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10368_ _04916_ u2.mem\[52\]\[13\] _04981_ _04983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06946__A2 _02422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12107_ _01490_ clknet_leaf_47_clock u2.active_mem\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10940__I _04126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13087_ _00966_ clknet_5_19_0_clock u2.mem\[60\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10299_ _04072_ _04863_ _04943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09196__I0 _04254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12038_ col_select_trans\[0\].A clknet_leaf_316_clock col_select_trans\[0\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08943__I0 _04039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07026__I _02504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12205__CLK clknet_leaf_267_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06530_ _02014_ _02015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07659__B1 _03054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07123__A2 _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06461_ u2.mem\[0\]\[8\] _01954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08200_ _03610_ _00051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09180_ _04171_ u2.mem\[24\]\[13\] _04241_ _04243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_18_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06392_ _01891_ _01892_ _01893_ _01894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08131_ _03520_ _03566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08062_ _01951_ _03504_ _03515_ _00008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07831__B1 _03138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07977__A4 _03440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07013_ _02473_ _02370_ _02374_ _02393_ _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__09423__I1 u2.mem\[30\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09617__S _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06105__I _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06937__A2 _02415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08964_ _04021_ u2.mem\[20\]\[3\] _04097_ _04101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_25_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09416__I _04395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07915_ u2.mem\[1\]\[14\] _03263_ _03264_ u2.mem\[7\]\[14\] _03380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_102_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08320__I _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08895_ _04030_ u2.mem\[18\]\[7\] _04056_ _04060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08934__I0 _04030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_341_clock clknet_5_7_0_clock clknet_leaf_341_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_56_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07846_ _02590_ _03313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_20_0_clock_I clknet_4_10_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09352__S _04351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06165__A3 _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input17_I data_in_a[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13130__CLK clknet_5_6_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07901__A4 _03366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07777_ u2.mem\[39\]\[11\] _03090_ _03091_ u2.mem\[48\]\[11\] _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_44_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09516_ _04378_ u2.mem\[32\]\[9\] _04453_ _04455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06728_ u2.mem\[155\]\[2\] _02030_ _02035_ u2.mem\[174\]\[2\] u2.mem\[181\]\[2\]
+ _02039_ _02211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_37_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09447_ _04413_ _00495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06659_ _02143_ _02144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_169_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13280__CLK clknet_leaf_380_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09378_ _04144_ _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08329_ data_in_trans\[10\].data_sync _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11122__S _05453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11340_ _05592_ _01209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06625__A1 u2.mem\[159\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06625__B2 u2.mem\[149\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06443__C _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11271_ _05549_ _01183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13010_ _00889_ clknet_leaf_251_clock u2.mem\[55\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_165_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09527__S _04458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10222_ _04894_ _00789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06389__B1 _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11856__I _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10153_ _04852_ _00762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10760__I _03720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09178__I0 _04167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12228__CLK clknet_leaf_73_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10980__I0 _05340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10084_ _04810_ u2.mem\[45\]\[12\] _04811_ _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_309_clock clknet_5_20_0_clock clknet_leaf_309_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09878__A1 _04249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08925__I0 _04021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11685__A1 _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10732__I0 _05209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12378__CLK clknet_leaf_60_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11591__I _05667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11288__I1 u2.mem\[155\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10986_ _05349_ u2.mem\[136\]\[4\] _05364_ _05370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07105__A2 _02570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12725_ _00604_ clknet_leaf_24_clock u2.mem\[37\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08606__S _03871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12656_ _00535_ clknet_leaf_235_clock u2.mem\[33\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06864__B2 row_select_trans\[1\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09102__I0 _04167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10935__I _05334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11607_ _05760_ _05761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_12587_ _00466_ clknet_leaf_205_clock u2.mem\[29\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09802__A1 _03751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11032__S _05395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06616__A1 _01992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08405__I _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11538_ _05717_ u2.mem\[170\]\[4\] _05708_ _05718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_128_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11967__S _05980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06092__A2 _01592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13003__CLK clknet_leaf_266_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11469_ _05673_ _05674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09437__S _04406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13208_ _01087_ clknet_leaf_297_clock u2.mem\[138\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06919__A2 _02385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11912__A2 _05929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13139_ _01018_ clknet_leaf_34_clock u2.mem\[63\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09169__I0 _04154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input9_I data_in_a[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13153__CLK clknet_leaf_283_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08140__I _03527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07700_ _03165_ _03166_ _03167_ _03168_ _03169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_66_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08680_ _03922_ u2.mem\[13\]\[8\] _03923_ _03924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07631_ u2.mem\[45\]\[9\] _03099_ _03100_ u2.mem\[34\]\[9\] _03101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11207__S _05502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07562_ _02464_ _03033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11279__I1 u2.mem\[154\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09301_ _04267_ u2.mem\[27\]\[7\] _04318_ _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06513_ row_select_trans\[5\].data_sync _01997_ _01998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07493_ u2.mem\[18\]\[6\] _02852_ _02853_ u2.mem\[19\]\[6\] _02966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_146_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_134_clock_I clknet_5_15_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11006__I _05381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09232_ _04278_ u2.mem\[25\]\[12\] _04279_ _04280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_146_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06444_ _01844_ _01938_ _01939_ _01940_ _01468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_107_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06855__B2 u2.mem\[147\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08516__S _03817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09163_ _04233_ _00391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06375_ u2.mem\[0\]\[5\] _01877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_148_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08114_ _03506_ _03554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09094_ _04193_ _00362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08315__I _03687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06083__A2 _01583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08045_ _03502_ _03493_ _03503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09347__S _04346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11203__I1 u2.mem\[150\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09996_ _04709_ u2.mem\[43\]\[12\] _04755_ _04756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_280_clock clknet_5_23_0_clock clknet_leaf_280_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_59_clock_I clknet_5_12_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08050__I _03492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08947_ _04090_ _00318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06791__B1 _02244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08907__I0 _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12520__CLK clknet_leaf_124_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08878_ _03583_ _03988_ _04050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07829_ _02538_ _03296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07886__A3 _03346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_295_clock clknet_5_21_0_clock clknet_leaf_295_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_72_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10840_ _05275_ _05276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12670__CLK clknet_leaf_217_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09810__S _04639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10771_ _05202_ u2.mem\[62\]\[3\] _05232_ _05236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12510_ _00389_ clknet_leaf_193_clock u2.mem\[24\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13490_ _01369_ clknet_leaf_307_clock u2.mem\[185\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12441_ _00320_ clknet_leaf_119_clock u2.mem\[19\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13026__CLK clknet_leaf_265_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12372_ _00251_ clknet_leaf_79_clock u2.mem\[15\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11442__I1 u2.mem\[165\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_233_clock clknet_5_28_0_clock clknet_leaf_233_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_165_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11323_ _05554_ u2.mem\[157\]\[4\] _05575_ _05581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_336_clock_I clknet_5_18_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11254_ _05505_ u2.mem\[153\]\[1\] _05537_ _05539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10205_ _04815_ u2.mem\[48\]\[14\] _04880_ _04883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_79_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11185_ _05464_ u2.mem\[149\]\[1\] _05492_ _05494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_248_clock clknet_5_18_0_clock clknet_leaf_248_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_45_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09056__I _04123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10136_ _04786_ u2.mem\[47\]\[1\] _04841_ _04843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06782__B1 _02019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10067_ _04799_ u2.mem\[45\]\[7\] _04793_ _04800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10866__S _05286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08826__A2 _04013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11130__I0 _05432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10969_ _05346_ u2.mem\[135\]\[3\] _05356_ _05360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_43_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06837__A1 u2.mem\[159\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12708_ _00587_ clknet_leaf_69_clock u2.mem\[36\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06837__B2 u2.mem\[149\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12639_ _00518_ clknet_leaf_159_clock u2.mem\[32\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06160_ _01666_ _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13519__CLK clknet_leaf_13_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11697__S _05809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06065__A2 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06091_ _01576_ _01597_ _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_172_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11496__I _05691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12543__CLK clknet_leaf_189_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09850_ _04660_ _04666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08801_ _03998_ _00264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_60_clock_I clknet_5_12_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06993_ _02453_ _02462_ _02468_ _02471_ _02472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09781_ _04626_ _00616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08732_ _03940_ _03956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_6_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07317__A2 _02638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12693__CLK clknet_leaf_82_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08663_ _03911_ u2.mem\[13\]\[3\] _03905_ _03912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07614_ _02603_ _03085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08594_ _03868_ _00187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07545_ _01951_ _02784_ _02995_ _03016_ _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_39_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10776__S _05237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13049__CLK clknet_leaf_343_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_12_0_clock clknet_3_6_0_clock clknet_4_12_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_34_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_285_clock_I clknet_5_20_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06828__A1 u2.mem\[184\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07476_ u2.mem\[49\]\[6\] _02817_ _02818_ u2.mem\[46\]\[6\] _02949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11672__I1 u2.mem\[179\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09215_ _04267_ u2.mem\[25\]\[7\] _04261_ _04268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06427_ _01916_ _01927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09146_ _04222_ _00385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12073__CLK clknet_2_0__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13199__CLK clknet_leaf_292_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06358_ u2.mem\[166\]\[4\] _01757_ _01758_ u2.mem\[161\]\[4\] _01860_ _01861_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_135_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07089__C _02562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06056__A2 col_select_trans\[1\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09077_ _04128_ u2.mem\[22\]\[1\] _04182_ _04184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_162_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06289_ u2.mem\[190\]\[2\] _01703_ _01705_ u2.mem\[194\]\[2\] _01794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11400__S _05625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09077__S _04182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08028_ _03488_ _03489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10016__S _04767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09979_ _04746_ _00694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12990_ _00869_ clknet_leaf_275_clock u2.mem\[54\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09553__I0 _04478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11941_ _05949_ _05965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_3645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10163__I1 u2.mem\[47\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11872_ _05924_ _01409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09540__S _04465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10823_ _05265_ _01019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10686__S _05179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06819__A1 u2.mem\[154\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13542_ _01421_ clknet_leaf_18_clock u2.mem\[192\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10754_ _03712_ _05225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07492__A1 u2.mem\[52\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13473_ _01352_ clknet_leaf_308_clock u2.mem\[182\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10685_ _05180_ _00966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_172_clock clknet_5_26_0_clock clknet_leaf_172_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_12_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12424_ _00303_ clknet_leaf_121_clock u2.mem\[18\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11415__I1 u2.mem\[163\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12355_ _00234_ clknet_leaf_91_clock u2.mem\[14\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07794__I _02451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11306_ _05571_ _01196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12286_ _00165_ clknet_leaf_199_clock u2.mem\[10\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11179__I0 _05472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_187_clock clknet_5_30_0_clock clknet_leaf_187_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_153_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11237_ _05528_ _05529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_150_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10926__I0 _05301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07547__A2 _02866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06203__I _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11168_ _05483_ _05484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_110_clock clknet_5_11_0_clock clknet_leaf_110_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10119_ _04806_ u2.mem\[46\]\[10\] _04830_ _04833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11099_ _05440_ _01120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11351__I0 _05587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11980__S _05985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07180__B1 _02657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_125_clock clknet_5_15_0_clock clknet_leaf_125_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_23_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07330_ _02796_ _02799_ _02802_ _02804_ _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12096__CLK clknet_leaf_246_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06873__I _02340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13341__CLK clknet_leaf_1_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07261_ u2.mem\[6\]\[2\] _02694_ _02695_ u2.mem\[47\]\[2\] _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06286__A2 _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09000_ _04123_ _04124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__12909__CLK clknet_leaf_202_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06212_ _01613_ _01614_ _01597_ _01719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_121_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06691__C1 u2.mem\[159\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07192_ u2.mem\[37\]\[1\] _02537_ _02539_ u2.mem\[59\]\[1\] _02670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_157_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07235__A1 u2.mem\[58\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06143_ _01649_ _01650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13491__CLK clknet_leaf_307_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10090__I0 _04815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06074_ _01580_ _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09902_ _04698_ u2.mem\[41\]\[7\] _04692_ _04699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09625__S _04522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09833_ _04609_ u2.mem\[39\]\[13\] _04654_ _04656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_150_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06746__B1 _02130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09764_ _04616_ _00609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06976_ _02362_ _02455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_39_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08715_ _03913_ u2.mem\[14\]\[4\] _03946_ _03947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09695_ _04563_ _00593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08646_ _03898_ _00209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12439__CLK clknet_leaf_119_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07171__B1 _02648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08577_ _03803_ u2.mem\[11\]\[2\] _03856_ _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07528_ _02996_ _02997_ _02998_ _02999_ _03000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_74_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07459_ u2.mem\[45\]\[6\] _02866_ _02867_ u2.mem\[34\]\[6\] _02932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12589__CLK clknet_leaf_205_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10470_ _03751_ _04964_ _05050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09129_ _04202_ _04213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_159_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11130__S _05452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12140_ _00019_ clknet_leaf_225_clock u2.mem\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07777__A2 _03090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07241__A4 _02717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12071_ net9 clknet_2_0__leaf_clock_a data_in_trans\[11\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10908__I0 _05294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07529__A2 _02908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11022_ _05392_ u2.mem\[138\]\[5\] _05381_ _05393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_77_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06737__C2 _02081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13214__CLK clknet_leaf_297_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08741__A4 _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12973_ _00852_ clknet_leaf_273_clock u2.mem\[53\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_42_clock clknet_5_6_0_clock clknet_leaf_42_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_17_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11333__I0 _05587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11924_ _05913_ u2.mem\[193\]\[4\] _05955_ _05956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07162__B1 _02639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07701__A2 _03027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13364__CLK clknet_leaf_363_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11855_ _05914_ _01402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07789__I _02409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06693__I _02105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10806_ u2.mem\[63\]\[2\] _03499_ _05253_ _05256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_57_clock clknet_5_12_0_clock clknet_leaf_57_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11786_ _05871_ _01376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13525_ _01404_ clknet_leaf_329_clock u2.mem\[191\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10737_ _03690_ _05213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13456_ _01335_ clknet_leaf_320_clock u2.mem\[179\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08614__S _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10668_ _05126_ u2.mem\[59\]\[14\] _05167_ _05170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12407_ _00286_ clknet_leaf_121_clock u2.mem\[17\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13387_ _01266_ clknet_leaf_364_clock u2.mem\[168\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10599_ _05130_ _05131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_115_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07768__A2 _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12338_ _00217_ clknet_leaf_159_clock u2.mem\[13\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_233_clock_I clknet_5_28_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12082__D net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06440__A2 _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12269_ _00148_ clknet_leaf_194_clock u2.mem\[9\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07029__I _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06830_ u2.mem\[150\]\[5\] _02192_ _02310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06868__I _02346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09244__I _04287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07940__A2 _02594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06761_ _02240_ _02241_ _02242_ _02243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_55_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08500_ _03810_ u2.mem\[9\]\[5\] _03808_ _03811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_64_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09480_ _04382_ u2.mem\[31\]\[11\] _04429_ _04433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06692_ _02109_ _02176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09180__S _04241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08431_ _03767_ _00125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12731__CLK clknet_leaf_266_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11215__S _05501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08362_ _03657_ _03725_ _03632_ _03726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_23_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07313_ u2.mem\[32\]\[4\] _02786_ _02787_ u2.mem\[2\]\[4\] _02788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_71_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08293_ _03669_ _03670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07244_ u2.mem\[60\]\[2\] _02542_ _02544_ u2.mem\[62\]\[2\] _02721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07208__A1 u2.mem\[52\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07175_ u2.mem\[53\]\[1\] _02476_ _02483_ u2.mem\[56\]\[1\] _02653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07759__A2 _03224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08956__A1 _04095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06126_ _01581_ _01609_ _01633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_127_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10763__A1 _04394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11885__S _05932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12111__CLK clknet_leaf_348_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13237__CLK clknet_leaf_302_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06057_ _01563_ _01564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06431__A2 _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11684__I _05768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09816_ _04646_ _00631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12261__CLK clknet_leaf_23_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13387__CLK clknet_leaf_364_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09747_ _04603_ _00605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06959_ _02398_ _02411_ _02427_ _02437_ _02438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__11315__I0 _05544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08993__I data_in_trans\[0\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09678_ _04543_ _04554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_28_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09090__S _04187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08629_ _03878_ _03889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07695__A1 _01958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06498__A2 _01924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11640_ _05750_ u2.mem\[177\]\[1\] _05779_ _05781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_182_clock_I clknet_5_27_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11571_ _05737_ _01295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13310_ _01189_ clknet_leaf_363_clock u2.mem\[155\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10522_ _05080_ _00903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10453_ _05011_ u2.mem\[54\]\[8\] _05040_ _05041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13241_ _01120_ clknet_leaf_288_clock u2.mem\[143\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06670__A2 _02052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10054__I0 _04790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13172_ _01051_ clknet_leaf_278_clock u2.mem\[132\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10384_ _04130_ _04994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06958__B1 _02436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12123_ _01458_ clknet_leaf_37_clock u2.driver_mem\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09265__S _04300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12054_ data_in_trans\[2\].A clknet_leaf_379_clock data_in_trans\[2\].data_sync vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12604__CLK clknet_leaf_216_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11594__I _05670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11005_ _04288_ _05363_ _05381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_120_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06186__A1 _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09064__I _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12754__CLK clknet_leaf_247_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12956_ _00835_ clknet_leaf_197_clock u2.mem\[52\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11907_ u2.mem\[192\]\[13\] _03530_ _05942_ _05946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12887_ _00766_ clknet_leaf_57_clock u2.mem\[47\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11838_ _05902_ _01397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07312__I _02396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07438__B2 u2.mem\[25\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10874__S _05297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11769_ _05860_ _01370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10293__I0 _04916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13508_ _01387_ clknet_leaf_345_clock u2.mem\[188\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06110__A1 _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12134__CLK clknet_leaf_12_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13439_ _01318_ clknet_leaf_353_clock u2.mem\[176\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10045__I0 _04782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_384_clock_I clknet_5_0_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08980_ _04037_ u2.mem\[20\]\[10\] _04107_ _04110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09175__S _04236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09738__I0 _04596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07931_ u2.mem\[60\]\[14\] _03292_ _03293_ u2.mem\[62\]\[14\] _03396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11545__I0 _05707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08410__I0 _03667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07862_ u2.mem\[6\]\[12\] _03160_ _03161_ u2.mem\[47\]\[12\] _03329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_64_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07913__A2 _03375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09601_ _04480_ u2.mem\[34\]\[7\] _04506_ _04510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06813_ _02291_ _02292_ _02293_ _02294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_68_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07793_ _02444_ _03260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11009__I _05339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09532_ _04013_ _04441_ _04464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06744_ u2.mem\[194\]\[2\] _02198_ _02199_ u2.mem\[190\]\[2\] _02227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08519__S _03817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09702__I _04126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09463_ _04423_ _00501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06675_ _02149_ _02154_ _02159_ _02160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_97_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08414_ _03752_ _03758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_12_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08318__I data_in_trans\[8\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09394_ _04160_ _04380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08477__I0 _03718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08345_ data_in_trans\[13\].data_sync _03712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10284__I0 _04907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08276_ _03655_ _03656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07227_ u2.mem\[15\]\[2\] _02445_ _02452_ u2.mem\[13\]\[2\] _02704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06652__A2 _02001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10036__I0 _04712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07158_ u2.mem\[32\]\[1\] _02385_ _02397_ u2.mem\[2\]\[1\] _02636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08053__I data_in_trans\[5\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12627__CLK clknet_leaf_111_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06109_ _01562_ _01574_ _01548_ _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_106_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06404__A2 _01691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07089_ _02560_ _02561_ _02485_ _02562_ _02568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_161_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09729__I0 _04589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_129_clock_I clknet_5_15_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12777__CLK clknet_leaf_147_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06168__A1 _01612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12810_ _00689_ clknet_leaf_130_clock u2.mem\[42\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12007__CLK clknet_2_1__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09612__I _04500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12741_ _00620_ clknet_leaf_24_clock u2.mem\[38\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12672_ _00551_ clknet_leaf_156_clock u2.mem\[34\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08468__I0 _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11623_ _05770_ _05771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10275__I0 _04898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06971__I _02394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08164__S _03585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11554_ _05727_ _01288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10505_ _05027_ u2.mem\[55\]\[15\] _05066_ _05070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06643__A2 _02041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11485_ _05685_ _01261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10027__I0 _04703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09059__I data_in_trans\[13\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13224_ _01103_ clknet_leaf_291_clock u2.mem\[140\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10436_ _05031_ _00866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13552__CLK clknet_leaf_10_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13155_ _01034_ clknet_leaf_281_clock u2.mem\[129\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10367_ _04982_ _00846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12106_ _01489_ clknet_leaf_47_clock u2.active_mem\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10298_ _04942_ _00817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13086_ _00965_ clknet_leaf_274_clock u2.mem\[60\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09196__I1 u2.mem\[25\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12037_ net1 clknet_2_2__leaf_clock_a col_select_trans\[0\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06159__A1 _01612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11152__A1 _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09522__I _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12939_ _00818_ clknet_leaf_225_clock u2.mem\[51\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06460_ _01951_ _01938_ _01952_ _01953_ _01471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_61_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06331__A1 u2.mem\[173\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07042__I _02520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06331__B2 u2.mem\[185\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08459__I0 _03684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06391_ u2.mem\[159\]\[5\] _01603_ _01594_ u2.mem\[149\]\[5\] _01893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_57_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08130_ _03565_ _00026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10266__I0 _04889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06881__I _02359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08084__A1 _01973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08061_ _03514_ _03507_ _03515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_147_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10018__I0 _04694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07012_ u2.mem\[58\]\[0\] _02487_ _02490_ u2.mem\[36\]\[0\] _02491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09959__I0 _04709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11766__I0 _05829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09584__A1 _03583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_130_clock_I clknet_5_15_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08963_ _04100_ _00324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07914_ u2.mem\[15\]\[14\] _03260_ _03261_ u2.mem\[13\]\[14\] _03379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_97_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08894_ _04059_ _00296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07217__I _02623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07845_ _02585_ _03312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07776_ u2.mem\[5\]\[11\] _03155_ _03156_ u2.mem\[38\]\[11\] _03244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_17_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06570__A1 u2.mem\[164\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06570__B2 u2.mem\[178\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09515_ _04454_ _00522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06727_ u2.mem\[150\]\[2\] _02192_ _02210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_24_0_clock_I clknet_4_12_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13425__CLK clknet_leaf_365_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09446_ _04387_ u2.mem\[30\]\[13\] _04411_ _04413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08048__I data_in_trans\[4\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06658_ _02045_ _02077_ _02143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09377_ _04368_ _00470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06589_ _02055_ _02063_ _02069_ _02073_ _02074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_127_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_55_clock_I clknet_5_12_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11403__S _05625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10257__I0 _04918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08328_ _03698_ _00091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08075__A1 _03524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13575__CLK clknet_leaf_33_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08870__I0 _04044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08259_ _03566_ u2.mem\[4\]\[9\] _03644_ _03646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10009__I0 _04685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11202__I _05504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09808__S _04639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08712__S _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11270_ _05548_ u2.mem\[154\]\[1\] _05546_ _05549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10221_ _04893_ u2.mem\[49\]\[3\] _04887_ _04894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06389__A1 u2.mem\[187\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06389__B2 u2.mem\[192\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10152_ _04801_ u2.mem\[47\]\[8\] _04851_ _04852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_160_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10083_ _04783_ _04811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_94_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07127__I _02605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09543__S _04465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09878__A2 _04659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07889__A1 u2.mem\[37\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11685__A2 _05808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10732__I1 u2.mem\[61\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06966__I _02444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09342__I _04335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_332_clock_I clknet_5_18_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08689__I0 _03929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10985_ _05369_ _01077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12724_ _00603_ clknet_leaf_25_clock u2.mem\[37\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06313__A1 u2.mem\[189\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06313__B2 u2.mem\[176\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12655_ _00534_ clknet_leaf_236_clock u2.mem\[33\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07797__I _02460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11606_ _04416_ _05729_ _05760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__08066__A1 _03517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12586_ _00465_ clknet_leaf_117_clock u2.mem\[28\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09802__A2 _04542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11537_ _05676_ _05717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06616__A2 _02001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12942__CLK clknet_leaf_220_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06206__I _01712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11468_ _03501_ _05673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13207_ _01086_ clknet_leaf_300_clock u2.mem\[138\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10419_ _05019_ _00861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07577__B1 _02890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11399_ _05507_ _05629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13138_ _01017_ clknet_leaf_330_clock u2.mem\[63\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12090__D output_active_trans.A vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13069_ _00948_ clknet_leaf_274_clock u2.mem\[59\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12322__CLK clknet_leaf_167_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07630_ _02435_ _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07561_ u2.mem\[1\]\[8\] _03030_ _03031_ u2.mem\[7\]\[8\] _03032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10398__I _05004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09300_ _04321_ _00440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10487__I0 _05009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06512_ row_select_trans\[4\].data_sync _01997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_94_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07492_ u2.mem\[52\]\[6\] _02849_ _02850_ u2.mem\[21\]\[6\] _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12472__CLK clknet_leaf_123_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07501__B1 _02952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09231_ _04251_ _04279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06855__A2 _02141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06443_ u2.mem\[193\]\[4\] _01928_ _01929_ u2.mem\[192\]\[4\] _01934_ _01940_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_166_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11223__S _05520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09162_ _04145_ u2.mem\[24\]\[5\] _04231_ _04233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_159_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06374_ _01844_ _01555_ _01876_ _01484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08113_ _03553_ _00021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07804__A1 _03262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09093_ _04154_ u2.mem\[22\]\[8\] _04192_ _04193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_159_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06116__I _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08044_ _03501_ _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07280__A2 _02753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11739__I0 _05831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11957__I _05971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08604__I0 _03830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07568__B1 _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08331__I _03700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_281_clock_I clknet_5_23_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09995_ _04739_ _04755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08946_ _04041_ u2.mem\[19\]\[12\] _04089_ _04090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_170_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06791__A1 _01809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09363__S _04358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06791__B2 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08877_ _04049_ _00289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07828_ _02536_ _03295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07740__B1 _03020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12815__CLK clknet_leaf_167_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07886__A4 _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07759_ _03223_ _03224_ _03225_ _03226_ _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_25_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07099__A2 _02572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10770_ _05235_ _00996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09429_ _04403_ _00487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06846__A2 _02136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12965__CLK clknet_leaf_105_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12440_ _00319_ clknet_leaf_119_clock u2.mem\[19\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07410__I _02500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11978__I0 _05220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12371_ _00250_ clknet_leaf_80_clock u2.mem\[15\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11322_ _05580_ _01203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10650__I0 _05108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07271__A2 _02457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07566__B _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11253_ _05538_ _01176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10204_ _04882_ _00783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10402__I0 _05007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07023__A2 _02499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11184_ _05493_ _01152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10135_ _04842_ _00754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06782__A1 u2.mem\[176\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06782__B2 u2.mem\[189\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10066_ _04588_ _04799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10212__S _04887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12495__CLK clknet_leaf_176_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09072__I _04179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10968_ _05359_ _01070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11130__I1 u2.mem\[145\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12707_ _00586_ clknet_leaf_65_clock u2.mem\[36\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11043__S _05404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10899_ _05303_ u2.mem\[131\]\[3\] _05310_ _05314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12638_ _00517_ clknet_leaf_215_clock u2.mem\[32\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07320__I _02451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06364__C _01866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11969__I0 _05211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11978__S _05985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_340_clock clknet_5_7_0_clock clknet_leaf_340_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08834__I0 _04019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12569_ _00448_ clknet_leaf_128_clock u2.mem\[27\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10641__I0 _05099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06090_ _01596_ _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_172_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08800_ _03918_ u2.mem\[16\]\[6\] _03995_ _03998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13270__CLK clknet_leaf_5_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09780_ _04586_ u2.mem\[38\]\[6\] _04623_ _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06992_ u2.mem\[3\]\[0\] _02470_ _02359_ _02471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08731_ _03955_ _00237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12838__CLK clknet_leaf_87_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09011__I0 _04132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08662_ _03670_ _03911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07722__B1 _03142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07613_ u2.mem\[52\]\[8\] _03082_ _03083_ u2.mem\[21\]\[8\] _03084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_93_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08593_ _03819_ u2.mem\[11\]\[9\] _03866_ _03868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_121_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12988__CLK clknet_leaf_274_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07544_ _03000_ _03005_ _03010_ _03015_ _03016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA_clkbuf_leaf_228_clock_I clknet_5_28_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09710__I _04134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07475_ u2.mem\[14\]\[6\] _02892_ _02893_ u2.mem\[12\]\[6\] _02948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09214_ _04150_ _04267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12218__CLK clknet_leaf_54_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10880__I0 _05301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06426_ u2.mem\[194\]\[1\] _01924_ _01926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08326__I _03696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_308_clock clknet_5_20_0_clock clknet_leaf_308_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09145_ _04177_ u2.mem\[23\]\[15\] _04218_ _04222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06357_ _01857_ _01858_ _01859_ _01860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10792__S _05247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09358__S _04351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09076_ _04183_ _00354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07253__A2 _02682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06288_ _01789_ _01790_ _01791_ _01792_ _01793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_136_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08027_ _03487_ _03488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07005__A2 _02476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09978_ _04691_ u2.mem\[43\]\[4\] _04745_ _04746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06764__A1 u2.mem\[194\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09093__S _04192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08929_ _04080_ _00310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11128__S _05452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10699__I0 _05119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11940_ _05964_ _01437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07713__B1 _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10967__S _05356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11871_ _05915_ u2.mem\[191\]\[5\] _05917_ _05924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10822_ u2.mem\[63\]\[9\] _03520_ _05263_ _05265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08437__S _03768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11112__I1 u2.mem\[144\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13541_ _01420_ clknet_leaf_18_clock u2.mem\[192\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10753_ _05224_ _00990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09069__I0 _04177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13472_ _01351_ clknet_leaf_308_clock u2.mem\[182\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10684_ _05103_ u2.mem\[60\]\[4\] _05179_ _05180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13143__CLK clknet_leaf_40_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07140__I _02618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12423_ _00302_ clknet_leaf_120_clock u2.mem\[18\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08816__I0 _03934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12354_ _00233_ clknet_leaf_162_clock u2.mem\[14\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07244__A2 _02542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11597__I _05673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11305_ _05550_ u2.mem\[156\]\[2\] _05568_ _05571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13293__CLK clknet_leaf_384_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12285_ _00164_ clknet_leaf_194_clock u2.mem\[10\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11328__A1 _04393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09067__I data_in_trans\[15\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11236_ _04223_ _05527_ _05528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__08900__S _04061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09241__I0 _04285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06204__B1 _01710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10006__I _04761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11167_ _04094_ _05482_ _05483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_67_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_177_clock_I clknet_5_27_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07952__B1 _02436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10118_ _04832_ _00747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11098_ _05430_ u2.mem\[143\]\[4\] _05434_ _05440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_76_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10049_ _04787_ _00723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06507__A1 row_select_trans\[5\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07315__I _02409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11351__I1 u2.mem\[159\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10877__S _05297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07260_ u2.mem\[8\]\[2\] _02610_ _02612_ u2.mem\[4\]\[2\] _02737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10862__I0 _05200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06140__C1 u2.mem\[165\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07483__A2 _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06211_ u2.mem\[154\]\[0\] _01699_ _01701_ u2.mem\[162\]\[0\] _01717_ _01718_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__06691__B1 _02098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07191_ u2.mem\[60\]\[1\] _02542_ _02544_ u2.mem\[62\]\[1\] _02669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08807__I0 _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06691__C2 _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12510__CLK clknet_leaf_193_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11501__S _05692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09178__S _04241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06142_ _01613_ _01622_ _01644_ _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__09480__I0 _04382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07235__A2 _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06443__B1 _01929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_294_clock clknet_5_21_0_clock clknet_leaf_294_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06073_ _01550_ _01579_ _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10117__S _04830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11300__I _05567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09901_ _04588_ _04698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09906__S _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09232__I0 _04278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12660__CLK clknet_leaf_83_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09832_ _04655_ _00638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06746__B2 u2.mem\[152\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09763_ _04615_ u2.mem\[37\]\[15\] _04606_ _04616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06975_ _02428_ _02390_ _02381_ _02454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_100_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13016__CLK clknet_leaf_339_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08714_ _03940_ _03946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_41_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09694_ _04498_ u2.mem\[36\]\[15\] _04559_ _04563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09641__S _04532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11342__I1 u2.mem\[158\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08645_ _03832_ u2.mem\[12\]\[15\] _03894_ _03898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_232_clock clknet_5_28_0_clock clknet_leaf_232_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_26_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10787__S _05242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07710__A3 _03177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08576_ _03858_ _00179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09299__I0 _04265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08257__S _03644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_379_clock_I clknet_5_0_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12040__CLK clknet_leaf_316_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13166__CLK clknet_leaf_277_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_168_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10586__I _05094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07527_ u2.mem\[57\]\[7\] _02904_ _02905_ u2.mem\[41\]\[7\] _02999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_74_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_247_clock clknet_5_18_0_clock clknet_leaf_247_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10853__I0 _05207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07474__A2 _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07458_ _01877_ _02784_ _02898_ _02931_ _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06409_ _01878_ _01554_ _01910_ _01485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__12190__CLK clknet_leaf_267_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07389_ _02856_ _02859_ _02862_ _02863_ _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_109_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11558__A1 _04333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09088__S _04187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09128_ _04212_ _00377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09471__I0 _04373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10027__S _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09059_ data_in_trans\[13\].data_sync _04170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06985__A1 _02412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11210__I _05510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12070_ data_in_trans\[10\].A clknet_leaf_379_clock data_in_trans\[10\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11030__I0 _05386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11021_ _05351_ _05392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06737__A1 u2.mem\[165\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06737__B2 u2.mem\[163\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12972_ _00851_ clknet_leaf_223_clock u2.mem\[53\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11333__I1 u2.mem\[158\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13509__CLK clknet_leaf_347_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11923_ _05949_ _05955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_4199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10697__S _05184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07162__A1 u2.mem\[27\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11854_ _05913_ u2.mem\[190\]\[4\] _05904_ _05914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10805_ _05255_ _01011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11785_ _05870_ u2.mem\[186\]\[2\] _05866_ _05871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12533__CLK clknet_leaf_104_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13524_ _01403_ clknet_leaf_7_clock u2.mem\[190\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10736_ _05212_ _00985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13455_ _01334_ clknet_leaf_321_clock u2.mem\[179\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_174_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10667_ _05169_ _00959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11321__S _05576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12406_ _00285_ clknet_leaf_103_clock u2.mem\[17\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09462__I0 _04364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12683__CLK clknet_leaf_211_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13386_ _01265_ clknet_leaf_323_clock u2.mem\[167\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10598_ _04288_ _05071_ _05130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12337_ _00216_ clknet_leaf_209_clock u2.mem\[13\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12268_ _00147_ clknet_leaf_194_clock u2.mem\[9\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08630__S _03889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13039__CLK clknet_leaf_335_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11219_ _05517_ u2.mem\[150\]\[5\] _05501_ _05518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12199_ _00078_ clknet_leaf_42_clock u2.mem\[4\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06728__A1 u2.mem\[155\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07925__B1 _02525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06728__B2 u2.mem\[174\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06760_ u2.mem\[188\]\[3\] _02185_ _02177_ u2.mem\[175\]\[3\] _02242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12063__CLK clknet_2_1__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06691_ u2.mem\[166\]\[1\] _02096_ _02098_ u2.mem\[161\]\[1\] u2.mem\[159\]\[1\]
+ _02174_ _02175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_58_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07153__A1 _02557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11790__I _03673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08430_ _03705_ u2.mem\[7\]\[11\] _03763_ _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06884__I _02362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_380_clock_I clknet_5_0_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06900__A1 _02352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08361_ _03724_ _03605_ _03725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_75_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07312_ _02396_ _02787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10835__I0 u2.mem\[63\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08292_ _03501_ _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08805__S _04000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06664__B1 _02148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07243_ u2.mem\[61\]\[2\] _02666_ _02667_ u2.mem\[63\]\[2\] _02720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11231__S _05519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07208__A2 _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07174_ u2.mem\[54\]\[1\] _02650_ _02651_ u2.mem\[55\]\[1\] _02652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06125_ _01631_ _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08540__S _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06056_ _01562_ col_select_trans\[1\].data_sync _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_160_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12406__CLK clknet_leaf_103_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09815_ _04583_ u2.mem\[39\]\[5\] _04644_ _04646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06195__A2 _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09746_ _04602_ u2.mem\[37\]\[11\] _04593_ _04603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_171_clock clknet_5_26_0_clock clknet_leaf_171_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06958_ u2.mem\[45\]\[0\] _02432_ _02436_ u2.mem\[34\]\[0\] _02437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11315__I1 u2.mem\[157\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09677_ _04553_ _00585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07144__A1 _02443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06889_ _02365_ _02366_ _02367_ _02368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12556__CLK clknet_leaf_202_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11406__S _05624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08628_ _03888_ _00201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10310__S _04949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07695__A2 _03017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06352__C1 _01732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08559_ _03848_ _00172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_186_clock clknet_5_30_0_clock clknet_leaf_186_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_125_clock_I clknet_5_15_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11205__I _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11570_ _05719_ u2.mem\[172\]\[5\] _05730_ _05737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09692__I0 _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06655__B1 _02127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10521_ _05005_ u2.mem\[56\]\[5\] _05078_ _05080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11141__S _05462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13240_ _01119_ clknet_leaf_289_clock u2.mem\[143\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10452_ _05029_ _05040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_13_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09444__I0 _04384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10980__S _05365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13171_ _01050_ clknet_leaf_281_clock u2.mem\[132\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_163_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10383_ _04993_ _00851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12122_ _01485_ clknet_leaf_343_clock u2.select_mem_col\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_124_clock clknet_5_15_0_clock clknet_leaf_124_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08450__S _03777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12053_ net15 clknet_2_0__leaf_clock_a data_in_trans\[2\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06969__I _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11004_ _05334_ _05380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13331__CLK clknet_leaf_2_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_139_clock clknet_5_12_0_clock clknet_leaf_139_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_120_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12955_ _00834_ clknet_leaf_194_clock u2.mem\[52\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13481__CLK clknet_leaf_306_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11906_ _05945_ _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12886_ _00765_ clknet_leaf_71_clock u2.mem\[47\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11837_ _05876_ u2.mem\[189\]\[5\] _05895_ _05902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09683__I0 _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11768_ _05831_ u2.mem\[185\]\[2\] _05857_ _05860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11490__I0 _05677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13507_ _01386_ clknet_leaf_353_clock u2.mem\[188\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10719_ _05200_ u2.mem\[61\]\[2\] _05196_ _05201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11699_ _04120_ _05808_ _05817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06110__A2 _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11051__S _05403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13438_ _01317_ clknet_leaf_366_clock u2.mem\[176\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09435__I0 _04375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11242__I0 _05508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13369_ _01248_ clknet_leaf_371_clock u2.mem\[165\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06949__A1 _02348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_327_clock_I clknet_5_17_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09456__S _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12429__CLK clknet_leaf_192_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07610__A2 _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07930_ u2.mem\[61\]\[14\] _02553_ _02555_ u2.mem\[63\]\[14\] _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_170_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06879__I _02357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09255__I _04289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11545__I1 u2.mem\[171\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07861_ u2.mem\[8\]\[12\] _03326_ _03327_ u2.mem\[4\]\[12\] _03328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_60_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08410__I1 u2.mem\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12579__CLK clknet_leaf_111_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09600_ _04509_ _00552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06812_ u2.mem\[179\]\[4\] _02151_ _02153_ u2.mem\[191\]\[4\] _02293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07792_ _03251_ _03254_ _03257_ _03258_ _03259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_84_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09531_ _04118_ _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06743_ _02127_ _02226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_97_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09462_ _04364_ u2.mem\[31\]\[3\] _04419_ _04423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10130__S _04835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06674_ u2.mem\[146\]\[0\] _02156_ _02158_ u2.mem\[186\]\[0\] _02159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08413_ _03757_ _00117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09393_ _04379_ _00475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11025__I _05394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10808__I0 u2.mem\[63\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08344_ _03711_ _00094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09674__I0 _04478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10433__A1 _04180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08275_ _03654_ _03655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13204__CLK clknet_leaf_293_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07226_ _02699_ _02700_ _02701_ _02702_ _02703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09426__I0 _04366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08334__I data_in_trans\[11\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11896__S _05937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11233__I0 _05517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_41_clock clknet_5_6_0_clock clknet_leaf_41_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_164_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07157_ u2.mem\[45\]\[1\] _02633_ _02634_ u2.mem\[34\]\[1\] _02635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_3_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09366__S _04358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06108_ _01612_ _01613_ _01614_ _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_65_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13354__CLK clknet_leaf_377_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07088_ _02566_ _02567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_154_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06039_ col_select_trans\[0\].data_sync col_select_trans\[1\].data_sync _01546_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10305__S _04944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_56_clock clknet_5_12_0_clock clknet_leaf_56_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_59_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_51_clock_I clknet_5_13_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06168__A2 _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07365__B2 u2.mem\[25\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09729_ _04589_ u2.mem\[37\]\[7\] _04580_ _04590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07380__A4 _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10040__S _04777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12740_ _00619_ clknet_leaf_24_clock u2.mem\[38\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08509__I _03798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12671_ _00550_ clknet_leaf_156_clock u2.mem\[34\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_276_clock_I clknet_5_23_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11622_ _03486_ _05769_ _05770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09665__I0 _04469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11553_ _05717_ u2.mem\[171\]\[4\] _05721_ _05727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10504_ _05069_ _00896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09417__I0 _04356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11484_ _05668_ u2.mem\[167\]\[1\] _05683_ _05685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13223_ _01102_ clknet_leaf_301_clock u2.mem\[140\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10435_ _04987_ u2.mem\[54\]\[0\] _05030_ _05031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_7_0_clock clknet_0_clock clknet_3_7_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_174_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08180__S _03595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13154_ _01033_ clknet_leaf_281_clock u2.mem\[129\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10366_ _04913_ u2.mem\[52\]\[12\] _04981_ _04982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_48_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12105_ _01488_ clknet_leaf_25_clock u2.active_mem\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10215__S _04887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06946__A4 _02424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13085_ _00964_ clknet_leaf_276_clock u2.mem\[60\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12721__CLK clknet_leaf_248_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10297_ _04920_ u2.mem\[50\]\[15\] _04938_ _04942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12036_ row_select_trans\[5\].A clknet_leaf_303_clock row_select_trans\[5\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06159__A2 _01665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09803__I _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12871__CLK clknet_leaf_134_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10949__I _05345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07659__A2 _03053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12938_ _00817_ clknet_leaf_148_clock u2.mem\[50\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06316__C1 u2.mem\[163\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07323__I _02460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12101__CLK clknet_leaf_246_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12869_ _00748_ clknet_leaf_85_clock u2.mem\[46\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13227__CLK clknet_leaf_300_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09656__I0 _04498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06390_ u2.mem\[175\]\[5\] _01601_ _01631_ u2.mem\[188\]\[5\] _01892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_72_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07292__B1 _02676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08060_ data_in_trans\[7\].data_sync _03514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09408__I0 _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12251__CLK clknet_leaf_228_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13377__CLK clknet_leaf_8_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07831__A2 _03137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07011_ _02489_ _02490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11766__I1 u2.mem\[185\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07595__A1 _03058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08962_ _04019_ u2.mem\[20\]\[2\] _04097_ _04100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07913_ _03374_ _03375_ _03376_ _03377_ _03378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_08893_ _04028_ u2.mem\[18\]\[6\] _04056_ _04059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08395__I0 _03718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07844_ u2.mem\[23\]\[12\] _03148_ _03149_ u2.mem\[22\]\[12\] _03311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06555__C1 u2.mem\[181\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_9_0_clock clknet_4_4_0_clock clknet_5_9_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_68_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07775_ _03239_ _03240_ _03241_ _03242_ _03243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09514_ _04375_ u2.mem\[32\]\[8\] _04453_ _04454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06726_ _02205_ _02206_ _02207_ _02208_ _02209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__08329__I data_in_trans\[10\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09445_ _04412_ _00494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06657_ _02141_ _02142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09376_ _04366_ u2.mem\[29\]\[4\] _04367_ _04368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09647__I0 _04489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_28_0_clock_I clknet_4_14_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06588_ u2.mem\[184\]\[0\] _02072_ _01995_ _02073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10257__I1 u2.mem\[49\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08327_ _03697_ u2.mem\[5\]\[9\] _03693_ _03698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08075__A2 _03518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07283__B1 _02532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08258_ _03645_ _00074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08064__I data_in_trans\[8\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07822__A2 _03282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07209_ u2.mem\[18\]\[1\] _02604_ _02606_ u2.mem\[19\]\[1\] _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_10_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08189_ _03577_ u2.mem\[2\]\[14\] _03600_ _03603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12744__CLK clknet_leaf_43_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10220_ _04575_ _04893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10151_ _04840_ _04851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06794__C1 u2.mem\[159\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09824__S _04649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10082_ _04604_ _04810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12894__CLK clknet_leaf_224_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07338__A1 u2.mem\[58\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08386__I0 _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07338__B2 u2.mem\[36\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12124__CLK clknet_leaf_37_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08138__I0 _03570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10984_ _05346_ u2.mem\[136\]\[3\] _05365_ _05369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09886__I0 _04687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07143__I _02621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12723_ _00602_ clknet_leaf_25_clock u2.mem\[37\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11693__I0 _05794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12654_ _00533_ clknet_leaf_218_clock u2.mem\[33\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06982__I _02460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12274__CLK clknet_leaf_176_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09638__I0 _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11605_ _05759_ _01307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_169_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12585_ _00464_ clknet_leaf_117_clock u2.mem\[28\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08066__A2 _03518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11536_ _05716_ _01281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11467_ _05672_ _01256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13206_ _01085_ clknet_leaf_287_clock u2.mem\[137\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10418_ _05018_ u2.mem\[53\]\[11\] _05012_ _05019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09810__I0 _04576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11398_ _05628_ _01231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13137_ _01016_ clknet_leaf_335_clock u2.mem\[63\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10349_ _04972_ _00838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09734__S _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06222__I _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13068_ _00947_ clknet_leaf_275_clock u2.mem\[59\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_152_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08377__I0 _03684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12019_ net31 clknet_2_3__leaf_clock_a mem_address_trans\[7\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09533__I _04464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08129__I0 _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07560_ _02460_ _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07053__I _02531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12617__CLK clknet_leaf_134_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06511_ _01995_ _01996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07491_ u2.mem\[17\]\[6\] _02846_ _02847_ u2.mem\[24\]\[6\] _02964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07501__A1 _01945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09230_ _04166_ _04278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07501__B2 _02973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06442_ u2.mem\[194\]\[4\] _01924_ _01939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09629__I0 _04471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09161_ _04232_ _00390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11436__I0 _05633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06373_ _01848_ _01853_ _01862_ _01875_ _01876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_124_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08301__I0 _03675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08112_ _03552_ u2.mem\[1\]\[3\] _03546_ _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07265__B1 _02634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09909__S _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09092_ _04181_ _04192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_124_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08043_ data_in_trans\[3\].data_sync _03501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11739__I1 u2.mem\[183\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07017__B1 _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_224_clock_I clknet_5_29_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09994_ _04754_ _00701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08945_ _04073_ _04089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_83_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08368__I0 _03667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06791__A2 _01995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08876_ _04048_ u2.mem\[17\]\[15\] _04042_ _04049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09443__I _04395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input22_I data_in_a[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07827_ u2.mem\[60\]\[12\] _03292_ _03293_ u2.mem\[62\]\[12\] _03294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10589__I _03712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07740__A1 u2.mem\[32\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07758_ u2.mem\[43\]\[11\] _03053_ _03054_ u2.mem\[20\]\[11\] _03226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_72_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06709_ u2.mem\[180\]\[1\] _02043_ _02192_ u2.mem\[150\]\[1\] _02193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__13542__CLK clknet_leaf_18_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07689_ u2.mem\[8\]\[9\] _03093_ _03094_ u2.mem\[4\]\[9\] _03159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08540__I0 _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09428_ _04369_ u2.mem\[30\]\[5\] _04401_ _04403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09359_ _04355_ _00465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09245__A1 _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11213__I _03505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07256__B1 _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11978__I1 u2.mem\[194\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12370_ _00249_ clknet_leaf_158_clock u2.mem\[15\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11321_ _05552_ u2.mem\[157\]\[3\] _05576_ _05580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08522__I _03798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11252_ _05500_ u2.mem\[153\]\[0\] _05537_ _05538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10203_ _04813_ u2.mem\[48\]\[13\] _04880_ _04882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11183_ _05460_ u2.mem\[149\]\[0\] _05492_ _05493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07138__I _02616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06231__A1 u2.mem\[158\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10134_ _04782_ u2.mem\[47\]\[0\] _04841_ _04842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06231__B2 u2.mem\[151\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13072__CLK clknet_leaf_335_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10065_ _04798_ _00728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07731__A1 _03196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06534__A2 _02018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10967_ _05343_ u2.mem\[135\]\[2\] _05356_ _05359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06298__A1 u2.mem\[146\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12706_ _00585_ clknet_leaf_237_clock u2.mem\[36\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07495__B1 _02923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06298__B2 u2.mem\[186\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10898_ _05313_ _01046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07601__I _02576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_173_clock_I clknet_5_26_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12637_ _00516_ clknet_leaf_214_clock u2.mem\[32\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12568_ _00447_ clknet_leaf_135_clock u2.mem\[27\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11519_ _05677_ u2.mem\[169\]\[4\] _05699_ _05705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10962__I _05355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12499_ _00378_ clknet_leaf_119_clock u2.mem\[23\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06470__A1 _01958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08432__I _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06991_ _02469_ _02470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11793__I _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08730_ _03929_ u2.mem\[14\]\[11\] _03951_ _03955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_98_clock_I clknet_5_10_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08661_ _03910_ _00212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13565__CLK clknet_leaf_13_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07722__A1 u2.mem\[26\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07612_ _02600_ _03083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08592_ _03867_ _00186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07543_ _03011_ _03012_ _03013_ _03014_ _03015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_35_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08278__A2 _03544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06289__B2 u2.mem\[194\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07474_ u2.mem\[44\]\[6\] _02889_ _02890_ u2.mem\[42\]\[6\] _02947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_161_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09213_ _04266_ _00408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11409__I0 _05635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06425_ _01545_ _01915_ _01921_ _01925_ _01458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_72_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09144_ _04221_ _00384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07238__B1 _02660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06356_ u2.mem\[159\]\[4\] _01603_ _01594_ u2.mem\[149\]\[4\] _01859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_163_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09075_ _04119_ u2.mem\[22\]\[0\] _04182_ _04183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_159_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06287_ u2.mem\[193\]\[2\] _01731_ _01734_ u2.mem\[177\]\[2\] _01792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08026_ _03479_ _03486_ _03487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08342__I _03658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_375_clock_I clknet_5_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09977_ _04739_ _04745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11409__S _05624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08928_ _04023_ u2.mem\[19\]\[4\] _04079_ _04080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08859_ _03700_ _04037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08761__I0 _03922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_4_6_0_clock clknet_3_3_0_clock clknet_4_6_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12932__CLK clknet_leaf_64_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11870_ _05923_ _01408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10821_ _05264_ _01018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11648__I0 _05758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08513__I0 _03819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11144__S _05462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13540_ _01419_ clknet_leaf_12_clock u2.mem\[192\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10752_ _05222_ u2.mem\[61\]\[12\] _05223_ _05224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_77_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13471_ _01350_ clknet_leaf_309_clock u2.mem\[182\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10683_ _05173_ _05179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_71_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12422_ _00301_ clknet_leaf_101_clock u2.mem\[18\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07229__B1 _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12353_ _00232_ clknet_leaf_160_clock u2.mem\[14\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10782__I _05231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12312__CLK clknet_leaf_117_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11304_ _05570_ _01195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12284_ _00163_ clknet_leaf_199_clock u2.mem\[10\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11235_ _05442_ _05527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_136_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06204__A1 u2.mem\[153\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12462__CLK clknet_leaf_193_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06204__B2 u2.mem\[160\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11166_ _05442_ _05482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_121_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11319__S _05576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06755__A2 _02231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10117_ _04804_ u2.mem\[46\]\[9\] _04830_ _04832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11097_ _05439_ _01119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09083__I _04181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10048_ _04786_ u2.mem\[45\]\[1\] _04784_ _04787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11887__I0 u2.mem\[192\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06507__A2 row_select_trans\[4\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08752__I0 _03913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07180__A2 _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10957__I _05351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11999_ _00011_ clknet_leaf_18_clock u2.mem\[0\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12096__D _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10893__S _05310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06140__B1 _01643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06210_ _01706_ _01711_ _01716_ _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_125_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06691__A1 u2.mem\[166\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06691__B2 u2.mem\[161\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07190_ u2.mem\[61\]\[1\] _02666_ _02667_ u2.mem\[63\]\[1\] _02668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_160_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06141_ _01606_ _01629_ _01638_ _01647_ _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__10692__I _05173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06443__A1 u2.mem\[193\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07640__B1 _03034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06072_ _01551_ _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06443__B2 u2.mem\[192\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12805__CLK clknet_leaf_88_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09900_ _04697_ _00664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10378__I0 _04987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09831_ _04605_ u2.mem\[39\]\[12\] _04654_ _04655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_8_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06746__A2 _02128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08991__I0 _04048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11229__S _05520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12955__CLK clknet_leaf_194_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06974_ u2.mem\[15\]\[0\] _02445_ _02452_ u2.mem\[13\]\[0\] _02453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09762_ _04614_ _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09922__S _04710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08713_ _03945_ _00229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09693_ _04562_ _00592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11878__I0 u2.mem\[192\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08743__I0 _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08644_ _03897_ _00208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08538__S _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07171__A2 _02647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08575_ _03801_ u2.mem\[11\]\[1\] _03856_ _03858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09299__I1 u2.mem\[27\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07459__B1 _02867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07526_ u2.mem\[37\]\[7\] _02829_ _02830_ u2.mem\[59\]\[7\] _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_74_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07457_ _02907_ _02914_ _02921_ _02930_ _02931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_22_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12335__CLK clknet_leaf_159_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06131__C2 u2.mem\[192\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09369__S _04358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06682__A1 u2.mem\[185\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06408_ _01882_ _01887_ _01896_ _01909_ _01910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_07388_ u2.mem\[6\]\[4\] _02694_ _02695_ u2.mem\[47\]\[4\] _02863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_13_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11558__A2 _05729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09127_ _04151_ u2.mem\[23\]\[7\] _04208_ _04212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11802__I0 _05870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06339_ _01809_ _01555_ _01842_ _01483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09168__I _04225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12485__CLK clknet_leaf_109_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09058_ _04169_ _00350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07631__B1 _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06985__A2 _02413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08009_ u2.active_mem\[3\] _03461_ _03462_ u2.active_mem\[2\] _03472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_132_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11020_ _05391_ _01090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_121_clock_I clknet_5_14_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08982__I0 _04039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07416__I _02517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11869__I0 _05913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12971_ _00850_ clknet_leaf_266_clock u2.mem\[53\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10978__S _05365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11922_ _05954_ _01429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08448__S _03777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10541__I0 _05025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07162__A2 _02638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09631__I _04521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13110__CLK clknet_leaf_20_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11853_ _03673_ _05913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10804_ u2.mem\[63\]\[1\] _03496_ _05253_ _05255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08247__I _03633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11784_ _03665_ _05870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_354_clock clknet_5_5_0_clock clknet_leaf_354_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_14_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13523_ _01402_ clknet_leaf_13_clock u2.mem\[190\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06122__B1 _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10735_ _05211_ u2.mem\[61\]\[7\] _05205_ _05212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13260__CLK clknet_leaf_311_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13454_ _01333_ clknet_leaf_320_clock u2.mem\[179\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10666_ _05124_ u2.mem\[59\]\[13\] _05167_ _05169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_167_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12828__CLK clknet_leaf_203_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12405_ _00284_ clknet_leaf_103_clock u2.mem\[17\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10218__S _04887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_369_clock clknet_5_1_0_clock clknet_leaf_369_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13385_ _01264_ clknet_leaf_323_clock u2.mem\[167\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10597_ _05129_ _00929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06425__A1 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07100__B _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12336_ _00215_ clknet_leaf_159_clock u2.mem\[13\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08911__S _04066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12267_ _00146_ clknet_leaf_194_clock u2.mem\[9\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12978__CLK clknet_leaf_265_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11218_ _05516_ _05517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12198_ _00077_ clknet_leaf_22_clock u2.mem\[4\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07925__A1 u2.mem\[14\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11049__S _05403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08973__I0 _04030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11149_ _05351_ _05472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12208__CLK clknet_leaf_241_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10780__I0 _05211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07326__I _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09742__S _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_307_clock clknet_5_20_0_clock clknet_leaf_307_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_37_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06690_ _02108_ _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10532__I0 _05016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07153__A2 _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_323_clock_I clknet_5_16_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12358__CLK clknet_leaf_92_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06361__B1 _01710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08360_ _03542_ _03724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08157__I _03584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07311_ _02384_ _02786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08291_ _03668_ _00084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10835__I1 _05229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07456__A3 _02926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06113__B1 _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07996__I _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07242_ _02703_ _02708_ _02713_ _02718_ _02719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__06664__A1 u2.mem\[170\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06664__B2 u2.mem\[156\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07173_ _02500_ _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10128__S _04835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06124_ _01581_ _01630_ _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07613__B1 _03083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06055_ col_select_trans\[0\].data_sync _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09716__I _04566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08620__I _03878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07916__A1 u2.mem\[16\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08964__I0 _04021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09814_ _04645_ _00630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10771__I0 _05202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06195__A3 _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13133__CLK clknet_leaf_282_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09745_ _04601_ _04602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10798__S _05247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06957_ _02435_ _02436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09676_ _04480_ u2.mem\[36\]\[7\] _04549_ _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06888_ _02353_ _02367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10523__I0 _05007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07144__A2 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08627_ _03814_ u2.mem\[12\]\[7\] _03884_ _03888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13283__CLK clknet_leaf_384_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08558_ _03821_ u2.mem\[10\]\[10\] _03845_ _03848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09141__I0 _04171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07509_ u2.mem\[16\]\[7\] _02800_ _02801_ u2.mem\[33\]\[7\] _02981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_11_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10826__I1 _03524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08489_ _03666_ _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09692__I1 u2.mem\[36\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09099__S _04192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06655__A1 u2.mem\[154\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10520_ _05079_ _00902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06655__B2 u2.mem\[162\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10451_ _05039_ _00873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10038__S _04777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09444__I1 u2.mem\[30\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06407__A1 _01901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13170_ _01049_ clknet_leaf_283_clock u2.mem\[131\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10382_ _04992_ u2.mem\[53\]\[1\] _04989_ _04993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06958__A2 _02432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12121_ _01484_ clknet_leaf_348_clock u2.select_mem_col\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_174_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_272_clock_I clknet_5_23_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12052_ data_in_trans\[1\].A clknet_leaf_378_clock data_in_trans\[1\].data_sync vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07907__A1 _03357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11003_ _05379_ _01085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06186__A3 _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11891__I _05928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10501__S _05066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08178__S _03595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12954_ _00833_ clknet_leaf_146_clock u2.mem\[51\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10514__I0 _04995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11905_ u2.mem\[192\]\[12\] _03527_ _05942_ _05945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_3_3_0_clock clknet_0_clock clknet_3_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12885_ _00764_ clknet_leaf_75_clock u2.mem\[47\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06343__B1 _01658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_293_clock clknet_5_21_0_clock clknet_leaf_293_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10300__I _04943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11836_ _05901_ _01396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09132__I0 _04158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12650__CLK clknet_leaf_114_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10817__I1 _03514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11767_ _05859_ _01369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13506_ _01385_ clknet_leaf_333_clock u2.mem\[187\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08705__I _03940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10718_ _04994_ _05200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11698_ _05816_ _01343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13437_ _01316_ clknet_leaf_366_clock u2.mem\[176\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13006__CLK clknet_leaf_270_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10649_ _05159_ _00951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09435__I1 u2.mem\[30\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11242__I1 u2.mem\[152\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06225__I _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08641__S _03894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13368_ _01247_ clknet_leaf_372_clock u2.mem\[164\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_231_clock clknet_5_28_0_clock clknet_leaf_231_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06949__A2 _02415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12319_ _00198_ clknet_leaf_161_clock u2.mem\[12\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13299_ _01178_ clknet_leaf_382_clock u2.mem\[153\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09199__I0 _04256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09536__I _04127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12030__CLK clknet_leaf_303_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13156__CLK clknet_leaf_283_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08946__I0 _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07860_ _02611_ _03327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_246_clock clknet_5_18_0_clock clknet_leaf_246_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_64_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08571__A1 _03480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06811_ u2.mem\[170\]\[4\] _02146_ _02148_ u2.mem\[156\]\[4\] _02292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_42_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07791_ u2.mem\[27\]\[12\] _03104_ _03105_ u2.mem\[35\]\[12\] _03258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11507__S _05691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09530_ _04462_ _00529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06742_ _02126_ _02225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_49_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06895__I _02373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10505__I0 _05027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09461_ _04422_ _00500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06673_ _02157_ _02158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08412_ _03671_ u2.mem\[7\]\[3\] _03753_ _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_169_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09392_ _04378_ u2.mem\[29\]\[9\] _04376_ _04379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_24_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09123__I0 _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08343_ _03709_ u2.mem\[5\]\[12\] _03710_ _03711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10808__I1 _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11242__S _05529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08274_ _03490_ _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07225_ u2.mem\[27\]\[2\] _02638_ _02639_ u2.mem\[35\]\[2\] _02702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_5_0_clock clknet_4_2_0_clock clknet_5_5_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__09426__I1 u2.mem\[30\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09647__S _04532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07156_ _02435_ _02634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08551__S _03840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11233__I1 u2.mem\[151\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06107_ _01593_ _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07062__A1 _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07087_ _02522_ _02523_ _02485_ _02408_ _02566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_161_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10992__I0 _05335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06038_ _01544_ _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08350__I data_in_trans\[14\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08937__I0 _04032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12523__CLK clknet_leaf_187_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07989_ u2.mem\[39\]\[15\] _03323_ _03324_ u2.mem\[48\]\[15\] _03453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11417__S _05638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09728_ _04588_ _04589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10321__S _04954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09659_ _04095_ _04542_ _04543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06876__A1 _02339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12670_ _00549_ clknet_leaf_217_clock u2.mem\[34\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08726__S _03951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_219_clock_I clknet_5_29_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09114__I0 _04128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11621_ _05768_ _05769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13029__CLK clknet_leaf_29_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08525__I _03713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11552_ _05726_ _01287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10503_ _05025_ u2.mem\[55\]\[14\] _05066_ _05069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11483_ _05684_ _01260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09417__I1 u2.mem\[30\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12053__CLK clknet_2_0__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13222_ _01101_ clknet_leaf_300_clock u2.mem\[140\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13179__CLK clknet_leaf_279_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10434_ _05029_ _05030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08461__S _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10365_ _04965_ _04981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_152_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13153_ _01032_ clknet_leaf_283_clock u2.mem\[129\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12104_ _01487_ clknet_leaf_25_clock u2.active_mem\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13084_ _00963_ clknet_leaf_277_clock u2.mem\[60\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10296_ _04941_ _00816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08928__I0 _04023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12035_ net42 clknet_2_3__leaf_clock_a row_select_trans\[5\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08002__B1 _03462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10735__I0 _05211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09292__S _04313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06159__A3 _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_2_0_clock_I clknet_4_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10231__S _04896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07604__I _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12937_ _00816_ clknet_leaf_148_clock u2.mem\[50\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11160__I0 _05468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06316__C2 _01643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06867__A1 _02338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08636__S _03889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12868_ _00747_ clknet_leaf_85_clock u2.mem\[46\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11819_ _05872_ u2.mem\[188\]\[3\] _05888_ _05892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12799_ _00678_ clknet_leaf_167_clock u2.mem\[42\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11062__S _05413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07010_ _02455_ _02479_ _02481_ _02488_ _02489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_31_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_170_clock clknet_5_26_0_clock clknet_leaf_170_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_127_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11215__I1 u2.mem\[150\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12546__CLK clknet_leaf_189_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08961_ _04099_ _00323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08919__I0 _04010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_185_clock clknet_5_30_0_clock clknet_leaf_185_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07912_ u2.mem\[27\]\[14\] _02420_ _02426_ u2.mem\[35\]\[14\] _03377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08892_ _04058_ _00295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10726__I0 _05204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_168_clock_I clknet_5_26_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12696__CLK clknet_leaf_140_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09592__I0 _04471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07843_ _03300_ _03303_ _03306_ _03309_ _03310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07774_ u2.mem\[18\]\[11\] _03085_ _03086_ u2.mem\[19\]\[11\] _03242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_42_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09513_ _04442_ _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06725_ u2.mem\[184\]\[2\] _02072_ _01994_ _02208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_25_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06858__A1 _01878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09444_ _04384_ u2.mem\[30\]\[12\] _04411_ _04412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06656_ _02064_ _02119_ _02141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_220_clock_I clknet_5_29_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_123_clock clknet_5_15_0_clock clknet_leaf_123_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09375_ _04357_ _04367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06587_ _02071_ _02072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12076__CLK clknet_leaf_39_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08326_ _03696_ _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08345__I data_in_trans\[13\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_28_0_clock clknet_4_14_0_clock clknet_5_28_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_71_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13321__CLK clknet_leaf_321_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06293__C _01797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07283__A1 u2.mem\[49\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08257_ _03563_ u2.mem\[4\]\[8\] _03644_ _03645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_138_clock clknet_5_14_0_clock clknet_leaf_138_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_20_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07208_ u2.mem\[52\]\[1\] _02599_ _02601_ u2.mem\[21\]\[1\] _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_140_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08188_ _03602_ _00047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07139_ _02506_ _02614_ _02615_ _02383_ _02618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10316__S _04949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13471__CLK clknet_leaf_309_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10965__I0 _05340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07586__A2 _03038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10150_ _04850_ _00761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06794__B1 _02098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06794__C2 _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10081_ _04809_ _00733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09904__I _04591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08386__I1 u2.mem\[6\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11147__S _05461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10051__S _04784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10986__S _05364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10983_ _05368_ _01076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12722_ _00601_ clknet_leaf_249_clock u2.mem\[37\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06849__B2 u2.mem\[162\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12419__CLK clknet_leaf_104_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11693__I1 u2.mem\[180\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12653_ _00532_ clknet_leaf_218_clock u2.mem\[33\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11604_ _05758_ u2.mem\[174\]\[5\] _05747_ _05759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_168_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12584_ _00463_ clknet_leaf_110_clock u2.mem\[28\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12569__CLK clknet_leaf_128_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11535_ _05715_ u2.mem\[170\]\[3\] _05709_ _05716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_8_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11610__S _05761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08191__S _03600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11466_ _05671_ u2.mem\[166\]\[2\] _05665_ _05672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_172_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13205_ _01084_ clknet_leaf_292_clock u2.mem\[137\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10417_ _03703_ _05018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11397_ _05627_ u2.mem\[162\]\[1\] _05625_ _05628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07577__A2 _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06503__I row_select_trans\[2\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13136_ _01015_ clknet_leaf_330_clock u2.mem\[63\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10348_ _04895_ u2.mem\[52\]\[4\] _04971_ _04972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10279_ _04902_ u2.mem\[50\]\[7\] _04928_ _04932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13067_ _00946_ clknet_leaf_263_clock u2.mem\[59\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_152_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10708__I0 _05128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12018_ mem_address_trans\[6\].A clknet_leaf_315_clock mem_address_trans\[6\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11381__I0 _05587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07334__I _02482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_40_clock clknet_5_6_0_clock clknet_leaf_40_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06510_ _01994_ _01995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12099__CLK clknet_leaf_247_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07490_ u2.mem\[23\]\[6\] _02915_ _02916_ u2.mem\[22\]\[6\] _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_34_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08366__S _03727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13344__CLK clknet_leaf_6_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06441_ _01914_ _01938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09160_ _04140_ u2.mem\[24\]\[4\] _04231_ _04232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_128_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_55_clock clknet_5_12_0_clock clknet_leaf_55_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06372_ _01867_ _01868_ _01869_ _01874_ _01875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__11436__I1 u2.mem\[164\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08111_ _03502_ _03552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_147_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09091_ _04191_ _00361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_94_clock_I clknet_5_10_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07265__B2 u2.mem\[34\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13494__CLK clknet_leaf_309_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08042_ _01773_ _03489_ _03500_ _00003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_159_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07017__A1 u2.mem\[50\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07017__B2 u2.mem\[51\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10136__S _04841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07568__A2 _02880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09925__S _04710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06413__I _01913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09993_ _04707_ u2.mem\[43\]\[11\] _04750_ _04754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06776__B1 _02078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08944_ _04088_ _00317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08875_ _03721_ _04048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07826_ _02543_ _03293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09317__I0 _04283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input15_I data_in_a[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07740__A2 _03019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07757_ u2.mem\[49\]\[11\] _03050_ _03051_ u2.mem\[46\]\[11\] _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_44_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06708_ _02047_ _02192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_371_clock_I clknet_5_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07688_ u2.mem\[39\]\[9\] _03090_ _03091_ u2.mem\[48\]\[9\] _03158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_13_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09427_ _04402_ _00486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06639_ u2.mem\[185\]\[0\] _02121_ _02123_ u2.mem\[173\]\[0\] _02124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_157_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09358_ _04285_ u2.mem\[28\]\[15\] _04351_ _04355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08309_ _03682_ _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09289_ _04315_ _00435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11430__S _05647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11320_ _05579_ _01202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_4_2_0_clock clknet_3_1_0_clock clknet_4_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_165_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12861__CLK clknet_leaf_203_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11251_ _05536_ _05537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10938__I0 _05335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10202_ _04881_ _00782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09835__S _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11182_ _05491_ _05492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_171_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10133_ _04840_ _04841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__13217__CLK clknet_leaf_295_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09556__I0 _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10064_ _04797_ u2.mem\[45\]\[6\] _04793_ _04798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_121_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07192__B1 _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09308__I0 _04274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13367__CLK clknet_leaf_371_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10966_ _05358_ _01069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12705_ _00584_ clknet_leaf_242_clock u2.mem\[36\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12391__CLK clknet_leaf_140_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10897_ _05301_ u2.mem\[131\]\[2\] _05310_ _05313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_116_clock_I clknet_5_14_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12636_ _00515_ clknet_leaf_215_clock u2.mem\[32\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08295__I0 _03671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12567_ _00446_ clknet_leaf_116_clock u2.mem\[27\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_10_0_clock_I clknet_4_5_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11518_ _05704_ _01275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12498_ _00377_ clknet_leaf_175_clock u2.mem\[23\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06470__A2 _01955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11449_ _05659_ _01251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_160_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13119_ _00998_ clknet_leaf_257_clock u2.mem\[62\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06990_ _02387_ _02389_ _02424_ _02459_ _02469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09547__I0 _04473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input7_I data_in_a[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08660_ _03909_ u2.mem\[13\]\[2\] _03905_ _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07183__B1 _02660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07722__A2 _03141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09480__S _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07611_ _02598_ _03082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08591_ _03816_ u2.mem\[11\]\[8\] _03866_ _03867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11106__I0 _05420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07999__I _01665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12734__CLK clknet_leaf_270_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11515__S _05700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07542_ u2.mem\[6\]\[7\] _02927_ _02928_ u2.mem\[47\]\[7\] _03014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_35_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08278__A3 _03632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07473_ _02942_ _02943_ _02944_ _02945_ _02946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_74_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11314__I _05575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09212_ _04265_ u2.mem\[25\]\[6\] _04261_ _04266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11409__I1 u2.mem\[162\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06424_ u2.mem\[194\]\[0\] _01924_ _01925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09143_ _04174_ u2.mem\[23\]\[14\] _04218_ _04221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06355_ u2.mem\[175\]\[4\] _01601_ _01631_ u2.mem\[188\]\[4\] _01858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07238__B2 u2.mem\[12\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10093__I0 _04817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09719__I _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09074_ _04181_ _04182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_148_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06286_ u2.mem\[158\]\[2\] _01565_ _01572_ u2.mem\[151\]\[2\] _01589_ u2.mem\[168\]\[2\]
+ _01791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_147_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_163_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12114__CLK clknet_leaf_349_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08025_ _03485_ _03486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_162_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_318_clock_I clknet_5_17_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06143__I _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09976_ _04744_ _00693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12264__CLK clknet_leaf_55_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08927_ _04073_ _04079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_162_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11345__I0 _05595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08210__I0 _03559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08858_ _04036_ _00283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11896__I1 _03517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07174__B1 _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07713__A2 _03050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07809_ u2.mem\[53\]\[12\] _03274_ _03275_ u2.mem\[56\]\[12\] _03276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_84_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08789_ _03907_ u2.mem\[16\]\[1\] _03990_ _03992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10820_ u2.mem\[63\]\[8\] _03517_ _05263_ _05264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07477__B2 u2.mem\[20\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10751_ _05195_ _05223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13470_ _01349_ clknet_leaf_360_clock u2.mem\[181\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10682_ _05178_ _00965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12421_ _00300_ clknet_leaf_102_clock u2.mem\[18\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07229__B2 u2.mem\[33\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11160__S _05475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10084__I0 _04810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12352_ _00231_ clknet_leaf_161_clock u2.mem\[14\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_166_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11303_ _05548_ u2.mem\[156\]\[1\] _05568_ _05570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_4_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06452__A2 _01946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12283_ _00162_ clknet_leaf_188_clock u2.mem\[10\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12607__CLK clknet_leaf_159_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11234_ _05526_ _01169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11584__I0 _05719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06204__A2 _01708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06988__I _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11165_ _05481_ _01145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09529__I0 _04391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07952__A2 _02432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10116_ _04831_ _00746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_42_clock_I clknet_5_6_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11096_ _05428_ u2.mem\[143\]\[3\] _05435_ _05439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11336__I0 _05589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10047_ _04569_ _04786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08201__I0 _03550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12757__CLK clknet_leaf_71_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08909__S _04066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07165__B1 _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11887__I1 _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07704__A2 _03036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07612__I _02600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11998_ _00010_ clknet_5_3_0_clock u2.mem\[0\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07468__A1 _02937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10949_ _05345_ _05346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11134__I _05461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_267_clock_I clknet_5_22_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06228__I _01583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06140__A1 u2.mem\[145\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06140__B2 u2.mem\[163\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12619_ _00498_ clknet_leaf_206_clock u2.mem\[31\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08268__I0 _03575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12137__CLK clknet_leaf_38_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06691__A2 _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09539__I _04131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06140_ u2.mem\[145\]\[0\] _01640_ _01643_ u2.mem\[163\]\[0\] u2.mem\[165\]\[0\]
+ _01646_ _01647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_34_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08443__I _03774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06071_ u2.mem\[158\]\[0\] _01565_ _01572_ u2.mem\[151\]\[0\] _01577_ u2.mem\[193\]\[0\]
+ _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_145_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07640__B2 u2.mem\[33\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12287__CLK clknet_leaf_178_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13532__CLK clknet_leaf_349_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09830_ _04638_ _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_141_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06898__I _02376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09761_ data_in_trans\[15\].data_sync _04614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06973_ _02451_ _02452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08712_ _03911_ u2.mem\[14\]\[3\] _03941_ _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09692_ _04496_ u2.mem\[36\]\[14\] _04559_ _04562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11878__I1 _03491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08643_ _03830_ u2.mem\[12\]\[14\] _03894_ _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08574_ _03857_ _00178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_78_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07525_ u2.mem\[60\]\[7\] _02826_ _02827_ u2.mem\[62\]\[7\] _02997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_35_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08554__S _03845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07456_ _02924_ _02925_ _02926_ _02929_ _02930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06131__A1 u2.mem\[188\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06131__B2 u2.mem\[187\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08259__I0 _03566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06407_ _01901_ _01902_ _01903_ _01908_ _01909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__13062__CLK clknet_leaf_30_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07387_ u2.mem\[8\]\[4\] _02860_ _02861_ u2.mem\[4\]\[4\] _02862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_41_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09126_ _04211_ _00376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06338_ _01814_ _01819_ _01828_ _01841_ _01842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_159_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11802__I1 u2.mem\[187\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07226__A4 _02702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09057_ _04167_ u2.mem\[21\]\[12\] _04168_ _04169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_159_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06269_ _01615_ _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08008_ _03469_ _03470_ _03471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09759__I0 _04612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11566__I0 _05715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09959_ _04709_ u2.mem\[42\]\[12\] _04734_ _04735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_4102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10123__I _04819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12970_ _00849_ clknet_leaf_127_clock u2.mem\[52\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11869__I1 u2.mem\[191\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07698__A1 u2.mem\[40\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11921_ _05911_ u2.mem\[193\]\[3\] _05950_ _05954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_4179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07698__B2 u2.mem\[30\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06757__B _02239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08528__I _03717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11852_ _05912_ _01401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10803_ _05254_ _01010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10994__S _05373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11783_ _05869_ _01375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13405__CLK clknet_leaf_320_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13522_ _01401_ clknet_leaf_4_clock u2.mem\[190\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06048__I _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10734_ _03686_ _05211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06122__A1 u2.mem\[171\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06122__B2 u2.mem\[157\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13453_ _01332_ clknet_leaf_320_clock u2.mem\[179\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10665_ _05168_ _00958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12404_ _00283_ clknet_leaf_103_clock u2.mem\[17\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09998__I0 _04712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13384_ _01263_ clknet_leaf_318_clock u2.mem\[167\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10596_ _05128_ u2.mem\[57\]\[15\] _05122_ _05129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12335_ _00214_ clknet_leaf_159_clock u2.mem\[13\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06425__A2 _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08670__I0 _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07100__C _02408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09295__S _04318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12266_ _00145_ clknet_leaf_54_clock u2.mem\[8\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11217_ _03509_ _05516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10234__S _04896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06189__A1 _01685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12197_ _00076_ clknet_leaf_23_clock u2.mem\[4\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07925__A2 _02521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08973__I1 u2.mem\[20\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06511__I _01995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11148_ _05471_ _01138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11309__I0 _05554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10033__I _04761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08639__S _03894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11079_ _05345_ _05428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09922__I0 _04712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07153__A3 _02608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07342__I _02527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13085__CLK clknet_leaf_276_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07310_ u2.mem\[45\]\[4\] _02633_ _02634_ u2.mem\[34\]\[4\] _02785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_36_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08290_ _03667_ u2.mem\[5\]\[2\] _03659_ _03668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06113__A1 u2.mem\[178\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07310__B1 _02634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06113__B2 u2.mem\[164\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07241_ _02714_ _02715_ _02716_ _02717_ _02718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_108_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10409__S _05012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06664__A2 _02146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10048__I0 _04786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09989__I0 _04703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07172_ _02498_ _02650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_157_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06123_ _01558_ _01559_ _01585_ _01630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_145_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06054_ _01560_ _01561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09813_ _04579_ u2.mem\[39\]\[4\] _04644_ _04645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06421__I _01911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10920__A1 _04121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09744_ data_in_trans\[11\].data_sync _04601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06956_ _02421_ _02433_ _02434_ _02393_ _02435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_100_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08549__S _03840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09732__I _04591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_1_0_clock clknet_4_0_0_clock clknet_5_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_09675_ _04552_ _00584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06887_ _02339_ _02338_ _02344_ _02366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07144__A3 _02615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13428__CLK clknet_leaf_352_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08626_ _03887_ _00200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06352__A1 u2.mem\[158\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06352__B2 u2.mem\[151\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08557_ _03847_ _00171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11703__S _05818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07508_ u2.mem\[1\]\[7\] _02797_ _02798_ u2.mem\[7\]\[7\] _02980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_165_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08488_ _03802_ _00147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12452__CLK clknet_leaf_90_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07447__A4 _02920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13578__CLK clknet_leaf_35_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07439_ u2.mem\[28\]\[5\] _02841_ _02842_ u2.mem\[31\]\[5\] _02913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_10_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06655__A2 _02126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10319__S _04954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10450_ _05009_ u2.mem\[54\]\[7\] _05035_ _05039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_109_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09109_ _04201_ _00369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06407__A2 _01902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10381_ _04991_ _04992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12120_ _01483_ clknet_leaf_348_clock u2.select_mem_col\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_215_clock_I clknet_5_29_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10054__S _04784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12051_ net14 clknet_2_1__leaf_clock_a data_in_trans\[1\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07907__A2 _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_4_2_0_clock_I clknet_3_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11002_ _05352_ u2.mem\[137\]\[5\] _05372_ _05379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08459__S _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12953_ _00832_ clknet_leaf_148_clock u2.mem\[51\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11711__I0 _05798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11904_ _05944_ _01421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12884_ _00763_ clknet_leaf_75_clock u2.mem\[47\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06343__B2 u2.mem\[155\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11835_ _05874_ u2.mem\[189\]\[4\] _05895_ _05901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08096__A1 _03478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11766_ _05829_ u2.mem\[185\]\[1\] _05857_ _05859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13505_ _01384_ clknet_leaf_333_clock u2.mem\[187\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10717_ _05199_ _00979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08891__I0 _04026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11412__I _05637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11697_ _05798_ u2.mem\[180\]\[5\] _05809_ _05816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12945__CLK clknet_leaf_151_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07111__B _02401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13436_ _01315_ clknet_leaf_353_clock u2.mem\[176\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10648_ _05106_ u2.mem\[59\]\[5\] _05157_ _05159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08643__I0 _03830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13367_ _01246_ clknet_leaf_371_clock u2.mem\[164\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10579_ _03699_ _05117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10450__I0 _05009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12318_ _00197_ clknet_leaf_185_clock u2.mem\[12\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06803__C1 u2.mem\[145\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13298_ _01177_ clknet_leaf_382_clock u2.mem\[153\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09199__I1 u2.mem\[25\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12249_ _00128_ clknet_leaf_55_clock u2.mem\[7\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07359__B1 _02676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07337__I _02489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06241__I _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10899__S _05310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06810_ u2.mem\[146\]\[4\] _02156_ _02158_ u2.mem\[186\]\[4\] _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_95_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07790_ u2.mem\[40\]\[12\] _03255_ _03256_ u2.mem\[30\]\[12\] _03257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09552__I _04147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06741_ u2.mem\[144\]\[2\] _02115_ _02117_ u2.mem\[182\]\[2\] _02224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_36_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09460_ _04362_ u2.mem\[31\]\[2\] _04419_ _04422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06672_ _02125_ _02014_ _02157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06334__A1 u2.mem\[146\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06334__B2 u2.mem\[186\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08411_ _03756_ _00116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09391_ _04157_ _04378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06885__A2 _01997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09123__I1 u2.mem\[23\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08342_ _03658_ _03710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08087__A1 _01976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07800__I _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_164_clock_I clknet_5_26_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08273_ _03653_ _00081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06637__A2 _02018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08882__I0 _04017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07224_ u2.mem\[40\]\[2\] _02403_ _02410_ u2.mem\[30\]\[2\] _02701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09928__S _04710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08634__I0 _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07155_ _02431_ _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09727__I data_in_trans\[7\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06106_ _01561_ _01613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_161_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07086_ u2.mem\[29\]\[0\] _02559_ _02564_ u2.mem\[11\]\[0\] _02565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13100__CLK clknet_leaf_281_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06270__B1 _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06037_ u2.mem\[0\]\[0\] _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_160_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09663__S _04544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_353_clock clknet_5_5_0_clock clknet_leaf_353_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08011__A1 _03472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_5_24_0_clock clknet_4_12_0_clock clknet_5_24_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13250__CLK clknet_leaf_295_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10602__S _05131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07988_ u2.mem\[5\]\[15\] _02627_ _02629_ u2.mem\[38\]\[15\] _03452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06573__A1 _02056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_89_clock_I clknet_5_11_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09727_ data_in_trans\[7\].data_sync _04588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06939_ _02407_ _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_41_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_368_clock clknet_5_1_0_clock clknet_leaf_368_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_16_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10401__I _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09658_ _04440_ _04542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08078__I data_in_trans\[12\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06325__A1 u2.mem\[144\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06325__B2 u2.mem\[182\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08609_ _03876_ _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06876__A2 _02354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09589_ _04503_ _00547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12968__CLK clknet_leaf_128_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11620_ _04861_ _05274_ _05768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_70_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11551_ _05715_ u2.mem\[171\]\[3\] _05722_ _05726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06628__A2 _02090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08873__I0 _04046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10502_ _05068_ _00895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11482_ _05663_ u2.mem\[167\]\[0\] _05683_ _05684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_306_clock clknet_5_20_0_clock clknet_leaf_306_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13221_ _01100_ clknet_leaf_300_clock u2.mem\[140\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08625__I0 _03812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10433_ _04180_ _04964_ _05029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13152_ _01031_ clknet_leaf_260_clock u2.mem\[128\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10364_ _04980_ _00845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12348__CLK clknet_leaf_207_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12103_ _01501_ clknet_leaf_29_clock u2.active_mem\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_366_clock_I clknet_5_4_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06261__B1 _01710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06261__C2 u2.mem\[194\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13083_ _00962_ clknet_leaf_261_clock u2.mem\[60\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10295_ _04918_ u2.mem\[50\]\[14\] _04938_ _04941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08002__A1 u2.active_mem\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12034_ row_select_trans\[4\].A clknet_leaf_301_clock row_select_trans\[4\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06061__I col_select_trans\[3\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08002__B2 u2.active_mem\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10735__I1 u2.mem\[61\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11608__S _05761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10512__S _05073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08189__S _03600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12498__CLK clknet_leaf_175_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07761__B1 _03133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_6_0_clock_I clknet_4_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10499__I0 _05020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07106__B _02454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12936_ _00815_ clknet_leaf_147_clock u2.mem\[50\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06316__A1 u2.mem\[177\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07513__B1 _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06316__B2 u2.mem\[165\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11160__I1 u2.mem\[147\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12867_ _00746_ clknet_leaf_86_clock u2.mem\[46\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11818_ _05891_ _01388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08069__A1 _03520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12798_ _00677_ clknet_leaf_208_clock u2.mem\[42\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07620__I _02618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11749_ _05848_ _05849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_144_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07292__A2 _02675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13123__CLK clknet_leaf_21_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_146_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13419_ _01298_ clknet_leaf_318_clock u2.mem\[173\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08616__I0 _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08960_ _04017_ u2.mem\[20\]\[1\] _04097_ _04099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13273__CLK clknet_leaf_7_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07911_ u2.mem\[40\]\[14\] _03255_ _03256_ u2.mem\[30\]\[14\] _03376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08891_ _04026_ u2.mem\[18\]\[5\] _04056_ _04058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10726__I1 u2.mem\[61\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07842_ u2.mem\[28\]\[12\] _03307_ _03308_ u2.mem\[31\]\[12\] _03309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09592__I1 u2.mem\[34\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10422__S _05021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_90_clock_I clknet_5_10_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06555__A1 u2.mem\[155\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07752__B1 _03042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06839__C _02318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07773_ u2.mem\[52\]\[11\] _03082_ _03083_ u2.mem\[21\]\[11\] _03241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09512_ _04452_ _00521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06724_ u2.mem\[171\]\[2\] _02066_ _02068_ u2.mem\[157\]\[2\] _02207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_77_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06307__A1 u2.mem\[167\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06307__B2 u2.mem\[183\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09443_ _04395_ _04411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_25_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06655_ u2.mem\[154\]\[0\] _02126_ _02127_ u2.mem\[162\]\[0\] _02139_ _02140_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_24_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09374_ _04139_ _04366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06586_ _02060_ _02070_ _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08325_ _03695_ _03696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07283__A2 _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08256_ _03633_ _03644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07207_ u2.mem\[17\]\[1\] _02586_ _02591_ u2.mem\[24\]\[1\] _02685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06491__B1 _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08187_ _03575_ u2.mem\[2\]\[13\] _03600_ _03602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07138_ _02616_ _02617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08232__A1 mem_address_trans\[1\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09280__I0 _04285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07586__A3 _03047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_292_clock clknet_5_21_0_clock clknet_leaf_292_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07069_ _02547_ _02548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06794__A1 u2.mem\[166\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07991__B1 _02624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06794__B2 u2.mem\[161\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12640__CLK clknet_leaf_157_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10080_ _04808_ u2.mem\[45\]\[11\] _04802_ _04809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11428__S _05647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10332__S _04959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09192__I _04251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12790__CLK clknet_leaf_33_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10982_ _05343_ u2.mem\[136\]\[2\] _05365_ _05368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12721_ _00600_ clknet_leaf_248_clock u2.mem\[37\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_230_clock clknet_5_28_0_clock clknet_leaf_230_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_55_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09099__I0 _04164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12652_ _00531_ clknet_leaf_218_clock u2.mem\[33\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12020__CLK clknet_leaf_315_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13146__CLK clknet_leaf_40_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11603_ _05679_ _05758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12583_ _00462_ clknet_leaf_112_clock u2.mem\[28\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_245_clock clknet_5_24_0_clock clknet_leaf_245_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_8_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11534_ _05673_ _05715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07274__A2 _02470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12170__CLK clknet_leaf_59_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11465_ _05670_ _05671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13296__CLK clknet_leaf_370_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10405__I0 _05009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13204_ _01083_ clknet_leaf_293_clock u2.mem\[137\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10416_ _05017_ _00860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09271__I0 _04276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11396_ _05504_ _05627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13135_ _01014_ clknet_leaf_330_clock u2.mem\[63\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10347_ _04965_ _04971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_140_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06785__A1 u2.mem\[179\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06785__B2 u2.mem\[191\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_112_clock_I clknet_5_11_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13066_ _00945_ clknet_leaf_339_clock u2.mem\[58\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10278_ _04931_ _00808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10708__I1 u2.mem\[60\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12017_ net30 clknet_2_3__leaf_clock_a mem_address_trans\[6\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07615__I _02605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11381__I1 u2.mem\[161\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11137__I _05339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09830__I _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12919_ _00798_ clknet_leaf_134_clock u2.mem\[49\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06440_ _01809_ _01915_ _01936_ _01937_ _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_62_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08837__I0 _04021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06371_ u2.mem\[147\]\[4\] _01675_ _01679_ u2.mem\[169\]\[4\] _01873_ _01874_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__12513__CLK clknet_leaf_175_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09478__S _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08110_ _03551_ _00020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_37_clock_I clknet_5_6_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09090_ _04151_ u2.mem\[22\]\[7\] _04187_ _04191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07265__A2 _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08382__S _03737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08041_ _03499_ _03493_ _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_163_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07017__A2 _02493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09262__I0 _04267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09992_ _04753_ _00700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06776__A1 u2.mem\[165\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06776__B2 u2.mem\[163\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07973__B1 _02555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08943_ _04039_ u2.mem\[19\]\[11\] _04084_ _04088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13019__CLK clknet_leaf_266_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11248__S _05528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10152__S _04851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08874_ _04047_ _00288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07725__B1 _03075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09941__S _04724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07825_ _02541_ _03292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09317__I1 u2.mem\[27\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07756_ u2.mem\[14\]\[11\] _03125_ _03126_ u2.mem\[12\]\[11\] _03224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12043__CLK clknet_2_2__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09740__I data_in_trans\[10\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11124__I1 u2.mem\[145\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13169__CLK clknet_leaf_283_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_314_clock_I clknet_5_17_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06707_ u2.mem\[155\]\[1\] _02030_ _02035_ u2.mem\[174\]\[1\] u2.mem\[181\]\[1\]
+ _02039_ _02191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_07687_ u2.mem\[5\]\[9\] _03155_ _03156_ u2.mem\[38\]\[9\] _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_25_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09426_ _04366_ u2.mem\[30\]\[4\] _04401_ _04402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10883__I0 _05303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08356__I _03720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06638_ _02122_ _02123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06700__A1 u2.mem\[171\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06700__B2 u2.mem\[157\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08828__I0 _04010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09357_ _04354_ _00464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12193__CLK clknet_leaf_253_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06569_ _02053_ _02054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11711__S _05817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08308_ data_in_trans\[6\].data_sync _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07256__A2 _02604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09288_ _04254_ u2.mem\[27\]\[1\] _04313_ _04315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06464__B1 _01943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08239_ _03538_ u2.mem\[4\]\[0\] _03634_ _03635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_5_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11250_ _04248_ _05527_ _05536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__06604__I _02088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09253__I0 _04258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10201_ _04810_ u2.mem\[48\]\[12\] _04880_ _04881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11060__I0 _05386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11181_ _04120_ _05482_ _05491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06767__B2 u2.mem\[152\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10132_ _04417_ _04760_ _04840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11158__S _05475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10063_ _04585_ _04797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07435__I _02568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09308__I1 u2.mem\[27\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10965_ _05340_ u2.mem\[135\]\[1\] _05356_ _05358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12536__CLK clknet_leaf_109_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12704_ _00583_ clknet_leaf_238_clock u2.mem\[36\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10874__I0 _05294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07495__A2 _02922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10896_ _05312_ _01045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_184_clock clknet_5_30_0_clock clknet_leaf_184_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12635_ _00514_ clknet_leaf_211_clock u2.mem\[32\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12566_ _00445_ clknet_leaf_98_clock u2.mem\[27\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08444__A1 _03629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07247__A2 _02721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12686__CLK clknet_leaf_216_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11517_ _05674_ u2.mem\[169\]\[3\] _05700_ _05704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06455__B1 _01948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12497_ _00376_ clknet_leaf_175_clock u2.mem\[23\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_199_clock clknet_5_31_0_clock clknet_leaf_199_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_156_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11448_ _05631_ u2.mem\[165\]\[3\] _05655_ _05659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08930__S _04079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_5_14_0_clock_I clknet_4_7_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11051__I0 _05392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11379_ _05583_ u2.mem\[161\]\[0\] _05616_ _05617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06758__A1 u2.mem\[159\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07955__B1 _02426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06758__B2 u2.mem\[149\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13118_ _00997_ clknet_leaf_276_clock u2.mem\[62\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_122_clock clknet_5_14_0_clock clknet_leaf_122_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_263_clock_I clknet_5_22_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_2_2__f_clock_a_I clknet_0_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13049_ _00928_ clknet_leaf_343_clock u2.mem\[57\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07707__B1 _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12066__CLK clknet_leaf_374_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07345__I _02504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13311__CLK clknet_leaf_363_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07183__B2 u2.mem\[12\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07610_ u2.mem\[17\]\[8\] _03079_ _03080_ u2.mem\[24\]\[8\] _03081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_137_clock clknet_5_14_0_clock clknet_leaf_137_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08590_ _03855_ _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_82_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11106__I1 u2.mem\[144\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07541_ u2.mem\[8\]\[7\] _02860_ _02861_ u2.mem\[4\]\[7\] _03013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_90_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13461__CLK clknet_leaf_360_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07472_ u2.mem\[58\]\[6\] _02811_ _02812_ u2.mem\[36\]\[6\] _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07080__I _02558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09211_ _04147_ _04265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06694__B1 _02177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06423_ _01923_ _01924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09142_ _04220_ _00383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07238__A2 _02659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06354_ u2.mem\[187\]\[4\] _01634_ _01637_ u2.mem\[192\]\[4\] _01857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09483__I0 _04384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09001__S _04124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09073_ _04180_ _04122_ _04181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11290__I0 _05550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10147__S _04846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06285_ u2.mem\[145\]\[2\] _01639_ _01642_ u2.mem\[163\]\[2\] u2.mem\[165\]\[2\]
+ _01645_ _01790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_129_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09936__S _04719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08024_ _03480_ _03481_ _03484_ _03485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__09235__I0 _04281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06749__A1 u2.mem\[185\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06749__B2 u2.mem\[173\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12409__CLK clknet_leaf_124_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09975_ _04689_ u2.mem\[43\]\[3\] _04740_ _04744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_77_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08926_ _04078_ _00309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11345__I1 u2.mem\[158\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08857_ _04035_ u2.mem\[17\]\[9\] _04033_ _04036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12559__CLK clknet_leaf_159_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07808_ _02482_ _03275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08788_ _03991_ _00258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07739_ u2.mem\[45\]\[11\] _03099_ _03100_ u2.mem\[34\]\[11\] _03207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10750_ _03707_ _05222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09409_ _04390_ _00480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10681_ _05101_ u2.mem\[60\]\[3\] _05174_ _05178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12420_ _00299_ clknet_leaf_102_clock u2.mem\[18\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07229__A2 _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09474__I0 _04375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12351_ _00230_ clknet_leaf_160_clock u2.mem\[14\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09846__S _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11302_ _05569_ _01194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12282_ _00161_ clknet_leaf_118_clock u2.mem\[9\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11233_ _05517_ u2.mem\[151\]\[5\] _05519_ _05526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07874__B _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11733__A1 _05354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12089__CLK clknet_2_2__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11164_ _05472_ u2.mem\[147\]\[5\] _05474_ _05481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13334__CLK clknet_leaf_3_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09529__I1 u2.mem\[32\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10115_ _04801_ u2.mem\[46\]\[8\] _04830_ _04831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11095_ _05438_ _01118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_54_clock clknet_5_12_0_clock clknet_leaf_54_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11336__I1 u2.mem\[158\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10046_ _04785_ _00722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13484__CLK clknet_leaf_306_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11616__S _05760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08197__S _03608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_69_clock clknet_5_9_0_clock clknet_leaf_69_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_17_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11997_ _00009_ clknet_leaf_34_clock u2.mem\[0\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07114__B _02458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10847__I0 _05200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10948_ _04134_ _05345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06509__I _01993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08925__S _04074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10879_ _04994_ _05301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06140__A2 _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12618_ _00497_ clknet_leaf_137_clock u2.mem\[30\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09465__I0 _04366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12549_ _00428_ clknet_leaf_100_clock u2.mem\[26\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08660__S _03905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06244__I _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06070_ _01552_ _01576_ _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07640__A2 _03033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_0_clock_I clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09555__I _04150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09760_ _04613_ _00608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06972_ _02447_ _02449_ _02430_ _02450_ _02451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_113_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12701__CLK clknet_leaf_222_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08711_ _03944_ _00228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09691_ _04561_ _00591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11526__S _05709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08642_ _03896_ _00207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08573_ _03797_ u2.mem\[11\]\[0\] _03856_ _03857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_165_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07524_ u2.mem\[61\]\[7\] _02899_ _02900_ u2.mem\[63\]\[7\] _02996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_63_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07459__A2 _02866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06419__I _01913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07455_ u2.mem\[6\]\[5\] _02927_ _02928_ u2.mem\[47\]\[5\] _02929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__13207__CLK clknet_leaf_300_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06131__A2 _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06406_ u2.mem\[147\]\[5\] _01675_ _01679_ u2.mem\[169\]\[5\] _01907_ _01908_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_10_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09456__I0 _04356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07386_ _02611_ _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09125_ _04148_ u2.mem\[23\]\[6\] _04208_ _04211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06337_ _01829_ _01834_ _01835_ _01840_ _01841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_124_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09056_ _04123_ _04168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__12231__CLK clknet_leaf_54_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06154__I _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07631__A2 _03099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06268_ _01772_ _01773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_163_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08007_ u2.active_mem\[15\] _03461_ _03462_ u2.active_mem\[14\] _03470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_116_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06199_ u2.mem\[190\]\[0\] _01703_ _01705_ u2.mem\[194\]\[0\] _01706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_150_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07919__B1 _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05993__I row_col_select_trans.data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11566__I1 u2.mem\[172\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_2_0_clock_I clknet_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07395__A1 u2.mem\[32\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12381__CLK clknet_leaf_232_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_6_clock_I clknet_5_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10404__I _03686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09958_ _04718_ _04734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_clkbuf_leaf_159_clock_I clknet_5_27_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08909_ _04044_ u2.mem\[18\]\[13\] _04066_ _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_4136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07147__A1 _02560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09889_ _04689_ u2.mem\[41\]\[3\] _04683_ _04690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_4147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11920_ _05953_ _01428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11851_ _05911_ u2.mem\[190\]\[3\] _05905_ _05912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11235__I _05442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10802_ u2.mem\[63\]\[0\] _03491_ _05253_ _05254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08745__S _03962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_211_clock_I clknet_5_28_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11782_ _05868_ u2.mem\[186\]\[1\] _05866_ _05869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13521_ _01400_ clknet_leaf_4_clock u2.mem\[190\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10733_ _05210_ _00984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06122__A2 _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11171__S _05484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13452_ _01331_ clknet_leaf_358_clock u2.mem\[178\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08544__I _03834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10664_ _05121_ u2.mem\[59\]\[12\] _05167_ _05168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07870__A2 _03333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_19_0_clock clknet_4_9_0_clock clknet_5_19_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_90_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12403_ _00282_ clknet_leaf_109_clock u2.mem\[17\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11254__I0 _05505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13383_ _01262_ clknet_leaf_318_clock u2.mem\[167\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_167_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10595_ _03720_ _05128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12334_ _00213_ clknet_leaf_234_clock u2.mem\[13\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06999__I _02368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12265_ _00144_ clknet_leaf_55_clock u2.mem\[8\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12724__CLK clknet_leaf_25_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09375__I _04357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11216_ _05515_ _01162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12196_ _00075_ clknet_leaf_22_clock u2.mem\[4\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_150_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11147_ _05470_ u2.mem\[146\]\[4\] _05461_ _05471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_1_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11309__I1 u2.mem\[156\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11078_ _05427_ _01112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10029_ _04705_ u2.mem\[44\]\[10\] _04772_ _04775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_48_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07623__I _02611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12104__CLK clknet_leaf_25_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06361__A2 _01708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07310__A1 u2.mem\[45\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06113__A2 _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07240_ u2.mem\[43\]\[2\] _02505_ _02508_ u2.mem\[20\]\[2\] _02717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_31_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08454__I _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07171_ u2.mem\[50\]\[1\] _02647_ _02648_ u2.mem\[51\]\[1\] _02649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06122_ u2.mem\[171\]\[0\] _01611_ _01615_ u2.mem\[157\]\[0\] _01628_ _01629_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_69_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07613__A2 _03082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06053_ _01558_ _01559_ _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10425__S _05021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09285__I _04312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06702__I _02100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09610__I0 _04489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10224__I _04886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09812_ _04638_ _04644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06719__A4 _02202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_160_clock_I clknet_5_27_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06955_ _02373_ _02434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_09743_ _04600_ _00604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11256__S _05537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06858__B _02337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09674_ _04478_ u2.mem\[36\]\[6\] _04549_ _04552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08629__I _03878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06886_ _02364_ _02365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08625_ _03812_ u2.mem\[12\]\[6\] _03884_ _03887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_54_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07144__A4 _02442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11055__I _05412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08556_ _03819_ u2.mem\[10\]\[9\] _03845_ _03847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08565__S _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07507_ u2.mem\[15\]\[7\] _02794_ _02795_ u2.mem\[13\]\[7\] _02979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_161_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11484__I0 _05668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08487_ _03801_ u2.mem\[9\]\[1\] _03799_ _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07438_ u2.mem\[9\]\[5\] _02838_ _02839_ u2.mem\[25\]\[5\] _02912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_168_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_20_0_clock clknet_4_10_0_clock clknet_5_20_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_126_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_85_clock_I clknet_5_9_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07369_ _02834_ _02837_ _02840_ _02843_ _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__12747__CLK clknet_leaf_271_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09108_ _04177_ u2.mem\[22\]\[15\] _04197_ _04201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10380_ _04126_ _04991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09039_ _04123_ _04155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_151_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09195__I _04127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12050_ data_in_trans\[0\].A clknet_leaf_378_clock data_in_trans\[0\].data_sync vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06612__I _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09601__I0 _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11001_ _05378_ _01084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07907__A3 _03367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12127__CLK clknet_leaf_36_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_6_0_clock_I clknet_3_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12952_ _00831_ clknet_leaf_148_clock u2.mem\[51\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11711__I1 u2.mem\[181\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06487__C _01964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11903_ u2.mem\[192\]\[11\] _03524_ _05942_ _05944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12883_ _00762_ clknet_leaf_69_clock u2.mem\[47\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07540__B2 u2.mem\[48\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12277__CLK clknet_leaf_104_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_362_clock_I clknet_5_4_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11834_ _05900_ _01395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13522__CLK clknet_leaf_4_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11765_ _05858_ _01368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13504_ _01383_ clknet_leaf_333_clock u2.mem\[187\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10716_ _05198_ u2.mem\[61\]\[1\] _05196_ _05199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08274__I _03490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11696_ _05815_ _01342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11227__I0 _05508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10309__I _04943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13435_ _01314_ clknet_leaf_366_clock u2.mem\[176\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10647_ _05158_ _00950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13366_ _01245_ clknet_leaf_373_clock u2.mem\[164\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10578_ _05116_ _00923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12317_ _00196_ clknet_leaf_186_clock u2.mem\[12\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13297_ _01176_ clknet_leaf_382_clock u2.mem\[153\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12248_ _00127_ clknet_leaf_56_clock u2.mem\[7\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10044__I _04783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12179_ _00058_ clknet_leaf_77_clock u2.mem\[3\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_150_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06031__B2 _01516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06582__A2 _02018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13052__CLK clknet_leaf_274_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06740_ _02219_ _02220_ _02221_ _02222_ _02223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06671_ _02155_ _02156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08410_ _03667_ u2.mem\[7\]\[2\] _03753_ _03756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_91_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09390_ _04377_ _00474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08341_ _03708_ _03709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11466__I0 _05671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09284__A1 _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_107_clock_I clknet_5_11_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06098__A1 u2.mem\[175\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07295__B1 _02582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08184__I _03584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08272_ _03579_ u2.mem\[4\]\[15\] _03649_ _03653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06098__B2 u2.mem\[159\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07223_ u2.mem\[32\]\[2\] _02385_ _02397_ u2.mem\[2\]\[2\] _02700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07047__B1 _02525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07154_ _01544_ _02361_ _02535_ _02632_ _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_146_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09831__I0 _04605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06105_ _01557_ _01612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_156_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07085_ _02563_ _02564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06270__A1 u2.mem\[171\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06036_ u3.data u3.enable net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06432__I _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06270__B2 u2.mem\[157\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08011__A2 _03473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input38_I row_select_a[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07987_ _03447_ _03448_ _03449_ _03450_ _03451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06588__B _01995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06938_ _02390_ _02400_ _02416_ _02417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_09726_ _04587_ _00600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13545__CLK clknet_leaf_40_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09657_ _04541_ _00577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06869_ _01579_ _01985_ _02348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_55_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08608_ _03630_ _03773_ _03876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09588_ _04467_ u2.mem\[34\]\[1\] _04501_ _04503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08295__S _03659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08539_ _03837_ _00163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08322__I0 _03692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11550_ _05725_ _01286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08094__I _03491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06607__I _02091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10501_ _05023_ u2.mem\[55\]\[13\] _05066_ _05068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11481_ _05682_ _05683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_155_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13220_ _01099_ clknet_leaf_299_clock u2.mem\[140\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09918__I _04682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10432_ _05028_ _00865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08822__I _03655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09822__I0 _04592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13151_ _01030_ clknet_leaf_260_clock u2.mem\[128\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_163_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10363_ _04911_ u2.mem\[52\]\[11\] _04976_ _04980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_309_clock_I clknet_5_20_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_174_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12102_ _01500_ clknet_leaf_43_clock u2.active_mem\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06261__B2 u2.mem\[160\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13082_ _00961_ clknet_leaf_341_clock u2.mem\[59\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10294_ _04940_ _00815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12033_ net41 clknet_2_3__leaf_clock_a row_select_trans\[4\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13075__CLK clknet_leaf_25_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10196__I0 _04806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08002__A2 _03461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07761__A1 u2.mem\[61\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09889__I0 _04689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07173__I _02500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12935_ _00814_ clknet_leaf_147_clock u2.mem\[50\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06316__A2 _01734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11624__S _05771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12912__CLK clknet_leaf_162_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12866_ _00745_ clknet_leaf_154_clock u2.mem\[46\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11448__I0 _05631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11817_ _05870_ u2.mem\[188\]\[2\] _05888_ _05891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08069__A2 _03518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12797_ _00676_ clknet_leaf_204_clock u2.mem\[42\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07277__B1 _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11748_ _04223_ _05847_ _05848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_18_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11679_ _05805_ _01335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08732__I _03940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13418_ _01297_ clknet_leaf_314_clock u2.mem\[173\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08616__I1 u2.mem\[12\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09813__I0 _04579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13418__CLK clknet_leaf_314_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13349_ _01228_ clknet_leaf_3_clock u2.mem\[161\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06252__I _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07595__A4 _03065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07910_ u2.mem\[32\]\[14\] _03252_ _03253_ u2.mem\[2\]\[14\] _03375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_29_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08890_ _04057_ _00294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10187__I0 _04797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07201__B1 _02577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07841_ _02581_ _03308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13568__CLK clknet_leaf_13_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_33_clock_I clknet_5_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07772_ u2.mem\[17\]\[11\] _03079_ _03080_ u2.mem\[24\]\[11\] _03240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07083__I _02363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09511_ _04373_ u2.mem\[32\]\[7\] _04448_ _04452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06723_ u2.mem\[167\]\[2\] _02059_ _02062_ u2.mem\[183\]\[2\] _02206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_65_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11687__I0 _05786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07504__A1 u2.mem\[40\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12592__CLK clknet_leaf_161_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07504__B2 u2.mem\[30\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09442_ _04410_ _00493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06654_ _02132_ _02135_ _02138_ _02139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_168_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07811__I _02489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09373_ _04365_ _00469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06585_ _02027_ _02000_ _02070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_258_clock_I clknet_5_19_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08324_ data_in_trans\[9\].data_sync _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07268__B1 _02639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08255_ _03643_ _00073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07206_ u2.mem\[23\]\[1\] _02682_ _02683_ u2.mem\[22\]\[1\] _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_105_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08186_ _03601_ _00046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09804__I0 _04565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07137_ _02459_ _02614_ _02615_ _02458_ _02616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__13098__CLK clknet_leaf_340_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_310_clock_I clknet_5_20_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08232__A2 mem_address_trans\[0\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07586__A4 _03056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07068_ _02418_ _02510_ _02511_ _02546_ _02547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06794__A2 _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11709__S _05817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06019_ _01514_ _01521_ _01527_ _01516_ _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_160_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10613__S _05136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10178__I0 _04788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09473__I _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07743__A1 _03207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08791__I0 _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12935__CLK clknet_leaf_147_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11678__I0 _05794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09709_ _04574_ _00596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10981_ _05367_ _01075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11444__S _05655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12720_ _00599_ clknet_leaf_248_clock u2.mem\[37\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10350__I0 _04898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12651_ _00530_ clknet_leaf_213_clock u2.mem\[33\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11602_ _05757_ _01306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12582_ _00461_ clknet_leaf_100_clock u2.mem\[28\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12315__CLK clknet_leaf_185_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11533_ _05714_ _01280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11464_ _03498_ _05670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10415_ _05016_ u2.mem\[53\]\[10\] _05012_ _05017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13203_ _01082_ clknet_leaf_294_clock u2.mem\[137\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11395_ _05626_ _01230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09271__I1 u2.mem\[26\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06234__A1 u2.mem\[170\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10346_ _04970_ _00837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12465__CLK clknet_leaf_173_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06234__B2 u2.mem\[156\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13134_ _01013_ clknet_leaf_262_clock u2.mem\[63\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13065_ _00944_ clknet_leaf_339_clock u2.mem\[58\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10277_ _04900_ u2.mem\[50\]\[6\] _04928_ _04931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_79_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10523__S _05078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12016_ mem_address_trans\[5\].A clknet_leaf_315_clock mem_address_trans\[5\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11905__I1 _03527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06537__A2 _01997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08928__S _04079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12918_ _00797_ clknet_leaf_87_clock u2.mem\[49\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07498__B1 _02928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10341__I0 _04889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12849_ _00728_ clknet_leaf_154_clock u2.mem\[45\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09759__S _04606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06247__I _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06370_ _01870_ _01871_ _01872_ _01873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_37_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08663__S _03905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_352_clock clknet_5_4_0_clock clknet_leaf_352_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08837__I1 u2.mem\[17\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13240__CLK clknet_leaf_289_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09558__I _04153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08040_ _03498_ _03499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12808__CLK clknet_leaf_130_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_367_clock clknet_5_1_0_clock clknet_leaf_367_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_31_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13390__CLK clknet_leaf_364_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09991_ _04705_ u2.mem\[43\]\[10\] _04750_ _04753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11529__S _05709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06776__A2 _02075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07973__B2 u2.mem\[63\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08942_ _04087_ _00316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12958__CLK clknet_leaf_197_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08873_ _04046_ u2.mem\[17\]\[14\] _04042_ _04047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07824_ u2.mem\[61\]\[12\] _03132_ _03133_ u2.mem\[63\]\[12\] _03291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_3809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10580__I0 _05117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07755_ u2.mem\[44\]\[11\] _03122_ _03123_ u2.mem\[42\]\[11\] _03223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_305_clock clknet_5_20_0_clock clknet_leaf_305_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_56_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06706_ _02184_ _02188_ _02189_ _02190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_65_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10332__I0 _04918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07686_ _02628_ _03156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_129_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09425_ _04395_ _04401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06637_ _02064_ _02018_ _02122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12338__CLK clknet_leaf_159_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06161__B1 _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06700__A2 _02065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06157__I _01663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09356_ _04283_ u2.mem\[28\]\[14\] _04351_ _04354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08573__S _03856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06568_ _02052_ _01999_ _02053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_139_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08307_ _03681_ _00087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09287_ _04314_ _00434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06499_ row_select_trans\[0\].data_sync _01984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08238_ _03633_ _03634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_14_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06464__A1 u2.mem\[193\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12488__CLK clknet_leaf_125_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08372__I _03726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06464__B2 u2.mem\[194\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08169_ _03557_ u2.mem\[2\]\[5\] _03590_ _03592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10407__I _03690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10399__I0 _05005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10200_ _04864_ _04880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06216__A1 u2.mem\[173\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06216__B2 u2.mem\[185\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11180_ _05490_ _01151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06767__A2 _02129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10131_ _04839_ _00753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10343__S _04966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10062_ _04796_ _00727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10142__I _04840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09931__I _04718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07192__A2 _02537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13113__CLK clknet_leaf_39_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08516__I0 _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10323__I0 _04909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10964_ _05357_ _01068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12703_ _00582_ clknet_leaf_238_clock u2.mem\[36\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13263__CLK clknet_leaf_286_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10895_ _05299_ u2.mem\[131\]\[1\] _05310_ _05312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12634_ _00513_ clknet_leaf_115_clock u2.mem\[31\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06067__I col_select_trans\[1\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11823__I0 _05876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12565_ _00444_ clknet_leaf_105_clock u2.mem\[27\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08444__A2 _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09378__I _04144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11516_ _05703_ _01274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08282__I _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12496_ _00375_ clknet_leaf_175_clock u2.mem\[23\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11447_ _05658_ _01250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06207__A1 _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_166_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11378_ _05615_ _05616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_125_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07955__A1 u2.mem\[27\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06758__A2 _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_206_clock_I clknet_5_31_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10329_ _04960_ _00830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13117_ _00996_ clknet_leaf_276_clock u2.mem\[62\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_18_0_clock_I clknet_4_9_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06530__I _02014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13048_ _00927_ clknet_leaf_344_clock u2.mem\[57\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07183__A2 _02659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09841__I _04660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06391__B1 _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07540_ u2.mem\[39\]\[7\] _02857_ _02858_ u2.mem\[48\]\[7\] _03012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_35_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10314__I0 _04900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07361__I _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09180__I0 _04171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07471_ u2.mem\[53\]\[6\] _02808_ _02809_ u2.mem\[56\]\[6\] _02944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_34_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_291_clock clknet_5_21_0_clock clknet_leaf_291_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_62_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09210_ _04264_ _00407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06422_ _01922_ _01916_ _01923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06694__A1 u2.mem\[149\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08393__S _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12630__CLK clknet_leaf_95_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09141_ _04171_ u2.mem\[23\]\[13\] _04218_ _04220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06353_ u2.mem\[193\]\[4\] _01731_ _01734_ u2.mem\[177\]\[4\] _01856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10428__S _05021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09072_ _04179_ _04180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11290__I1 u2.mem\[155\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06284_ u2.mem\[166\]\[2\] _01757_ _01758_ u2.mem\[161\]\[2\] _01788_ _01789_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_50_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08023_ _03482_ _03483_ _03484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09235__I1 u2.mem\[25\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12780__CLK clknet_leaf_268_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09974_ _04743_ _00692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12010__CLK clknet_leaf_315_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09952__S _04729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13136__CLK clknet_leaf_330_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08925_ _04021_ u2.mem\[19\]\[3\] _04074_ _04078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08856_ _03696_ _04035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input20_I data_in_a[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07174__A2 _02650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07807_ _02475_ _03274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08787_ _03899_ u2.mem\[16\]\[0\] _03990_ _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12160__CLK clknet_leaf_236_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05999_ _01507_ _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13286__CLK clknet_leaf_381_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10305__I0 _04891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07738_ _01962_ _03017_ _03185_ _03206_ _01487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09171__I0 _04158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_259_clock clknet_5_19_0_clock clknet_leaf_259_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_77_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07669_ u2.mem\[57\]\[9\] _03137_ _03138_ u2.mem\[41\]\[9\] _03139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_13_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11722__S _05827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09408_ _04389_ u2.mem\[29\]\[14\] _04385_ _04390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07882__B1 _02525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10680_ _05177_ _00964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_2_clock_I clknet_5_0_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_155_clock_I clknet_5_24_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09339_ _04344_ _00456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09198__I _04131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06437__A1 _01773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12350_ _00229_ clknet_leaf_208_clock u2.mem\[14\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06437__B2 _01935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11301_ _05544_ u2.mem\[156\]\[0\] _05568_ _05569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12281_ _00160_ clknet_leaf_118_clock u2.mem\[9\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11232_ _05525_ _01168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08830__I _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07937__B2 u2.mem\[25\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08985__I0 _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11733__A2 _05808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11169__S _05484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11163_ _05480_ _01144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10792__I0 _05222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10114_ _04819_ _04830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09862__S _04671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11094_ _05426_ u2.mem\[143\]\[2\] _05435_ _05438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08737__I0 _03936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12503__CLK clknet_leaf_125_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_15_0_clock clknet_4_7_0_clock clknet_5_15_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_10045_ _04782_ u2.mem\[45\]\[0\] _04784_ _04785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07165__A2 _02457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07181__I _02520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11996_ _00008_ clknet_leaf_334_clock u2.mem\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09162__I0 _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10947_ _05344_ _01064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11632__S _05770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06676__B2 u2.mem\[147\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10878_ _05300_ _01039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09102__S _04197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12617_ _00496_ clknet_leaf_134_clock u2.mem\[30\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13009__CLK clknet_leaf_253_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07130__B _02401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07625__B1 _02928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08941__S _04084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12548_ _00427_ clknet_leaf_100_clock u2.mem\[26\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06979__A2 _02391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12479_ _00358_ clknet_leaf_176_clock u2.mem\[22\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12033__CLK clknet_2_3__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07928__A1 _03389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08976__I0 _04032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_357_clock_I clknet_5_5_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10783__I0 _05213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06971_ _02394_ _02450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_100_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12183__CLK clknet_leaf_62_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08728__I0 _03927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08710_ _03909_ u2.mem\[14\]\[2\] _03941_ _03944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09690_ _04494_ u2.mem\[36\]\[13\] _04559_ _04561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08388__S _03737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09571__I _04166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08641_ _03828_ u2.mem\[12\]\[13\] _03894_ _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08572_ _03855_ _03856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_78_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09153__I0 _04128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07523_ _02978_ _02984_ _02989_ _02994_ _02995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_22_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08900__I0 _04035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07454_ _02623_ _02928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06667__A1 _02104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06405_ _01904_ _01905_ _01906_ _01907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06863__C col_select_trans\[4\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10158__S _04851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07385_ _02609_ _02860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11341__I _05513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09124_ _04210_ _00375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09947__S _04724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06336_ u2.mem\[147\]\[3\] _01676_ _01680_ u2.mem\[169\]\[3\] _01839_ _01840_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_52_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06435__I _01920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09055_ _04166_ _04167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07092__A1 _02439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06267_ u2.mem\[0\]\[2\] _01772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_11_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08006_ u2.active_mem\[12\] _03458_ _03459_ u2.active_mem\[13\] _03469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_104_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06198_ _01704_ _01705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08967__I0 _04023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12526__CLK clknet_leaf_198_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10774__I0 _05204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09957_ _04733_ _00685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07934__A4 _03398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_183_clock clknet_5_27_0_clock clknet_leaf_183_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08719__I0 _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08908_ _04067_ _00302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_3_6_0_clock_I clknet_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09888_ _04575_ _04689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07147__A2 _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_81_clock_I clknet_5_8_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09392__I0 _04378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12676__CLK clknet_leaf_83_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08839_ _03674_ _04023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06355__B1 _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10420__I _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11850_ _03669_ _05911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_198_clock clknet_5_31_0_clock clknet_leaf_198_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10801_ _05252_ _05253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10829__I1 _03527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11781_ _03661_ _05868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13520_ _01399_ clknet_leaf_5_clock u2.mem\[190\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07855__B1 _03156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11651__A1 _05295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10732_ _05209_ u2.mem\[61\]\[6\] _05205_ _05210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_121_clock clknet_5_14_0_clock clknet_leaf_121_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13451_ _01330_ clknet_leaf_322_clock u2.mem\[178\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10663_ _05151_ _05167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_139_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11251__I _05536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12402_ _00281_ clknet_leaf_171_clock u2.mem\[17\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12056__CLK clknet_leaf_376_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07607__B1 _02916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11254__I1 u2.mem\[153\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08761__S _03972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13382_ _01261_ clknet_leaf_319_clock u2.mem\[167\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10594_ _05127_ _00928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13301__CLK clknet_leaf_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12333_ _00212_ clknet_leaf_210_clock u2.mem\[13\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_136_clock clknet_5_14_0_clock clknet_leaf_136_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_126_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06830__A1 u2.mem\[150\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12264_ _00143_ clknet_leaf_55_clock u2.mem\[8\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08958__I0 _04010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11215_ _05514_ u2.mem\[150\]\[4\] _05501_ _05515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12195_ _00074_ clknet_leaf_22_clock u2.mem\[4\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13451__CLK clknet_leaf_322_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10765__I0 _05194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09592__S _04501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11146_ _05348_ _05470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11077_ _05426_ u2.mem\[142\]\[2\] _05422_ _05427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09391__I _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10028_ _04774_ _00715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06897__A1 _02352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11979_ _05987_ _01453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06649__A1 _02014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07310__A2 _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09767__S _04618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07170_ _02494_ _02648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06121_ _01620_ _01625_ _01627_ _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__12549__CLK clknet_leaf_100_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06821__A1 u2.mem\[185\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06052_ col_select_trans\[3\].data_sync _01559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_160_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09811_ _04643_ _00629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_103_clock_I clknet_5_10_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09742_ _04599_ u2.mem\[37\]\[10\] _04593_ _04600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10441__S _05030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06954_ _02369_ _02433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_132_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09673_ _04551_ _00583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06885_ _01988_ _01997_ _02364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08624_ _03886_ _00199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08555_ _03846_ _00170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07506_ _02974_ _02975_ _02976_ _02977_ _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__12079__CLK clknet_2_0__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08486_ _03662_ _03801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11484__I1 u2.mem\[167\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13324__CLK clknet_leaf_322_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07437_ u2.mem\[29\]\[5\] _02835_ _02836_ u2.mem\[11\]\[5\] _02911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_4_13_0_clock_I clknet_3_6_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_28_clock_I clknet_5_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_53_clock clknet_5_12_0_clock clknet_leaf_53_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_164_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07368_ u2.mem\[28\]\[4\] _02841_ _02842_ u2.mem\[31\]\[4\] _02843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_6_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09107_ _04200_ _00368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06319_ u2.mem\[175\]\[3\] _01602_ _01632_ u2.mem\[188\]\[3\] _01823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07299_ u2.mem\[52\]\[3\] _02599_ _02601_ u2.mem\[21\]\[3\] _02775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_108_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13474__CLK clknet_leaf_308_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06812__A1 u2.mem\[179\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09038_ _04153_ _04154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06812__B2 u2.mem\[191\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_68_clock clknet_5_9_0_clock clknet_leaf_68_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_85_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11000_ _05349_ u2.mem\[137\]\[4\] _05372_ _05378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12951_ _00830_ clknet_leaf_147_clock u2.mem\[51\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06328__B1 _01714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11902_ _05943_ _01420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08756__S _03967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12882_ _00761_ clknet_leaf_243_clock u2.mem\[47\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_305_clock_I clknet_5_20_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11833_ _05872_ u2.mem\[189\]\[3\] _05896_ _05900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11764_ _05825_ u2.mem\[185\]\[0\] _05857_ _05858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13503_ _01382_ clknet_leaf_346_clock u2.mem\[187\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10715_ _04991_ _05198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11695_ _05796_ u2.mem\[180\]\[4\] _05809_ _05815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11227__I1 u2.mem\[151\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06075__I _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13434_ _01313_ clknet_leaf_353_clock u2.mem\[175\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10646_ _05103_ u2.mem\[59\]\[4\] _05157_ _05158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07056__A1 _02438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13365_ _01244_ clknet_leaf_373_clock u2.mem\[164\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10577_ _05115_ u2.mem\[57\]\[9\] _05113_ _05116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12316_ _00195_ clknet_leaf_185_clock u2.mem\[12\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06803__A1 u2.mem\[165\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06803__B2 u2.mem\[163\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12841__CLK clknet_leaf_130_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13296_ _01175_ clknet_leaf_370_clock u2.mem\[152\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08005__B1 _03467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12247_ _00126_ clknet_leaf_56_clock u2.mem\[7\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07359__A2 _02675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12178_ _00057_ clknet_leaf_239_clock u2.mem\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11357__S _05597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11129_ _05458_ _01132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09356__I0 _04283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07634__I _02419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06319__B1 _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06670_ _02022_ _02052_ _02155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12221__CLK clknet_leaf_226_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10910__I0 _05299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09108__I0 _04177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13347__CLK clknet_leaf_14_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11092__S _05435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08340_ _03707_ _03708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08271_ _03652_ _00080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13497__CLK clknet_leaf_329_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07222_ u2.mem\[45\]\[2\] _02633_ _02634_ u2.mem\[34\]\[2\] _02699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_121_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07153_ _02557_ _02584_ _02608_ _02631_ _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06104_ _01610_ _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07084_ _02560_ _02561_ _02417_ _02562_ _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_161_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07062__A4 _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06035_ _01543_ _00000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06270__A2 _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10729__I0 _05207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09595__I0 _04473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_254_clock_I clknet_5_19_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11267__S _05546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07986_ u2.mem\[18\]\[15\] _03318_ _03319_ u2.mem\[19\]\[15\] _03450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_75_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09347__I0 _04274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09725_ _04586_ u2.mem\[37\]\[6\] _04580_ _04587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06937_ _02349_ _02415_ _02416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_27_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11154__I0 _05460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12102__D _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09656_ _04498_ u2.mem\[35\]\[15\] _04537_ _04541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06868_ _02346_ _02347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10901__I0 _05305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08607_ _03875_ _00193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09587_ _04502_ _00546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06799_ u2.mem\[184\]\[4\] _02071_ _01993_ _02280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12714__CLK clknet_leaf_146_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05999__I _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08538_ _03801_ u2.mem\[10\]\[1\] _03835_ _03837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_24_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11606__A1 _04416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07286__A1 _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08469_ _03790_ _00140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06628__A4 _02112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10500_ _05067_ _00894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11480_ _05354_ _05645_ _05682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__12864__CLK clknet_leaf_154_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07038__A1 _02395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10431_ _05027_ u2.mem\[53\]\[15\] _05021_ _05028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13150_ _01029_ clknet_leaf_281_clock u2.mem\[128\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10362_ _04979_ _00844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06797__B1 _02053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12101_ _01499_ clknet_leaf_246_clock u2.active_mem\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10293_ _04916_ u2.mem\[50\]\[13\] _04938_ _04940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13081_ _00960_ clknet_leaf_340_clock u2.mem\[59\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09586__I0 _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12032_ row_select_trans\[3\].A clknet_leaf_303_clock row_select_trans\[3\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11177__S _05483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12244__CLK clknet_leaf_73_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07454__I _02623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09338__I0 _04265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07761__A2 _03132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12012__D mem_address_trans\[3\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11905__S _05942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12934_ _00813_ clknet_leaf_63_clock u2.mem\[50\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07513__A2 _02880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12865_ _00744_ clknet_leaf_154_clock u2.mem\[46\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12394__CLK clknet_leaf_140_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06721__B1 _02171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11816_ _05890_ _01387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11448__I1 u2.mem\[165\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12796_ _00675_ clknet_leaf_204_clock u2.mem\[42\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11747_ _05768_ _05847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11640__S _05779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11678_ _05794_ u2.mem\[179\]\[3\] _05801_ _05805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_174_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13417_ _01296_ clknet_leaf_314_clock u2.mem\[173\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10629_ _05124_ u2.mem\[58\]\[13\] _05146_ _05148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07629__I _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13348_ _01227_ clknet_leaf_14_clock u2.mem\[161\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13279_ _01158_ clknet_leaf_380_clock u2.mem\[150\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06004__A2 _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07201__B2 u2.mem\[25\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07840_ _02579_ _03307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07364__I _02576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09329__I0 _04256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09780__S _04623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07752__A2 _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07771_ u2.mem\[23\]\[11\] _03148_ _03149_ u2.mem\[22\]\[11\] _03239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_133_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09510_ _04451_ _00520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12737__CLK clknet_leaf_247_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11815__S _05888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06722_ u2.mem\[164\]\[2\] _02051_ _02054_ u2.mem\[178\]\[2\] _02205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11687__I1 u2.mem\[180\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09441_ _04382_ u2.mem\[30\]\[11\] _04406_ _04410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06653_ u2.mem\[153\]\[0\] _02136_ _02137_ u2.mem\[160\]\[0\] _02138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09372_ _04364_ u2.mem\[29\]\[3\] _04358_ _04365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06708__I _02047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06584_ u2.mem\[171\]\[0\] _02066_ _02068_ u2.mem\[157\]\[0\] _02069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_36_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12887__CLK clknet_leaf_57_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07268__A1 u2.mem\[27\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08323_ _03694_ _00090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08254_ _03561_ u2.mem\[4\]\[7\] _03639_ _03643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07205_ _02595_ _02683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12117__CLK clknet_leaf_348_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08185_ _03572_ u2.mem\[2\]\[12\] _03600_ _03601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_174_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_146_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07136_ _02480_ _02615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_118_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06779__B1 _02012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07067_ _02428_ _02377_ _02429_ _02546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_160_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12267__CLK clknet_leaf_194_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09754__I _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06018_ _01504_ _01524_ _01526_ _01527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07991__A2 _02622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13512__CLK clknet_leaf_354_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11375__I0 _05595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07743__A2 _03208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07969_ u2.mem\[49\]\[15\] _03283_ _03284_ u2.mem\[46\]\[15\] _03433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11725__S _05827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09708_ _04573_ u2.mem\[37\]\[2\] _04567_ _04574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11678__I1 u2.mem\[179\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10980_ _05340_ u2.mem\[136\]\[1\] _05365_ _05367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09639_ _04531_ _00569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10350__I1 u2.mem\[52\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12650_ _00529_ clknet_leaf_114_clock u2.mem\[32\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11601_ _05756_ u2.mem\[174\]\[4\] _05747_ _05757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_169_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12581_ _00460_ clknet_leaf_100_clock u2.mem\[28\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11532_ _05713_ u2.mem\[170\]\[2\] _05709_ _05714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08833__I _03666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11463_ _05669_ _01255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06482__A2 _01929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13042__CLK clknet_leaf_336_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07449__I _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13202_ _01081_ clknet_leaf_297_clock u2.mem\[137\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10414_ _03699_ _05016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11394_ _05623_ u2.mem\[162\]\[0\] _05625_ _05626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_174_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13133_ _01012_ clknet_leaf_282_clock u2.mem\[63\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10345_ _04893_ u2.mem\[52\]\[3\] _04966_ _04970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10804__S _05253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13192__CLK clknet_leaf_293_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13064_ _00943_ clknet_leaf_49_clock u2.mem\[58\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10276_ _04930_ _00807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12015_ net29 clknet_2_3__leaf_clock_a mem_address_trans\[5\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07195__B1 _02672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12917_ _00796_ clknet_leaf_88_clock u2.mem\[49\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10341__I1 u2.mem\[52\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12848_ _00727_ clknet_leaf_155_clock u2.mem\[45\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06528__I _02012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_202_clock_I clknet_5_29_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12779_ _00658_ clknet_leaf_265_clock u2.mem\[41\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06972__B _02430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09839__I _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_159_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07670__A1 _03134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09798__I0 _04612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13535__CLK clknet_leaf_334_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07422__B2 u2.mem\[20\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09990_ _04752_ _00699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08470__I0 _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07973__A2 _02553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08941_ _04037_ u2.mem\[19\]\[10\] _04084_ _04087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_48_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08872_ _03717_ _04046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07094__I _02446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07725__A2 _03074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07823_ _03259_ _03271_ _03280_ _03289_ _03290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_85_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07754_ _03218_ _03219_ _03220_ _03221_ _03222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__08918__I _04073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06705_ u2.mem\[165\]\[1\] _02076_ _02079_ u2.mem\[163\]\[1\] _02092_ u2.mem\[177\]\[1\]
+ _02189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_53_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07685_ _02626_ _03155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09424_ _04400_ _00485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06636_ _02120_ _02121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08854__S _04033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06161__A1 u2.mem\[180\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06161__B2 u2.mem\[150\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09355_ _04353_ _00463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06567_ _01990_ _02032_ _02052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13065__CLK clknet_leaf_339_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09749__I _04604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08306_ _03680_ u2.mem\[5\]\[5\] _03676_ _03681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08653__I _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09286_ _04246_ u2.mem\[27\]\[0\] _04313_ _04314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06498_ _01979_ _01924_ _01970_ _01980_ _01983_ _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_142_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06464__A2 _01942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08237_ _03629_ _03541_ _03632_ _03633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_20_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09685__S _04554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09789__I0 _04599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06173__I _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08168_ _03591_ _00038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07119_ _02463_ _02529_ _02530_ _02488_ _02598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__07413__A1 u2.mem\[58\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08461__I0 _03688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10624__S _05141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12902__CLK clknet_leaf_71_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08099_ mem_address_trans\[0\].data_sync _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_136_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10130_ _04817_ u2.mem\[46\]\[15\] _04835_ _04839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10061_ _04795_ u2.mem\[45\]\[5\] _04793_ _04796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_151_clock_I clknet_5_24_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10020__I0 _04696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07716__A2 _03174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09961__I0 _04712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10963_ _05335_ u2.mem\[135\]\[0\] _05356_ _05357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13408__CLK clknet_leaf_319_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12702_ _00581_ clknet_leaf_224_clock u2.mem\[36\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06688__C1 u2.mem\[193\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10894_ _05311_ _01044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12633_ _00512_ clknet_leaf_115_clock u2.mem\[31\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10087__I0 _04813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12564_ _00443_ clknet_leaf_90_clock u2.mem\[27\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12432__CLK clknet_leaf_169_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_11_0_clock clknet_4_5_0_clock clknet_5_11_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__11823__I1 u2.mem\[188\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13558__CLK clknet_leaf_16_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11515_ _05671_ u2.mem\[169\]\[2\] _05700_ _05703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_76_clock_I clknet_5_8_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06455__A2 _01942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12495_ _00374_ clknet_leaf_176_clock u2.mem\[23\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07179__I _02517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11446_ _05629_ u2.mem\[165\]\[2\] _05655_ _05658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06207__A2 _01618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12582__CLK clknet_leaf_100_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10534__S _05083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08452__I0 _03671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11377_ _05285_ _05606_ _05615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_154_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09394__I _04160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07955__A2 _02420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13116_ _00995_ clknet_leaf_276_clock u2.mem\[62\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10328_ _04913_ u2.mem\[51\]\[12\] _04959_ _04960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11339__I0 _05591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13047_ _00926_ clknet_leaf_340_clock u2.mem\[57\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_152_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10259_ _04614_ _04920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08939__S _04084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10011__I0 _04687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07707__A2 _03116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09952__I0 _04703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10711__A1 _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11365__S _05608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06391__A1 u2.mem\[159\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06391__B2 u2.mem\[149\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09704__I0 _04570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11511__I0 _05663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07470_ u2.mem\[54\]\[6\] _02883_ _02884_ u2.mem\[55\]\[6\] _02943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_leaf_353_clock_I clknet_5_5_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07340__B1 _02657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06421_ _01911_ _01922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_61_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09140_ _04219_ _00382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06352_ u2.mem\[158\]\[4\] _01728_ _01729_ u2.mem\[151\]\[4\] _01732_ u2.mem\[168\]\[4\]
+ _01855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_147_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06283_ _01785_ _01786_ _01787_ _01788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09071_ _03581_ _03749_ _04179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_163_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12925__CLK clknet_leaf_221_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08022_ mem_write_n_trans.data_sync mem_address_trans\[9\].data_sync mem_address_trans\[8\].data_sync
+ _03483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_163_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11578__I0 _05713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10444__S _05035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07817__I _02531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09973_ _04687_ u2.mem\[43\]\[2\] _04740_ _04743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08924_ _04077_ _00308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10243__I _04598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07159__B1 _02410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10002__I0 _04716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09943__I0 _04694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08855_ _04034_ _00282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11750__I0 _05825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12305__CLK clknet_leaf_161_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07806_ u2.mem\[54\]\[12\] _03116_ _03117_ u2.mem\[55\]\[12\] _03273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08786_ _03989_ _03990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06382__A1 u2.mem\[167\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07552__I _02409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05998_ _01505_ row_col_select_trans.data_sync _01506_ _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06382__B2 u2.mem\[183\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input13_I data_in_a[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07737_ _03190_ _03195_ _03200_ _03205_ _03206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_26_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12110__D _05992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07668_ _02549_ _03138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12455__CLK clknet_leaf_135_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07331__B1 _02648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09407_ _04173_ _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06619_ _02026_ _02010_ _02104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07882__A1 u2.mem\[14\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06685__A2 _02168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07599_ u2.mem\[29\]\[8\] _03068_ _03069_ u2.mem\[11\]\[8\] _03070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07882__B2 u2.mem\[12\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09338_ _04265_ u2.mem\[28\]\[6\] _04341_ _04344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06437__A2 _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09269_ _04274_ u2.mem\[26\]\[10\] _04300_ _04303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11300_ _05567_ _05568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_12280_ _00159_ clknet_leaf_118_clock u2.mem\[9\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11231_ _05514_ u2.mem\[151\]\[4\] _05519_ _05525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10241__I0 _04907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11162_ _05470_ u2.mem\[147\]\[4\] _05474_ _05480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10113_ _04829_ _00745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11093_ _05437_ _01117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08737__I1 u2.mem\[14\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09934__I0 _04685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_351_clock clknet_5_4_0_clock clknet_leaf_351_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_49_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10044_ _04783_ _04784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_49_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11741__I0 _05833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11185__S _05492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11995_ _00007_ clknet_leaf_344_clock u2.mem\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_366_clock clknet_5_4_0_clock clknet_leaf_366_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09162__I1 u2.mem\[24\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12020__D mem_address_trans\[7\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10946_ _05343_ u2.mem\[134\]\[2\] _05337_ _05344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13380__CLK clknet_leaf_367_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10877_ _05299_ u2.mem\[130\]\[1\] _05297_ _05300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_43_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12948__CLK clknet_leaf_64_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12616_ _00495_ clknet_leaf_136_clock u2.mem\[30\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08293__I _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12547_ _00426_ clknet_leaf_110_clock u2.mem\[26\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08673__I0 _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07130__C _02450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06979__A3 _02416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12478_ _00357_ clknet_leaf_196_clock u2.mem\[22\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_304_clock clknet_5_20_0_clock clknet_leaf_304_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10264__S _04923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11429_ _05648_ _01242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11980__I0 _05222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10783__I1 u2.mem\[62\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12328__CLK clknet_leaf_136_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06970_ _02448_ _02449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xclkbuf_leaf_319_clock clknet_5_16_0_clock clknet_leaf_319_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_171_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08728__I1 u2.mem\[14\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input5_I col_select_a[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09925__I0 _04714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08640_ _03895_ _00206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06364__A1 u2.mem\[154\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07372__I _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07561__B1 _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08571_ _03480_ _03605_ _03606_ _03775_ _03855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_82_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11823__S _05887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07522_ _02990_ _02991_ _02992_ _02993_ _02994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_74_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07453_ _02621_ _02927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07864__A1 _03299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06667__A2 _02060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10439__S _05030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06404_ u2.mem\[146\]\[5\] _01691_ _01693_ u2.mem\[186\]\[5\] _01906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06716__I _02137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07384_ u2.mem\[39\]\[4\] _02857_ _02858_ u2.mem\[48\]\[4\] _02859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09123_ _04145_ u2.mem\[23\]\[5\] _04208_ _04210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06335_ _01836_ _01837_ _01838_ _01839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_136_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09054_ data_in_trans\[12\].data_sync _04166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06266_ _01727_ _01554_ _01737_ _01771_ _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08005_ _01591_ _03464_ _03467_ _01678_ _03468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_151_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06197_ _01552_ _01616_ _01704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09963__S _04734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07919__A2 _02493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06451__I _01923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08041__A1 _03499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11971__I0 _05213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13253__CLK clknet_leaf_307_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09956_ _04707_ u2.mem\[42\]\[11\] _04729_ _04733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08579__S _03856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09762__I _04614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08907_ _04041_ u2.mem\[18\]\[12\] _04066_ _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_4105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_24_clock_I clknet_5_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09887_ _04688_ _00660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08838_ _04022_ _00277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10701__I _05173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06355__A1 u2.mem\[175\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06355__B2 u2.mem\[188\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08769_ _03961_ _03977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10800_ _04416_ _05172_ _05252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_148_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11780_ _05867_ _01374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07304__B1 _02612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10731_ _03682_ _05209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06658__A2 _02077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_249_clock_I clknet_5_18_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13450_ _01329_ clknet_leaf_359_clock u2.mem\[178\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10662_ _05166_ _00957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12401_ _00280_ clknet_leaf_172_clock u2.mem\[17\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13381_ _01260_ clknet_leaf_319_clock u2.mem\[167\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_167_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10593_ _05126_ u2.mem\[57\]\[14\] _05122_ _05127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12332_ _00211_ clknet_5_28_0_clock u2.mem\[13\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10462__I0 _05020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06291__B1 _01715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10084__S _04811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12263_ _00142_ clknet_leaf_54_clock u2.mem\[8\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06830__A2 _02192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_301_clock_I clknet_5_21_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11167__A1 _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08958__I1 u2.mem\[20\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11214_ _05513_ _05514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12194_ _00073_ clknet_leaf_252_clock u2.mem\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11962__I0 _05913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_290_clock clknet_5_21_0_clock clknet_leaf_290_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11145_ _05469_ _01137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07791__B1 _03105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12620__CLK clknet_leaf_201_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11076_ _05342_ _05426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09532__A1 _04013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10027_ _04703_ u2.mem\[44\]\[9\] _04772_ _04774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08288__I _03665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06346__A1 u2.mem\[178\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06346__B2 u2.mem\[164\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06897__A2 _02375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11978_ _05220_ u2.mem\[194\]\[11\] _05985_ _05987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_75_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06649__A2 _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10929_ _05331_ _01059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12000__CLK clknet_leaf_19_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13126__CLK clknet_leaf_21_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_243_clock clknet_5_24_0_clock clknet_leaf_243_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10453__I0 _05011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06120_ u2.mem\[184\]\[0\] _01626_ _01553_ _01627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08751__I _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12150__CLK clknet_leaf_74_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06051_ col_select_trans\[2\].data_sync _01558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13276__CLK clknet_leaf_8_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07367__I _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10205__I0 _04815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08023__A1 _03482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11953__I0 _05903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_258_clock clknet_5_19_0_clock clknet_leaf_258_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_113_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09810_ _04576_ u2.mem\[39\]\[3\] _04639_ _04643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_59_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10722__S _05196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07782__B1 _03228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09741_ _04598_ _04599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06953_ _02431_ _02432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11705__I0 _05792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07129__A3 _02602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_198_clock_I clknet_5_31_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09672_ _04476_ u2.mem\[36\]\[5\] _04549_ _04551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06884_ _02362_ _02363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_41_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07534__B1 _02916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08623_ _03810_ u2.mem\[12\]\[5\] _03884_ _03886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11553__S _05721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08554_ _03816_ u2.mem\[10\]\[8\] _03845_ _03846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07505_ u2.mem\[27\]\[7\] _02871_ _02872_ u2.mem\[35\]\[7\] _02977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_78_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08485_ _03800_ _00146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_250_clock_I clknet_5_19_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07436_ u2.mem\[26\]\[5\] _02908_ _02909_ u2.mem\[10\]\[5\] _02910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06446__I _01927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07367_ _02581_ _02842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09106_ _04174_ u2.mem\[22\]\[14\] _04197_ _04200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09757__I data_in_trans\[14\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10444__I0 _05001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06318_ u2.mem\[145\]\[3\] _01640_ _01732_ u2.mem\[168\]\[3\] _01822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_87_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07298_ u2.mem\[17\]\[3\] _02586_ _02591_ u2.mem\[24\]\[3\] _02774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_108_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09037_ data_in_trans\[8\].data_sync _04153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06249_ _01748_ _01751_ _01752_ _01754_ _01755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_117_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12643__CLK clknet_leaf_93_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11944__I0 _05225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07773__B1 _03083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09939_ _04723_ _00677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12950_ _00829_ clknet_leaf_63_clock u2.mem\[51\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12793__CLK clknet_leaf_340_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06328__A1 u2.mem\[152\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11901_ u2.mem\[192\]\[10\] _03522_ _05942_ _05943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12881_ _00760_ clknet_leaf_245_clock u2.mem\[47\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11832_ _05899_ _01394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08836__I _03670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12023__CLK clknet_2_2__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13149__CLK clknet_leaf_277_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08876__I0 _04048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11763_ _05856_ _05857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_26_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13502_ _01381_ clknet_leaf_345_clock u2.mem\[187\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10714_ _05197_ _00978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08772__S _03977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11694_ _05814_ _01341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13433_ _01312_ clknet_leaf_352_clock u2.mem\[175\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12173__CLK clknet_leaf_231_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13299__CLK clknet_leaf_382_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10645_ _05151_ _05157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_158_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10435__I0 _04987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13364_ _01243_ clknet_leaf_363_clock u2.mem\[164\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10576_ _03695_ _05115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12315_ _00194_ clknet_leaf_185_clock u2.mem\[12\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13295_ _01174_ clknet_leaf_0_clock u2.mem\[152\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12246_ _00125_ clknet_leaf_73_clock u2.mem\[7\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08005__A1 _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08005__B2 _01678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11935__I0 _05216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11638__S _05779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08800__I0 _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12177_ _00056_ clknet_leaf_233_clock u2.mem\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_150_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07764__B1 _03138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09108__S _04197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11128_ _05430_ u2.mem\[145\]\[4\] _05452_ _05458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11059_ _05415_ _01105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06319__B2 u2.mem\[188\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11373__S _05607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08867__I0 _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12516__CLK clknet_leaf_107_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09778__S _04623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08270_ _03577_ u2.mem\[4\]\[14\] _03649_ _03652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07295__A2 _02580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07221_ _01726_ _02361_ _02665_ _02698_ _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_182_clock clknet_5_27_0_clock clknet_leaf_182_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_20_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11900__I _05927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08481__I _03655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07047__A2 _02521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07152_ _02613_ _02620_ _02625_ _02630_ _02631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_34_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09292__I0 _04258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12666__CLK clknet_leaf_60_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06103_ _01607_ _01609_ _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06255__B1 _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07083_ _02363_ _02562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_173_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_197_clock clknet_5_31_0_clock clknet_leaf_197_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_12_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06034_ inverter_select_trans.data_sync _01542_ _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09044__I0 _04158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11926__I0 _05915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10729__I1 u2.mem\[61\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07755__B1 _03123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07825__I _02541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_120_clock clknet_5_14_0_clock clknet_leaf_120_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07985_ u2.mem\[52\]\[15\] _03315_ _03316_ u2.mem\[21\]\[15\] _03449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09724_ _04585_ _04586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06936_ _02414_ _02350_ _02415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08857__S _04033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12046__CLK clknet_leaf_315_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11154__I1 u2.mem\[147\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09655_ _04540_ _00576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06867_ _02338_ _02345_ _02346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_28_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08606_ _03832_ u2.mem\[11\]\[15\] _03871_ _03875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_135_clock clknet_5_15_0_clock clknet_leaf_135_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_43_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08656__I _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09586_ _04463_ u2.mem\[34\]\[0\] _04501_ _04502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07560__I _02460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06798_ u2.mem\[167\]\[4\] _02058_ _02061_ u2.mem\[183\]\[4\] _02279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06730__A1 u2.mem\[180\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08537_ _03836_ _00162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12196__CLK clknet_leaf_22_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11606__A2 _05729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11082__I _05348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13441__CLK clknet_leaf_363_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08468_ _03701_ u2.mem\[8\]\[10\] _03787_ _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07419_ _02524_ _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_168_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08399_ _03542_ _03481_ _03747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__10627__S _05146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11810__I _05768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10430_ _03720_ _05027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06246__B1 _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11090__I0 _05420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10361_ _04909_ u2.mem\[52\]\[10\] _04976_ _04979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_128_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06797__A1 u2.mem\[164\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07994__B1 _03436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12100_ _01498_ clknet_leaf_246_clock u2.active_mem\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06797__B2 u2.mem\[178\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09035__I0 _04151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13080_ _00959_ clknet_leaf_341_clock u2.mem\[59\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10292_ _04939_ _00814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11917__I0 _05907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12031_ net40 clknet_2_3__leaf_clock_a row_select_trans\[3\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06549__A1 _02031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07746__B1 _03034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08767__S _03972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12933_ _00812_ clknet_leaf_63_clock u2.mem\[50\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12539__CLK clknet_leaf_187_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12864_ _00743_ clknet_leaf_154_clock u2.mem\[46\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06721__A1 _01727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11815_ _05868_ u2.mem\[188\]\[1\] _05888_ _05890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12795_ _00674_ clknet_leaf_184_clock u2.mem\[42\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11921__S _05950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07277__A2 _02650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11746_ _05846_ _01361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_146_clock_I clknet_5_13_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11677_ _05804_ _01334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09397__I _04163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13416_ _01295_ clknet_leaf_324_clock u2.mem\[172\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10628_ _05147_ _00942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09274__I0 _04278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10336__I _04862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13347_ _01226_ clknet_leaf_14_clock u2.mem\[161\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10559_ _05000_ _05103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13278_ _01157_ clknet_leaf_8_clock u2.mem\[149\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12229_ _00108_ clknet_leaf_73_clock u2.mem\[6\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12069__CLK clknet_2_1__leaf_clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13314__CLK clknet_5_5_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07201__A2 _02572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07770_ _03234_ _03235_ _03236_ _03237_ _03238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_110_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_52_clock clknet_5_13_0_clock clknet_leaf_52_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_133_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06721_ _01727_ _01995_ _02171_ _02204_ _01475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_49_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09440_ _04409_ _00492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13464__CLK clknet_leaf_360_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06652_ _02056_ _02001_ _02137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10895__I0 _05299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09371_ _04135_ _04364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06583_ _02067_ _02068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_67_clock clknet_5_9_0_clock clknet_leaf_67_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11831__S _05896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08322_ _03692_ u2.mem\[5\]\[8\] _03693_ _03694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07268__A2 _02638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09301__S _04318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08253_ _03642_ _00072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07204_ _02593_ _02682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_159_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09265__I0 _04269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08184_ _03584_ _03600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_20_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10246__I _04601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07135_ _02478_ _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_14_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06779__A1 u2.mem\[180\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06779__B2 u2.mem\[172\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07976__B1 _02550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07066_ u2.mem\[60\]\[0\] _02542_ _02544_ u2.mem\[62\]\[0\] _02545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_133_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06017_ u2.driver_mem\[4\] _01522_ _01525_ _01519_ _01526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA_clkbuf_leaf_348_clock_I clknet_5_7_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07728__B1 _03080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11524__A1 _04287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09971__S _04740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06400__B1 _01672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07968_ u2.mem\[14\]\[15\] _02521_ _02525_ u2.mem\[12\]\[15\] _03432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10910__S _05319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06951__A1 _02428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06919_ u2.mem\[32\]\[0\] _02385_ _02397_ u2.mem\[2\]\[0\] _02398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09707_ _04572_ _04573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07899_ u2.mem\[52\]\[13\] _03315_ _03316_ u2.mem\[21\]\[13\] _03365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_90_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10886__I0 _05305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09638_ _04480_ u2.mem\[35\]\[7\] _04527_ _04531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09569_ _04489_ u2.mem\[33\]\[11\] _04483_ _04490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11741__S _05840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11600_ _05676_ _05756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12580_ _00459_ clknet_leaf_96_clock u2.mem\[28\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11531_ _05670_ _05713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10357__S _04976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12981__CLK clknet_leaf_30_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11462_ _05668_ u2.mem\[166\]\[1\] _05665_ _05669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09256__I0 _04260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09010__I _04131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13201_ _01080_ clknet_leaf_295_clock u2.mem\[137\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10413_ _05015_ _00859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11393_ _05624_ _05625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_124_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07967__B1 _02518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13132_ _01011_ clknet_leaf_262_clock u2.mem\[63\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10344_ _04969_ _00836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13337__CLK clknet_leaf_4_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13063_ _00942_ clknet_leaf_47_clock u2.mem\[58\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07982__A3 _03444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10275_ _04898_ u2.mem\[50\]\[5\] _04928_ _04930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07719__B1 _03063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12014_ mem_address_trans\[4\].A clknet_leaf_315_clock mem_address_trans\[4\].data_sync
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12361__CLK clknet_leaf_136_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13487__CLK clknet_leaf_314_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10820__S _05263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08497__S _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_72_clock_I clknet_5_8_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10877__I0 _05299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12916_ _00795_ clknet_leaf_87_clock u2.mem\[49\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07498__A2 _02927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12847_ _00726_ clknet_leaf_155_clock u2.mem\[45\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10629__I0 _05124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12778_ _00657_ clknet_leaf_141_clock u2.mem\[40\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09121__S _04208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06972__C _02450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_297_clock_I clknet_5_21_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11729_ _05836_ _01354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09247__I0 _04246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08960__S _04097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11098__S _05434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08940_ _04086_ _00315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07375__I _02600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09791__S _04628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11357__I1 u2.mem\[159\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08871_ _04045_ _00287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07822_ _03281_ _03282_ _03285_ _03288_ _03289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_57_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07753_ u2.mem\[58\]\[11\] _03044_ _03045_ u2.mem\[36\]\[11\] _03221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_42_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06704_ u2.mem\[188\]\[1\] _02185_ _02186_ u2.mem\[187\]\[1\] _02187_ u2.mem\[192\]\[1\]
+ _02188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_168_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10868__I0 _05207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07684_ _03150_ _03151_ _03152_ _03153_ _03154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__07489__A2 _02959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09423_ _04364_ u2.mem\[30\]\[3\] _04396_ _04400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_77_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06697__B1 _02061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06635_ _02119_ _02015_ _02120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_168_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06161__A2 _01664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09354_ _04281_ u2.mem\[28\]\[13\] _04351_ _04353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06566_ _02050_ _02051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09031__S _04141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08305_ _03679_ _03680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09285_ _04312_ _04313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_138_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06497_ u2.mem\[193\]\[15\] _01917_ _01982_ _01911_ _01983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_166_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08236_ _03631_ _03632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09238__I0 _04283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06454__I _01913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07661__A2 _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11045__I0 _05386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08167_ _03554_ u2.mem\[2\]\[4\] _03590_ _03591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07118_ u2.mem\[23\]\[0\] _02594_ _02596_ u2.mem\[22\]\[0\] _02597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_162_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08098_ mem_address_trans\[1\].data_sync _03542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08610__A1 _03629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12384__CLK clknet_leaf_234_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06621__B1 _02105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07049_ _02527_ _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10060_ _04582_ _04795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07177__A1 _02649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07716__A3 _03179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10962_ _05355_ _05356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_56_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09005__I _04127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12701_ _00580_ clknet_leaf_222_clock u2.mem\[36\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06688__B1 _02087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06688__C2 _02089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10893_ _05294_ u2.mem\[131\]\[0\] _05310_ _05311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12632_ _00511_ clknet_leaf_112_clock u2.mem\[31\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12563_ _00442_ clknet_leaf_112_clock u2.mem\[27\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10087__S _04811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11514_ _05702_ _01273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_19_clock_I clknet_5_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12494_ _00373_ clknet_leaf_197_clock u2.mem\[23\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11036__I0 _05392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12018__D mem_address_trans\[6\].A vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11445_ _05657_ _01249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12727__CLK clknet_leaf_45_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11376_ _05614_ _01223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10327_ _04943_ _04959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_13115_ _00994_ clknet_leaf_261_clock u2.mem\[62\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11339__I1 u2.mem\[158\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13046_ _00925_ clknet_leaf_33_clock u2.mem\[57\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10258_ _04919_ _00800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12877__CLK clknet_leaf_224_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11646__S _05778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10189_ _04799_ u2.mem\[48\]\[7\] _04870_ _04874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09116__S _04203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12107__CLK clknet_leaf_47_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06391__A2 _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06539__I row_select_trans\[1\].data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06420_ u2.mem\[193\]\[0\] _01917_ _01919_ u2.mem\[192\]\[0\] _01920_ _01921_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_37_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06351_ u2.mem\[145\]\[4\] _01639_ _01642_ u2.mem\[163\]\[4\] u2.mem\[165\]\[4\]
+ _01646_ _01854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_37_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09070_ _04178_ _00353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06282_ u2.mem\[159\]\[2\] _01604_ _01595_ u2.mem\[149\]\[2\] _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_120_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08021_ mem_address_trans\[2\].data_sync mem_address_trans\[3\].data_sync _03482_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_50_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06851__B1 _02147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09585__I _04500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11578__I1 u2.mem\[173\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09972_ _04742_ _00691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08923_ _04019_ u2.mem\[19\]\[2\] _04074_ _04077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07159__B2 u2.mem\[30\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08854_ _04032_ u2.mem\[17\]\[8\] _04033_ _04034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11750__I1 u2.mem\[184\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07805_ u2.mem\[50\]\[12\] _03113_ _03114_ u2.mem\[51\]\[12\] _03272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_79_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08785_ _03982_ _03988_ _03989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05997_ u2.select_mem_row\[0\] row_col_select_trans.data_sync _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07736_ _03201_ _03202_ _03203_ _03204_ _03205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_84_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07667_ _02547_ _03137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_168_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06893__B _02353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09406_ _04388_ _00479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06618_ _02014_ _02011_ _02103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07598_ _02563_ _03069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07882__A2 _02521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09337_ _04343_ _00455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06549_ _02031_ _02033_ _02034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_20_clock_I clknet_5_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09268_ _04302_ _00427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08219_ _03568_ u2.mem\[3\]\[10\] _03618_ _03621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09199_ _04256_ u2.mem\[25\]\[2\] _04252_ _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09495__I _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11230_ _05524_ _01167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11161_ _05479_ _01143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10434__I _05029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10112_ _04799_ u2.mem\[46\]\[7\] _04825_ _04829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06070__A1 _01552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_245_clock_I clknet_5_24_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11092_ _05424_ u2.mem\[143\]\[1\] _05435_ _05437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_1_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10043_ _03903_ _04760_ _04783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08839__I _03674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11741__I1 u2.mem\[183\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08362__A3 _03632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06373__A2 _01853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11994_ _00006_ clknet_leaf_334_clock u2.mem\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13525__CLK clknet_leaf_329_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10945_ _05342_ _05343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08370__I0 _03671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10876_ _04991_ _05299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12615_ _00494_ clknet_leaf_137_clock u2.mem\[30\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08122__I0 _03559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07086__B1 _02564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12546_ _00425_ clknet_leaf_189_clock u2.mem\[26\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07625__A2 _02927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12477_ _00356_ clknet_leaf_196_clock u2.mem\[22\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11428_ _05623_ u2.mem\[164\]\[0\] _05647_ _05648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11359_ _05595_ u2.mem\[159\]\[5\] _05597_ _05604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08189__I0 _03577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13029_ _00908_ clknet_leaf_29_clock u2.mem\[56\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07653__I _02517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06364__A2 _01699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08570_ _03854_ _00177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06269__I _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07521_ u2.mem\[43\]\[7\] _02820_ _02821_ u2.mem\[20\]\[7\] _02993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_81_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07313__A1 u2.mem\[32\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07452_ u2.mem\[8\]\[5\] _02860_ _02861_ u2.mem\[4\]\[5\] _02926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_39_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07864__A2 _03310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06403_ u2.mem\[191\]\[5\] _01681_ _01683_ u2.mem\[179\]\[5\] _01905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_167_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11248__I0 _05517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07383_ _02618_ _02858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09122_ _04209_ _00374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06334_ u2.mem\[146\]\[3\] _01692_ _01694_ u2.mem\[186\]\[3\] _01838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07077__B1 _02555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_194_clock_I clknet_5_31_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09053_ _04165_ _00349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10455__S _05040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06265_ _01745_ _01755_ _01762_ _01770_ _01771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_129_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08004_ _03465_ _03466_ _03467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07828__I _02536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09613__I0 _04491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06196_ _01702_ _01703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11971__I1 u2.mem\[194\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09955_ _04732_ _00684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11286__S _05559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08906_ _04050_ _04066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_98_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08659__I _03666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09886_ _04687_ u2.mem\[41\]\[2\] _04683_ _04688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_4117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07563__I _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13548__CLK clknet_leaf_37_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08837_ _04021_ u2.mem\[17\]\[3\] _04015_ _04022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11085__I _05351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06355__A2 _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08595__S _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08768_ _03976_ _00253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07719_ u2.mem\[37\]\[10\] _03062_ _03063_ u2.mem\[59\]\[10\] _03188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_122_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12572__CLK clknet_leaf_201_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08699_ _03936_ u2.mem\[13\]\[14\] _03932_ _03937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10730_ _05208_ _00983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07855__A2 _03155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10661_ _05119_ u2.mem\[59\]\[11\] _05162_ _05166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12400_ _00279_ clknet_leaf_172_clock u2.mem\[17\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13380_ _01259_ clknet_leaf_367_clock u2.mem\[166\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07607__A2 _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10592_ _03716_ _05126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12331_ _00210_ clknet_leaf_234_clock u2.mem\[13\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06291__A1 u2.mem\[152\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12262_ _00141_ clknet_leaf_72_clock u2.mem\[8\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09604__I0 _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11213_ _03505_ _05513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13078__CLK clknet_leaf_22_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12193_ _00072_ clknet_leaf_253_clock u2.mem\[4\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07240__B1 _02508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11144_ _05468_ u2.mem\[146\]\[3\] _05462_ _05469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11962__I1 u2.mem\[194\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07791__A1 u2.mem\[27\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11075_ _05425_ _01111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10026_ _04773_ _00714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08591__I0 _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11924__S _05955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12915__CLK clknet_leaf_87_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06089__I _01587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11478__I0 _05680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11977_ _05986_ _01452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08343__I0 _03709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10928_ _05303_ u2.mem\[133\]\[3\] _05327_ _05331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_0_clock_a_I clock_a vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10859_ _05288_ _01032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13578_ _01457_ clknet_leaf_35_clock u2.mem\[194\]\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12529_ _00408_ clknet_leaf_178_clock u2.mem\[25\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10275__S _04928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06050_ _01556_ _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06282__A1 u2.mem\[159\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06282__B2 u2.mem\[149\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08023__A2 _03483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06034__A1 inverter_select_trans.data_sync vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12445__CLK clknet_leaf_187_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11953__I1 u2.mem\[194\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07782__A1 _01966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06952_ _02363_ _02370_ _02374_ _02430_ _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_09740_ data_in_trans\[10\].data_sync _04598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
.ends


* NGSPICE file created from clock_mux.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_1 I Z VDD VSS
.ends

.subckt clock_mux clock_out_a clock_out_b clock_out_c core_clock io_clock la_oenb
+ vdd vss
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_1_0__f_net2_I clknet_0_net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output2_I clknet_1_0__leaf_net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_0_core_clock core_clock clknet_0_core_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_37_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_0_net2 net2 clknet_0_net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_23_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input1_I la_oenb vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_1_1__f_core_clock clknet_0_core_clock clknet_1_1__leaf_core_clock vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_11_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_7_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5__I clknet_1_1__leaf_net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_1_1__f_net2 clknet_0_net2 clknet_1_1__leaf_net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput1 la_oenb net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3__D net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5_ clknet_1_1__leaf_net2 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4_ clknet_1_0__leaf_net2 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3_ net1 clknet_1_1__leaf_core_clock sel_reg vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1__I1 io_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2_ _0_ net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_1_0__f_core_clock clknet_0_core_clock clknet_1_0__leaf_core_clock vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_45_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1_ clknet_1_0__leaf_core_clock io_clock sel_reg _0_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_1_0__f_net2 clknet_0_net2 clknet_1_0__leaf_net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_43_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_46_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_37_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_0_core_clock_I core_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_1_1__f_net2_I clknet_0_net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput2 clknet_1_0__leaf_net2 clock_out_a vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput3 net3 clock_out_b vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4__I clknet_1_0__leaf_net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput4 net4 clock_out_c vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_45_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output4_I net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
.ends


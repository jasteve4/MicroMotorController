magic
tech gf180mcuC
magscale 1 5
timestamp 1670292224
<< obsm1 >>
rect 672 1538 24304 23158
<< metal2 >>
rect 1456 0 1512 400
rect 4200 0 4256 400
rect 6944 0 7000 400
rect 9688 0 9744 400
rect 12432 0 12488 400
rect 15176 0 15232 400
rect 17920 0 17976 400
rect 20664 0 20720 400
rect 23408 0 23464 400
<< obsm2 >>
rect 910 430 24066 24127
rect 910 400 1426 430
rect 1542 400 4170 430
rect 4286 400 6914 430
rect 7030 400 9658 430
rect 9774 400 12402 430
rect 12518 400 15146 430
rect 15262 400 17890 430
rect 18006 400 20634 430
rect 20750 400 23378 430
rect 23494 400 24066 430
<< metal3 >>
rect 24600 24080 25000 24136
rect 24600 23352 25000 23408
rect 0 23240 400 23296
rect 24600 22624 25000 22680
rect 24600 21896 25000 21952
rect 24600 21168 25000 21224
rect 24600 20440 25000 20496
rect 0 20160 400 20216
rect 24600 19712 25000 19768
rect 24600 18984 25000 19040
rect 24600 18256 25000 18312
rect 24600 17528 25000 17584
rect 0 17080 400 17136
rect 24600 16800 25000 16856
rect 24600 16072 25000 16128
rect 24600 15344 25000 15400
rect 24600 14616 25000 14672
rect 0 14000 400 14056
rect 24600 13888 25000 13944
rect 24600 13160 25000 13216
rect 24600 12432 25000 12488
rect 24600 11704 25000 11760
rect 0 10920 400 10976
rect 24600 10976 25000 11032
rect 24600 10248 25000 10304
rect 24600 9520 25000 9576
rect 24600 8792 25000 8848
rect 24600 8064 25000 8120
rect 0 7840 400 7896
rect 24600 7336 25000 7392
rect 24600 6608 25000 6664
rect 24600 5880 25000 5936
rect 24600 5152 25000 5208
rect 0 4760 400 4816
rect 24600 4424 25000 4480
rect 24600 3696 25000 3752
rect 24600 2968 25000 3024
rect 24600 2240 25000 2296
rect 0 1680 400 1736
rect 24600 1512 25000 1568
rect 24600 784 25000 840
<< obsm3 >>
rect 400 24050 24570 24122
rect 400 23438 24682 24050
rect 400 23326 24570 23438
rect 430 23322 24570 23326
rect 430 23210 24682 23322
rect 400 22710 24682 23210
rect 400 22594 24570 22710
rect 400 21982 24682 22594
rect 400 21866 24570 21982
rect 400 21254 24682 21866
rect 400 21138 24570 21254
rect 400 20526 24682 21138
rect 400 20410 24570 20526
rect 400 20246 24682 20410
rect 430 20130 24682 20246
rect 400 19798 24682 20130
rect 400 19682 24570 19798
rect 400 19070 24682 19682
rect 400 18954 24570 19070
rect 400 18342 24682 18954
rect 400 18226 24570 18342
rect 400 17614 24682 18226
rect 400 17498 24570 17614
rect 400 17166 24682 17498
rect 430 17050 24682 17166
rect 400 16886 24682 17050
rect 400 16770 24570 16886
rect 400 16158 24682 16770
rect 400 16042 24570 16158
rect 400 15430 24682 16042
rect 400 15314 24570 15430
rect 400 14702 24682 15314
rect 400 14586 24570 14702
rect 400 14086 24682 14586
rect 430 13974 24682 14086
rect 430 13970 24570 13974
rect 400 13858 24570 13970
rect 400 13246 24682 13858
rect 400 13130 24570 13246
rect 400 12518 24682 13130
rect 400 12402 24570 12518
rect 400 11790 24682 12402
rect 400 11674 24570 11790
rect 400 11062 24682 11674
rect 400 11006 24570 11062
rect 430 10946 24570 11006
rect 430 10890 24682 10946
rect 400 10334 24682 10890
rect 400 10218 24570 10334
rect 400 9606 24682 10218
rect 400 9490 24570 9606
rect 400 8878 24682 9490
rect 400 8762 24570 8878
rect 400 8150 24682 8762
rect 400 8034 24570 8150
rect 400 7926 24682 8034
rect 430 7810 24682 7926
rect 400 7422 24682 7810
rect 400 7306 24570 7422
rect 400 6694 24682 7306
rect 400 6578 24570 6694
rect 400 5966 24682 6578
rect 400 5850 24570 5966
rect 400 5238 24682 5850
rect 400 5122 24570 5238
rect 400 4846 24682 5122
rect 430 4730 24682 4846
rect 400 4510 24682 4730
rect 400 4394 24570 4510
rect 400 3782 24682 4394
rect 400 3666 24570 3782
rect 400 3054 24682 3666
rect 400 2938 24570 3054
rect 400 2326 24682 2938
rect 400 2210 24570 2326
rect 400 1766 24682 2210
rect 430 1650 24682 1766
rect 400 1598 24682 1650
rect 400 1482 24570 1598
rect 400 870 24682 1482
rect 400 798 24570 870
<< metal4 >>
rect 2224 1538 2384 23158
rect 9904 1538 10064 23158
rect 17584 1538 17744 23158
<< labels >>
rlabel metal2 s 1456 0 1512 400 6 clock
port 1 nsew signal input
rlabel metal3 s 24600 784 25000 840 6 clock_out
port 2 nsew signal output
rlabel metal3 s 24600 1512 25000 1568 6 data_out[0]
port 3 nsew signal output
rlabel metal3 s 24600 8792 25000 8848 6 data_out[10]
port 4 nsew signal output
rlabel metal3 s 24600 9520 25000 9576 6 data_out[11]
port 5 nsew signal output
rlabel metal3 s 24600 10248 25000 10304 6 data_out[12]
port 6 nsew signal output
rlabel metal3 s 24600 10976 25000 11032 6 data_out[13]
port 7 nsew signal output
rlabel metal3 s 24600 11704 25000 11760 6 data_out[14]
port 8 nsew signal output
rlabel metal3 s 24600 12432 25000 12488 6 data_out[15]
port 9 nsew signal output
rlabel metal3 s 24600 13160 25000 13216 6 data_out[16]
port 10 nsew signal output
rlabel metal3 s 24600 13888 25000 13944 6 data_out[17]
port 11 nsew signal output
rlabel metal3 s 24600 14616 25000 14672 6 data_out[18]
port 12 nsew signal output
rlabel metal3 s 24600 15344 25000 15400 6 data_out[19]
port 13 nsew signal output
rlabel metal3 s 24600 2240 25000 2296 6 data_out[1]
port 14 nsew signal output
rlabel metal3 s 24600 16072 25000 16128 6 data_out[20]
port 15 nsew signal output
rlabel metal3 s 24600 16800 25000 16856 6 data_out[21]
port 16 nsew signal output
rlabel metal3 s 24600 17528 25000 17584 6 data_out[22]
port 17 nsew signal output
rlabel metal3 s 24600 18256 25000 18312 6 data_out[23]
port 18 nsew signal output
rlabel metal3 s 24600 18984 25000 19040 6 data_out[24]
port 19 nsew signal output
rlabel metal3 s 24600 19712 25000 19768 6 data_out[25]
port 20 nsew signal output
rlabel metal3 s 24600 20440 25000 20496 6 data_out[26]
port 21 nsew signal output
rlabel metal3 s 24600 21168 25000 21224 6 data_out[27]
port 22 nsew signal output
rlabel metal3 s 24600 21896 25000 21952 6 data_out[28]
port 23 nsew signal output
rlabel metal3 s 24600 22624 25000 22680 6 data_out[29]
port 24 nsew signal output
rlabel metal3 s 24600 2968 25000 3024 6 data_out[2]
port 25 nsew signal output
rlabel metal3 s 24600 23352 25000 23408 6 data_out[30]
port 26 nsew signal output
rlabel metal3 s 24600 24080 25000 24136 6 data_out[31]
port 27 nsew signal output
rlabel metal3 s 24600 3696 25000 3752 6 data_out[3]
port 28 nsew signal output
rlabel metal3 s 24600 4424 25000 4480 6 data_out[4]
port 29 nsew signal output
rlabel metal3 s 24600 5152 25000 5208 6 data_out[5]
port 30 nsew signal output
rlabel metal3 s 24600 5880 25000 5936 6 data_out[6]
port 31 nsew signal output
rlabel metal3 s 24600 6608 25000 6664 6 data_out[7]
port 32 nsew signal output
rlabel metal3 s 24600 7336 25000 7392 6 data_out[8]
port 33 nsew signal output
rlabel metal3 s 24600 8064 25000 8120 6 data_out[9]
port 34 nsew signal output
rlabel metal2 s 15176 0 15232 400 6 la_data_in[0]
port 35 nsew signal input
rlabel metal2 s 17920 0 17976 400 6 la_data_in[1]
port 36 nsew signal input
rlabel metal2 s 20664 0 20720 400 6 la_data_in[2]
port 37 nsew signal input
rlabel metal2 s 23408 0 23464 400 6 la_data_in[3]
port 38 nsew signal input
rlabel metal2 s 4200 0 4256 400 6 la_oenb[0]
port 39 nsew signal output
rlabel metal2 s 6944 0 7000 400 6 la_oenb[1]
port 40 nsew signal output
rlabel metal2 s 9688 0 9744 400 6 la_oenb[2]
port 41 nsew signal output
rlabel metal2 s 12432 0 12488 400 6 la_oenb[3]
port 42 nsew signal output
rlabel metal3 s 0 20160 400 20216 6 miso
port 43 nsew signal output
rlabel metal3 s 0 23240 400 23296 6 miso_oeb
port 44 nsew signal output
rlabel metal3 s 0 7840 400 7896 6 mosi
port 45 nsew signal input
rlabel metal3 s 0 10920 400 10976 6 mosi_oeb
port 46 nsew signal output
rlabel metal3 s 0 1680 400 1736 6 sclk
port 47 nsew signal input
rlabel metal3 s 0 4760 400 4816 6 sclk_oeb
port 48 nsew signal output
rlabel metal3 s 0 14000 400 14056 6 ss_n
port 49 nsew signal input
rlabel metal3 s 0 17080 400 17136 6 ss_n_oeb
port 50 nsew signal output
rlabel metal4 s 2224 1538 2384 23158 6 vdd
port 51 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 23158 6 vdd
port 51 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 23158 6 vss
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 25000 25000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 525346
string GDS_FILE /home/jasteve4/Documents/MicroMotorController/openlane/spi_core/runs/22_12_05_21_02/results/signoff/spi_core.magic.gds
string GDS_START 100860
<< end >>


magic
tech gf180mcuC
magscale 1 10
timestamp 1670292224
<< metal1 >>
rect 1344 46282 48608 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 48608 46282
rect 1344 46196 48608 46230
rect 1822 46114 1874 46126
rect 1822 46050 1874 46062
rect 47842 45950 47854 46002
rect 47906 45950 47918 46002
rect 44930 45838 44942 45890
rect 44994 45838 45006 45890
rect 46722 45838 46734 45890
rect 46786 45838 46798 45890
rect 46050 45726 46062 45778
rect 46114 45726 46126 45778
rect 44158 45666 44210 45678
rect 44158 45602 44210 45614
rect 1344 45498 48608 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 48608 45498
rect 1344 45412 48608 45446
rect 44930 45054 44942 45106
rect 44994 45054 45006 45106
rect 44494 44994 44546 45006
rect 46622 44994 46674 45006
rect 45938 44942 45950 44994
rect 46002 44942 46014 44994
rect 44494 44930 44546 44942
rect 46622 44930 46674 44942
rect 1344 44714 48608 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 48608 44714
rect 1344 44628 48608 44662
rect 44718 44322 44770 44334
rect 45490 44270 45502 44322
rect 45554 44270 45566 44322
rect 44718 44258 44770 44270
rect 46610 44158 46622 44210
rect 46674 44158 46686 44210
rect 1344 43930 48608 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 48608 43930
rect 1344 43844 48608 43878
rect 1344 43146 48608 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 48608 43146
rect 1344 43060 48608 43094
rect 45490 42702 45502 42754
rect 45554 42702 45566 42754
rect 46610 42590 46622 42642
rect 46674 42590 46686 42642
rect 44718 42530 44770 42542
rect 44718 42466 44770 42478
rect 1344 42362 48608 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 48608 42362
rect 1344 42276 48608 42310
rect 1344 41578 48608 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 48608 41578
rect 1344 41492 48608 41526
rect 44718 41186 44770 41198
rect 3042 41134 3054 41186
rect 3106 41134 3118 41186
rect 45490 41134 45502 41186
rect 45554 41134 45566 41186
rect 44718 41122 44770 41134
rect 1922 41022 1934 41074
rect 1986 41022 1998 41074
rect 46610 41022 46622 41074
rect 46674 41022 46686 41074
rect 1344 40794 48608 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 48608 40794
rect 1344 40708 48608 40742
rect 3278 40626 3330 40638
rect 3278 40562 3330 40574
rect 3614 40402 3666 40414
rect 3614 40338 3666 40350
rect 4062 40402 4114 40414
rect 4062 40338 4114 40350
rect 1344 40010 48608 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 48608 40010
rect 1344 39924 48608 39958
rect 45490 39566 45502 39618
rect 45554 39566 45566 39618
rect 46610 39454 46622 39506
rect 46674 39454 46686 39506
rect 44718 39394 44770 39406
rect 44718 39330 44770 39342
rect 1344 39226 48608 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 48608 39226
rect 1344 39140 48608 39174
rect 44930 38782 44942 38834
rect 44994 38782 45006 38834
rect 46050 38670 46062 38722
rect 46114 38670 46126 38722
rect 1344 38442 48608 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 48608 38442
rect 1344 38356 48608 38390
rect 45714 37998 45726 38050
rect 45778 37998 45790 38050
rect 46610 37886 46622 37938
rect 46674 37886 46686 37938
rect 47182 37826 47234 37838
rect 47182 37762 47234 37774
rect 1344 37658 48608 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 48608 37658
rect 1344 37572 48608 37606
rect 39454 37490 39506 37502
rect 39454 37426 39506 37438
rect 39902 37490 39954 37502
rect 39902 37426 39954 37438
rect 43374 37490 43426 37502
rect 43374 37426 43426 37438
rect 42354 37326 42366 37378
rect 42418 37326 42430 37378
rect 42802 37326 42814 37378
rect 42866 37326 42878 37378
rect 42030 37266 42082 37278
rect 46162 37214 46174 37266
rect 46226 37214 46238 37266
rect 42030 37202 42082 37214
rect 45266 37102 45278 37154
rect 45330 37102 45342 37154
rect 41694 37042 41746 37054
rect 41694 36978 41746 36990
rect 1344 36874 48608 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 48608 36874
rect 1344 36788 48608 36822
rect 38334 36706 38386 36718
rect 38334 36642 38386 36654
rect 40238 36706 40290 36718
rect 40238 36642 40290 36654
rect 42142 36706 42194 36718
rect 42142 36642 42194 36654
rect 35646 36594 35698 36606
rect 35646 36530 35698 36542
rect 36878 36594 36930 36606
rect 36878 36530 36930 36542
rect 43486 36482 43538 36494
rect 46734 36482 46786 36494
rect 44482 36430 44494 36482
rect 44546 36430 44558 36482
rect 43486 36418 43538 36430
rect 46734 36418 46786 36430
rect 47630 36370 47682 36382
rect 38658 36318 38670 36370
rect 38722 36318 38734 36370
rect 39106 36318 39118 36370
rect 39170 36318 39182 36370
rect 40450 36318 40462 36370
rect 40514 36318 40526 36370
rect 41010 36318 41022 36370
rect 41074 36318 41086 36370
rect 42354 36318 42366 36370
rect 42418 36318 42430 36370
rect 42914 36318 42926 36370
rect 42978 36318 42990 36370
rect 46162 36318 46174 36370
rect 46226 36318 46238 36370
rect 46498 36318 46510 36370
rect 46562 36318 46574 36370
rect 47630 36306 47682 36318
rect 35198 36258 35250 36270
rect 35198 36194 35250 36206
rect 36206 36258 36258 36270
rect 36206 36194 36258 36206
rect 37998 36258 38050 36270
rect 37998 36194 38050 36206
rect 39902 36258 39954 36270
rect 39902 36194 39954 36206
rect 41806 36258 41858 36270
rect 41806 36194 41858 36206
rect 44718 36258 44770 36270
rect 44718 36194 44770 36206
rect 47070 36258 47122 36270
rect 47070 36194 47122 36206
rect 48078 36258 48130 36270
rect 48078 36194 48130 36206
rect 1344 36090 48608 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 48608 36090
rect 1344 36004 48608 36038
rect 42366 35922 42418 35934
rect 42366 35858 42418 35870
rect 40126 35810 40178 35822
rect 34290 35758 34302 35810
rect 34354 35758 34366 35810
rect 34850 35758 34862 35810
rect 34914 35758 34926 35810
rect 40126 35746 40178 35758
rect 40462 35810 40514 35822
rect 40462 35746 40514 35758
rect 41918 35810 41970 35822
rect 47742 35810 47794 35822
rect 45042 35758 45054 35810
rect 45106 35758 45118 35810
rect 41918 35746 41970 35758
rect 47742 35746 47794 35758
rect 35970 35646 35982 35698
rect 36034 35646 36046 35698
rect 41682 35646 41694 35698
rect 41746 35646 41758 35698
rect 44258 35646 44270 35698
rect 44322 35646 44334 35698
rect 47954 35646 47966 35698
rect 48018 35646 48030 35698
rect 32734 35586 32786 35598
rect 39230 35586 39282 35598
rect 36642 35534 36654 35586
rect 36706 35534 36718 35586
rect 38770 35534 38782 35586
rect 38834 35534 38846 35586
rect 32734 35522 32786 35534
rect 39230 35522 39282 35534
rect 43822 35586 43874 35598
rect 47170 35534 47182 35586
rect 47234 35534 47246 35586
rect 43822 35522 43874 35534
rect 33742 35474 33794 35486
rect 33742 35410 33794 35422
rect 34078 35474 34130 35486
rect 34078 35410 34130 35422
rect 1344 35306 48608 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 48608 35306
rect 1344 35220 48608 35254
rect 45950 35138 46002 35150
rect 45950 35074 46002 35086
rect 46286 35138 46338 35150
rect 46286 35074 46338 35086
rect 34862 35026 34914 35038
rect 32498 34974 32510 35026
rect 32562 34974 32574 35026
rect 34862 34962 34914 34974
rect 38334 35026 38386 35038
rect 47630 35026 47682 35038
rect 40114 34974 40126 35026
rect 40178 34974 40190 35026
rect 42242 34974 42254 35026
rect 42306 34974 42318 35026
rect 38334 34962 38386 34974
rect 47630 34962 47682 34974
rect 33518 34914 33570 34926
rect 37886 34914 37938 34926
rect 29698 34862 29710 34914
rect 29762 34862 29774 34914
rect 34290 34862 34302 34914
rect 34354 34862 34366 34914
rect 35858 34862 35870 34914
rect 35922 34862 35934 34914
rect 39442 34862 39454 34914
rect 39506 34862 39518 34914
rect 33518 34850 33570 34862
rect 37886 34850 37938 34862
rect 37550 34802 37602 34814
rect 30370 34750 30382 34802
rect 30434 34750 30446 34802
rect 34066 34750 34078 34802
rect 34130 34750 34142 34802
rect 37550 34738 37602 34750
rect 44382 34802 44434 34814
rect 46498 34750 46510 34802
rect 46562 34750 46574 34802
rect 46946 34750 46958 34802
rect 47010 34750 47022 34802
rect 44382 34738 44434 34750
rect 1822 34690 1874 34702
rect 1822 34626 1874 34638
rect 33182 34690 33234 34702
rect 33182 34626 33234 34638
rect 35646 34690 35698 34702
rect 35646 34626 35698 34638
rect 36766 34690 36818 34702
rect 36766 34626 36818 34638
rect 38782 34690 38834 34702
rect 38782 34626 38834 34638
rect 43822 34690 43874 34702
rect 43822 34626 43874 34638
rect 44718 34690 44770 34702
rect 44718 34626 44770 34638
rect 1344 34522 48608 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 48608 34522
rect 1344 34436 48608 34470
rect 30494 34354 30546 34366
rect 30494 34290 30546 34302
rect 32846 34354 32898 34366
rect 32846 34290 32898 34302
rect 39230 34354 39282 34366
rect 39230 34290 39282 34302
rect 40798 34354 40850 34366
rect 40798 34290 40850 34302
rect 30830 34242 30882 34254
rect 34738 34190 34750 34242
rect 34802 34190 34814 34242
rect 38434 34190 38446 34242
rect 38498 34190 38510 34242
rect 42354 34190 42366 34242
rect 42418 34190 42430 34242
rect 45826 34190 45838 34242
rect 45890 34190 45902 34242
rect 30830 34178 30882 34190
rect 34066 34078 34078 34130
rect 34130 34078 34142 34130
rect 38546 34078 38558 34130
rect 38610 34078 38622 34130
rect 41682 34078 41694 34130
rect 41746 34078 41758 34130
rect 45042 34078 45054 34130
rect 45106 34078 45118 34130
rect 37886 34018 37938 34030
rect 36866 33966 36878 34018
rect 36930 33966 36942 34018
rect 37886 33954 37938 33966
rect 39678 34018 39730 34030
rect 44482 33966 44494 34018
rect 44546 33966 44558 34018
rect 47954 33966 47966 34018
rect 48018 33966 48030 34018
rect 39678 33954 39730 33966
rect 37550 33906 37602 33918
rect 37550 33842 37602 33854
rect 1344 33738 48608 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 48608 33738
rect 1344 33652 48608 33686
rect 45950 33570 46002 33582
rect 45950 33506 46002 33518
rect 47630 33458 47682 33470
rect 34178 33406 34190 33458
rect 34242 33406 34254 33458
rect 40450 33406 40462 33458
rect 40514 33406 40526 33458
rect 44034 33406 44046 33458
rect 44098 33406 44110 33458
rect 47630 33394 47682 33406
rect 35870 33346 35922 33358
rect 46286 33346 46338 33358
rect 31266 33294 31278 33346
rect 31330 33294 31342 33346
rect 36530 33294 36542 33346
rect 36594 33294 36606 33346
rect 37650 33294 37662 33346
rect 37714 33294 37726 33346
rect 44706 33294 44718 33346
rect 44770 33294 44782 33346
rect 35870 33282 35922 33294
rect 46286 33282 46338 33294
rect 32050 33182 32062 33234
rect 32114 33182 32126 33234
rect 36642 33182 36654 33234
rect 36706 33182 36718 33234
rect 38322 33182 38334 33234
rect 38386 33182 38398 33234
rect 46498 33182 46510 33234
rect 46562 33182 46574 33234
rect 46834 33182 46846 33234
rect 46898 33182 46910 33234
rect 34638 33122 34690 33134
rect 34638 33058 34690 33070
rect 35534 33122 35586 33134
rect 35534 33058 35586 33070
rect 1344 32954 48608 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 48608 32954
rect 1344 32868 48608 32902
rect 32286 32786 32338 32798
rect 32286 32722 32338 32734
rect 32622 32674 32674 32686
rect 45378 32622 45390 32674
rect 45442 32622 45454 32674
rect 32622 32610 32674 32622
rect 34862 32562 34914 32574
rect 39118 32562 39170 32574
rect 35522 32510 35534 32562
rect 35586 32510 35598 32562
rect 34862 32498 34914 32510
rect 39118 32498 39170 32510
rect 39678 32562 39730 32574
rect 39678 32498 39730 32510
rect 40798 32562 40850 32574
rect 40798 32498 40850 32510
rect 41470 32562 41522 32574
rect 44034 32510 44046 32562
rect 44098 32510 44110 32562
rect 44594 32510 44606 32562
rect 44658 32510 44670 32562
rect 41470 32498 41522 32510
rect 42254 32450 42306 32462
rect 36194 32398 36206 32450
rect 36258 32398 36270 32450
rect 38322 32398 38334 32450
rect 38386 32398 38398 32450
rect 40338 32398 40350 32450
rect 40402 32398 40414 32450
rect 43250 32398 43262 32450
rect 43314 32398 43326 32450
rect 47506 32398 47518 32450
rect 47570 32398 47582 32450
rect 42254 32386 42306 32398
rect 1344 32170 48608 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 48608 32170
rect 1344 32084 48608 32118
rect 36878 31890 36930 31902
rect 36878 31826 36930 31838
rect 35982 31778 36034 31790
rect 43598 31778 43650 31790
rect 37650 31726 37662 31778
rect 37714 31726 37726 31778
rect 45714 31726 45726 31778
rect 45778 31726 45790 31778
rect 35982 31714 36034 31726
rect 43598 31714 43650 31726
rect 36318 31666 36370 31678
rect 36318 31602 36370 31614
rect 37886 31666 37938 31678
rect 37886 31602 37938 31614
rect 44382 31666 44434 31678
rect 46610 31614 46622 31666
rect 46674 31614 46686 31666
rect 44382 31602 44434 31614
rect 39902 31554 39954 31566
rect 39902 31490 39954 31502
rect 42478 31554 42530 31566
rect 42478 31490 42530 31502
rect 43038 31554 43090 31566
rect 43038 31490 43090 31502
rect 44718 31554 44770 31566
rect 44718 31490 44770 31502
rect 1344 31386 48608 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 48608 31386
rect 1344 31300 48608 31334
rect 43374 31218 43426 31230
rect 43374 31154 43426 31166
rect 44706 31054 44718 31106
rect 44770 31054 44782 31106
rect 43922 30942 43934 30994
rect 43986 30942 43998 30994
rect 46834 30830 46846 30882
rect 46898 30830 46910 30882
rect 1344 30602 48608 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 48608 30602
rect 1344 30516 48608 30550
rect 46174 30434 46226 30446
rect 46174 30370 46226 30382
rect 44034 30270 44046 30322
rect 44098 30270 44110 30322
rect 45838 30210 45890 30222
rect 44706 30158 44718 30210
rect 44770 30158 44782 30210
rect 45838 30146 45890 30158
rect 47518 30098 47570 30110
rect 46386 30046 46398 30098
rect 46450 30046 46462 30098
rect 46722 30046 46734 30098
rect 46786 30046 46798 30098
rect 47518 30034 47570 30046
rect 1344 29818 48608 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 48608 29818
rect 1344 29732 48608 29766
rect 43810 29374 43822 29426
rect 43874 29374 43886 29426
rect 43262 29314 43314 29326
rect 44594 29262 44606 29314
rect 44658 29262 44670 29314
rect 46722 29262 46734 29314
rect 46786 29262 46798 29314
rect 43262 29250 43314 29262
rect 1344 29034 48608 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 48608 29034
rect 1344 28948 48608 28982
rect 45950 28866 46002 28878
rect 45950 28802 46002 28814
rect 3266 28702 3278 28754
rect 3330 28702 3342 28754
rect 45614 28642 45666 28654
rect 43474 28590 43486 28642
rect 43538 28590 43550 28642
rect 45614 28578 45666 28590
rect 38446 28530 38498 28542
rect 1922 28478 1934 28530
rect 1986 28478 1998 28530
rect 38446 28466 38498 28478
rect 42590 28530 42642 28542
rect 44594 28478 44606 28530
rect 44658 28478 44670 28530
rect 46162 28478 46174 28530
rect 46226 28478 46238 28530
rect 46722 28478 46734 28530
rect 46786 28478 46798 28530
rect 42590 28466 42642 28478
rect 38110 28418 38162 28430
rect 38110 28354 38162 28366
rect 42926 28418 42978 28430
rect 42926 28354 42978 28366
rect 1344 28250 48608 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 48608 28250
rect 1344 28164 48608 28198
rect 1822 28082 1874 28094
rect 1822 28018 1874 28030
rect 46286 28082 46338 28094
rect 46286 28018 46338 28030
rect 37538 27918 37550 27970
rect 37602 27918 37614 27970
rect 43586 27918 43598 27970
rect 43650 27918 43662 27970
rect 41582 27858 41634 27870
rect 46622 27858 46674 27870
rect 36866 27806 36878 27858
rect 36930 27806 36942 27858
rect 42802 27806 42814 27858
rect 42866 27806 42878 27858
rect 41582 27794 41634 27806
rect 46622 27794 46674 27806
rect 40126 27746 40178 27758
rect 39666 27694 39678 27746
rect 39730 27694 39742 27746
rect 40126 27682 40178 27694
rect 40798 27746 40850 27758
rect 42018 27694 42030 27746
rect 42082 27694 42094 27746
rect 45714 27694 45726 27746
rect 45778 27694 45790 27746
rect 40798 27682 40850 27694
rect 1344 27466 48608 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 48608 27466
rect 1344 27380 48608 27414
rect 46398 27298 46450 27310
rect 46398 27234 46450 27246
rect 46734 27298 46786 27310
rect 46734 27234 46786 27246
rect 42814 27186 42866 27198
rect 40450 27134 40462 27186
rect 40514 27134 40526 27186
rect 42814 27122 42866 27134
rect 43262 27186 43314 27198
rect 43262 27122 43314 27134
rect 41134 27074 41186 27086
rect 30482 27022 30494 27074
rect 30546 27022 30558 27074
rect 37650 27022 37662 27074
rect 37714 27022 37726 27074
rect 41134 27010 41186 27022
rect 41470 27074 41522 27086
rect 41470 27010 41522 27022
rect 29934 26962 29986 26974
rect 33618 26910 33630 26962
rect 33682 26910 33694 26962
rect 38322 26910 38334 26962
rect 38386 26910 38398 26962
rect 41682 26910 41694 26962
rect 41746 26910 41758 26962
rect 42130 26910 42142 26962
rect 42194 26910 42206 26962
rect 45602 26910 45614 26962
rect 45666 26910 45678 26962
rect 46162 26910 46174 26962
rect 46226 26910 46238 26962
rect 29934 26898 29986 26910
rect 1344 26682 48608 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 48608 26682
rect 1344 26596 48608 26630
rect 38446 26514 38498 26526
rect 38446 26450 38498 26462
rect 39454 26514 39506 26526
rect 39454 26450 39506 26462
rect 38782 26402 38834 26414
rect 40562 26350 40574 26402
rect 40626 26350 40638 26402
rect 46162 26350 46174 26402
rect 46226 26350 46238 26402
rect 38782 26338 38834 26350
rect 39790 26290 39842 26302
rect 40226 26238 40238 26290
rect 40290 26238 40302 26290
rect 41570 26238 41582 26290
rect 41634 26238 41646 26290
rect 45042 26238 45054 26290
rect 45106 26238 45118 26290
rect 39790 26226 39842 26238
rect 42354 26126 42366 26178
rect 42418 26126 42430 26178
rect 44482 26126 44494 26178
rect 44546 26126 44558 26178
rect 1344 25898 48608 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 48608 25898
rect 1344 25812 48608 25846
rect 41246 25618 41298 25630
rect 41246 25554 41298 25566
rect 44482 25454 44494 25506
rect 44546 25454 44558 25506
rect 45490 25454 45502 25506
rect 45554 25454 45566 25506
rect 42590 25394 42642 25406
rect 42590 25330 42642 25342
rect 42926 25394 42978 25406
rect 46610 25342 46622 25394
rect 46674 25342 46686 25394
rect 42926 25330 42978 25342
rect 44718 25282 44770 25294
rect 44718 25218 44770 25230
rect 1344 25114 48608 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 48608 25114
rect 1344 25028 48608 25062
rect 45266 24782 45278 24834
rect 45330 24782 45342 24834
rect 44594 24670 44606 24722
rect 44658 24670 44670 24722
rect 43934 24610 43986 24622
rect 47394 24558 47406 24610
rect 47458 24558 47470 24610
rect 43934 24546 43986 24558
rect 43698 24446 43710 24498
rect 43762 24495 43774 24498
rect 43922 24495 43934 24498
rect 43762 24449 43934 24495
rect 43762 24446 43774 24449
rect 43922 24446 43934 24449
rect 43986 24446 43998 24498
rect 1344 24330 48608 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 48608 24330
rect 1344 24244 48608 24278
rect 43486 24162 43538 24174
rect 43486 24098 43538 24110
rect 43822 24162 43874 24174
rect 43822 24098 43874 24110
rect 45950 24162 46002 24174
rect 45950 24098 46002 24110
rect 46286 24162 46338 24174
rect 46286 24098 46338 24110
rect 44370 23886 44382 23938
rect 44434 23886 44446 23938
rect 44482 23774 44494 23826
rect 44546 23774 44558 23826
rect 46498 23774 46510 23826
rect 46562 23774 46574 23826
rect 46834 23774 46846 23826
rect 46898 23774 46910 23826
rect 1344 23546 48608 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 48608 23546
rect 1344 23460 48608 23494
rect 40462 23378 40514 23390
rect 40462 23314 40514 23326
rect 42254 23378 42306 23390
rect 42254 23314 42306 23326
rect 6402 23214 6414 23266
rect 6466 23214 6478 23266
rect 37650 23214 37662 23266
rect 37714 23214 37726 23266
rect 33742 23154 33794 23166
rect 40126 23154 40178 23166
rect 5730 23102 5742 23154
rect 5794 23102 5806 23154
rect 34290 23102 34302 23154
rect 34354 23102 34366 23154
rect 43922 23102 43934 23154
rect 43986 23102 43998 23154
rect 44594 23102 44606 23154
rect 44658 23102 44670 23154
rect 33742 23090 33794 23102
rect 40126 23090 40178 23102
rect 8990 23042 9042 23054
rect 8530 22990 8542 23042
rect 8594 22990 8606 23042
rect 43362 22990 43374 23042
rect 43426 22990 43438 23042
rect 45378 22990 45390 23042
rect 45442 22990 45454 23042
rect 47506 22990 47518 23042
rect 47570 22990 47582 23042
rect 8990 22978 9042 22990
rect 1344 22762 48608 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 48608 22762
rect 1344 22676 48608 22710
rect 44034 22430 44046 22482
rect 44098 22430 44110 22482
rect 46734 22370 46786 22382
rect 44706 22318 44718 22370
rect 44770 22318 44782 22370
rect 45938 22318 45950 22370
rect 46002 22318 46014 22370
rect 46734 22306 46786 22318
rect 47070 22370 47122 22382
rect 47954 22318 47966 22370
rect 48018 22318 48030 22370
rect 47070 22306 47122 22318
rect 46162 22206 46174 22258
rect 46226 22206 46238 22258
rect 1822 22146 1874 22158
rect 1822 22082 1874 22094
rect 39790 22146 39842 22158
rect 39790 22082 39842 22094
rect 47742 22146 47794 22158
rect 47742 22082 47794 22094
rect 1344 21978 48608 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 48608 21978
rect 1344 21892 48608 21926
rect 43374 21810 43426 21822
rect 43374 21746 43426 21758
rect 43922 21534 43934 21586
rect 43986 21534 43998 21586
rect 44706 21422 44718 21474
rect 44770 21422 44782 21474
rect 46834 21422 46846 21474
rect 46898 21422 46910 21474
rect 1344 21194 48608 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 48608 21194
rect 1344 21108 48608 21142
rect 46174 21026 46226 21038
rect 46174 20962 46226 20974
rect 45838 20802 45890 20814
rect 44482 20750 44494 20802
rect 44546 20750 44558 20802
rect 45838 20738 45890 20750
rect 44718 20690 44770 20702
rect 46386 20638 46398 20690
rect 46450 20638 46462 20690
rect 46722 20638 46734 20690
rect 46786 20638 46798 20690
rect 44718 20626 44770 20638
rect 1344 20410 48608 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 48608 20410
rect 1344 20324 48608 20358
rect 30258 20078 30270 20130
rect 30322 20078 30334 20130
rect 43262 20018 43314 20030
rect 26786 19966 26798 20018
rect 26850 19966 26862 20018
rect 43262 19954 43314 19966
rect 43822 20018 43874 20030
rect 43822 19954 43874 19966
rect 44382 20018 44434 20030
rect 46162 19966 46174 20018
rect 46226 19966 46238 20018
rect 44382 19954 44434 19966
rect 26350 19906 26402 19918
rect 45266 19854 45278 19906
rect 45330 19854 45342 19906
rect 26350 19842 26402 19854
rect 1344 19626 48608 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 48608 19626
rect 1344 19540 48608 19574
rect 45714 19182 45726 19234
rect 45778 19182 45790 19234
rect 44718 19122 44770 19134
rect 46610 19070 46622 19122
rect 46674 19070 46686 19122
rect 44718 19058 44770 19070
rect 44382 19010 44434 19022
rect 44382 18946 44434 18958
rect 1344 18842 48608 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 48608 18842
rect 1344 18756 48608 18790
rect 44482 18510 44494 18562
rect 44546 18510 44558 18562
rect 43150 18450 43202 18462
rect 43698 18398 43710 18450
rect 43762 18398 43774 18450
rect 43150 18386 43202 18398
rect 46610 18286 46622 18338
rect 46674 18286 46686 18338
rect 1344 18058 48608 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 48608 18058
rect 1344 17972 48608 18006
rect 45614 17890 45666 17902
rect 45614 17826 45666 17838
rect 45950 17890 46002 17902
rect 45950 17826 46002 17838
rect 42926 17778 42978 17790
rect 42926 17714 42978 17726
rect 41806 17666 41858 17678
rect 44606 17666 44658 17678
rect 42466 17614 42478 17666
rect 42530 17614 42542 17666
rect 43698 17614 43710 17666
rect 43762 17614 43774 17666
rect 41806 17602 41858 17614
rect 44606 17602 44658 17614
rect 46162 17502 46174 17554
rect 46226 17502 46238 17554
rect 46498 17502 46510 17554
rect 46562 17502 46574 17554
rect 1344 17274 48608 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 48608 17274
rect 1344 17188 48608 17222
rect 38782 17106 38834 17118
rect 38782 17042 38834 17054
rect 47630 16994 47682 17006
rect 46274 16942 46286 16994
rect 46338 16942 46350 16994
rect 47630 16930 47682 16942
rect 37886 16882 37938 16894
rect 37886 16818 37938 16830
rect 38446 16882 38498 16894
rect 43586 16830 43598 16882
rect 43650 16830 43662 16882
rect 47058 16830 47070 16882
rect 47122 16830 47134 16882
rect 47842 16830 47854 16882
rect 47906 16830 47918 16882
rect 38446 16818 38498 16830
rect 42914 16718 42926 16770
rect 42978 16718 42990 16770
rect 44146 16718 44158 16770
rect 44210 16718 44222 16770
rect 1344 16490 48608 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 48608 16490
rect 1344 16404 48608 16438
rect 46398 16322 46450 16334
rect 46398 16258 46450 16270
rect 46734 16322 46786 16334
rect 46734 16258 46786 16270
rect 44494 16210 44546 16222
rect 3266 16158 3278 16210
rect 3330 16158 3342 16210
rect 44034 16158 44046 16210
rect 44098 16158 44110 16210
rect 44494 16146 44546 16158
rect 41234 16046 41246 16098
rect 41298 16046 41310 16098
rect 1922 15934 1934 15986
rect 1986 15934 1998 15986
rect 41906 15934 41918 15986
rect 41970 15934 41982 15986
rect 45602 15934 45614 15986
rect 45666 15934 45678 15986
rect 46162 15934 46174 15986
rect 46226 15934 46238 15986
rect 40574 15874 40626 15886
rect 40574 15810 40626 15822
rect 1344 15706 48608 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 48608 15706
rect 1344 15620 48608 15654
rect 1822 15538 1874 15550
rect 1822 15474 1874 15486
rect 42478 15538 42530 15550
rect 42478 15474 42530 15486
rect 21982 15426 22034 15438
rect 45042 15374 45054 15426
rect 45106 15374 45118 15426
rect 45490 15374 45502 15426
rect 45554 15374 45566 15426
rect 21982 15362 22034 15374
rect 21422 15314 21474 15326
rect 42814 15314 42866 15326
rect 21746 15262 21758 15314
rect 21810 15262 21822 15314
rect 21422 15250 21474 15262
rect 42814 15250 42866 15262
rect 44382 15314 44434 15326
rect 44382 15250 44434 15262
rect 44718 15314 44770 15326
rect 46162 15262 46174 15314
rect 46226 15262 46238 15314
rect 44718 15250 44770 15262
rect 20302 15202 20354 15214
rect 20302 15138 20354 15150
rect 20974 15202 21026 15214
rect 20974 15138 21026 15150
rect 22094 15202 22146 15214
rect 47282 15150 47294 15202
rect 47346 15150 47358 15202
rect 22094 15138 22146 15150
rect 1344 14922 48608 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 48608 14922
rect 1344 14836 48608 14870
rect 22094 14754 22146 14766
rect 22094 14690 22146 14702
rect 45950 14754 46002 14766
rect 45950 14690 46002 14702
rect 19954 14590 19966 14642
rect 20018 14590 20030 14642
rect 44706 14590 44718 14642
rect 44770 14590 44782 14642
rect 20526 14530 20578 14542
rect 17042 14478 17054 14530
rect 17106 14478 17118 14530
rect 20526 14466 20578 14478
rect 20862 14530 20914 14542
rect 41794 14478 41806 14530
rect 41858 14478 41870 14530
rect 20862 14466 20914 14478
rect 20638 14418 20690 14430
rect 17826 14366 17838 14418
rect 17890 14366 17902 14418
rect 20638 14354 20690 14366
rect 22206 14418 22258 14430
rect 42578 14366 42590 14418
rect 42642 14366 42654 14418
rect 46274 14366 46286 14418
rect 46338 14366 46350 14418
rect 46498 14366 46510 14418
rect 46562 14366 46574 14418
rect 22206 14354 22258 14366
rect 41246 14306 41298 14318
rect 41246 14242 41298 14254
rect 45614 14306 45666 14318
rect 45614 14242 45666 14254
rect 1344 14138 48608 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 48608 14138
rect 1344 14052 48608 14086
rect 10446 13970 10498 13982
rect 10446 13906 10498 13918
rect 43486 13970 43538 13982
rect 43486 13906 43538 13918
rect 43822 13858 43874 13870
rect 6850 13806 6862 13858
rect 6914 13806 6926 13858
rect 11778 13806 11790 13858
rect 11842 13806 11854 13858
rect 20178 13806 20190 13858
rect 20242 13806 20254 13858
rect 43822 13794 43874 13806
rect 14366 13746 14418 13758
rect 6178 13694 6190 13746
rect 6242 13694 6254 13746
rect 10994 13694 11006 13746
rect 11058 13694 11070 13746
rect 19394 13694 19406 13746
rect 19458 13694 19470 13746
rect 46162 13694 46174 13746
rect 46226 13694 46238 13746
rect 14366 13682 14418 13694
rect 9662 13634 9714 13646
rect 18846 13634 18898 13646
rect 22766 13634 22818 13646
rect 8978 13582 8990 13634
rect 9042 13582 9054 13634
rect 13906 13582 13918 13634
rect 13970 13582 13982 13634
rect 22306 13582 22318 13634
rect 22370 13582 22382 13634
rect 45266 13582 45278 13634
rect 45330 13582 45342 13634
rect 9662 13570 9714 13582
rect 18846 13570 18898 13582
rect 22766 13570 22818 13582
rect 1344 13354 48608 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 48608 13354
rect 1344 13268 48608 13302
rect 45714 12910 45726 12962
rect 45778 12910 45790 12962
rect 46610 12798 46622 12850
rect 46674 12798 46686 12850
rect 1344 12570 48608 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 48608 12570
rect 1344 12484 48608 12518
rect 16718 12402 16770 12414
rect 16718 12338 16770 12350
rect 33742 12402 33794 12414
rect 33742 12338 33794 12350
rect 43262 12290 43314 12302
rect 14130 12238 14142 12290
rect 14194 12238 14206 12290
rect 39330 12238 39342 12290
rect 39394 12238 39406 12290
rect 43262 12226 43314 12238
rect 24894 12178 24946 12190
rect 13458 12126 13470 12178
rect 13522 12126 13534 12178
rect 24434 12126 24446 12178
rect 24498 12126 24510 12178
rect 34290 12126 34302 12178
rect 34354 12126 34366 12178
rect 43810 12126 43822 12178
rect 43874 12126 43886 12178
rect 24894 12114 24946 12126
rect 16258 12014 16270 12066
rect 16322 12014 16334 12066
rect 21634 12014 21646 12066
rect 21698 12014 21710 12066
rect 44594 12014 44606 12066
rect 44658 12014 44670 12066
rect 46722 12014 46734 12066
rect 46786 12014 46798 12066
rect 1344 11786 48608 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 48608 11786
rect 1344 11700 48608 11734
rect 45950 11618 46002 11630
rect 45950 11554 46002 11566
rect 46722 11342 46734 11394
rect 46786 11342 46798 11394
rect 43822 11282 43874 11294
rect 43822 11218 43874 11230
rect 44382 11282 44434 11294
rect 44382 11218 44434 11230
rect 44718 11282 44770 11294
rect 44718 11218 44770 11230
rect 45614 11282 45666 11294
rect 46498 11230 46510 11282
rect 46562 11230 46574 11282
rect 45614 11218 45666 11230
rect 43486 11170 43538 11182
rect 43486 11106 43538 11118
rect 1344 11002 48608 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 48608 11002
rect 1344 10916 48608 10950
rect 42366 10834 42418 10846
rect 42366 10770 42418 10782
rect 46510 10834 46562 10846
rect 46510 10770 46562 10782
rect 39118 10722 39170 10734
rect 43698 10670 43710 10722
rect 43762 10670 43774 10722
rect 47058 10670 47070 10722
rect 47122 10670 47134 10722
rect 47394 10670 47406 10722
rect 47458 10670 47470 10722
rect 39118 10658 39170 10670
rect 39454 10610 39506 10622
rect 46846 10610 46898 10622
rect 42914 10558 42926 10610
rect 42978 10558 42990 10610
rect 39454 10546 39506 10558
rect 46846 10546 46898 10558
rect 45826 10446 45838 10498
rect 45890 10446 45902 10498
rect 1344 10218 48608 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 48608 10218
rect 1344 10132 48608 10166
rect 43598 9938 43650 9950
rect 38994 9886 39006 9938
rect 39058 9886 39070 9938
rect 41122 9886 41134 9938
rect 41186 9886 41198 9938
rect 43598 9874 43650 9886
rect 44718 9938 44770 9950
rect 46050 9886 46062 9938
rect 46114 9886 46126 9938
rect 44718 9874 44770 9886
rect 38210 9774 38222 9826
rect 38274 9774 38286 9826
rect 46610 9774 46622 9826
rect 46674 9774 46686 9826
rect 1822 9602 1874 9614
rect 1822 9538 1874 9550
rect 37662 9602 37714 9614
rect 37662 9538 37714 9550
rect 44158 9602 44210 9614
rect 44158 9538 44210 9550
rect 1344 9434 48608 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 48608 9434
rect 1344 9348 48608 9382
rect 39118 9266 39170 9278
rect 39118 9202 39170 9214
rect 39678 9266 39730 9278
rect 39678 9202 39730 9214
rect 46734 9154 46786 9166
rect 46734 9090 46786 9102
rect 47070 9042 47122 9054
rect 46050 8990 46062 9042
rect 46114 8990 46126 9042
rect 47070 8978 47122 8990
rect 38658 8878 38670 8930
rect 38722 8878 38734 8930
rect 45266 8878 45278 8930
rect 45330 8878 45342 8930
rect 1344 8650 48608 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 48608 8650
rect 1344 8564 48608 8598
rect 47070 8482 47122 8494
rect 47070 8418 47122 8430
rect 25790 8370 25842 8382
rect 16594 8318 16606 8370
rect 16658 8318 16670 8370
rect 25218 8318 25230 8370
rect 25282 8318 25294 8370
rect 25790 8306 25842 8318
rect 39454 8370 39506 8382
rect 39454 8306 39506 8318
rect 17054 8258 17106 8270
rect 26014 8258 26066 8270
rect 13794 8206 13806 8258
rect 13858 8206 13870 8258
rect 22306 8206 22318 8258
rect 22370 8206 22382 8258
rect 17054 8194 17106 8206
rect 26014 8194 26066 8206
rect 39790 8258 39842 8270
rect 46734 8258 46786 8270
rect 43586 8206 43598 8258
rect 43650 8206 43662 8258
rect 46274 8206 46286 8258
rect 46338 8206 46350 8258
rect 39790 8194 39842 8206
rect 46734 8194 46786 8206
rect 21758 8146 21810 8158
rect 38334 8146 38386 8158
rect 14466 8094 14478 8146
rect 14530 8094 14542 8146
rect 23090 8094 23102 8146
rect 23154 8094 23166 8146
rect 40002 8094 40014 8146
rect 40066 8094 40078 8146
rect 40450 8094 40462 8146
rect 40514 8094 40526 8146
rect 44594 8094 44606 8146
rect 44658 8094 44670 8146
rect 46050 8094 46062 8146
rect 46114 8094 46126 8146
rect 21758 8082 21810 8094
rect 38334 8082 38386 8094
rect 37998 8034 38050 8046
rect 26338 7982 26350 8034
rect 26402 7982 26414 8034
rect 37998 7970 38050 7982
rect 41134 8034 41186 8046
rect 41134 7970 41186 7982
rect 42926 8034 42978 8046
rect 42926 7970 42978 7982
rect 1344 7866 48608 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 48608 7866
rect 1344 7780 48608 7814
rect 21758 7698 21810 7710
rect 21758 7634 21810 7646
rect 25678 7698 25730 7710
rect 25678 7634 25730 7646
rect 37986 7534 37998 7586
rect 38050 7534 38062 7586
rect 45154 7534 45166 7586
rect 45218 7534 45230 7586
rect 40574 7474 40626 7486
rect 37314 7422 37326 7474
rect 37378 7422 37390 7474
rect 40574 7410 40626 7422
rect 43822 7474 43874 7486
rect 44370 7422 44382 7474
rect 44434 7422 44446 7474
rect 43822 7410 43874 7422
rect 40114 7310 40126 7362
rect 40178 7310 40190 7362
rect 47282 7310 47294 7362
rect 47346 7310 47358 7362
rect 1344 7082 48608 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 48608 7082
rect 1344 6996 48608 7030
rect 38558 6914 38610 6926
rect 38558 6850 38610 6862
rect 38894 6914 38946 6926
rect 38894 6850 38946 6862
rect 46734 6802 46786 6814
rect 46734 6738 46786 6750
rect 34862 6690 34914 6702
rect 34862 6626 34914 6638
rect 35870 6690 35922 6702
rect 47070 6690 47122 6702
rect 36642 6638 36654 6690
rect 36706 6638 36718 6690
rect 39554 6638 39566 6690
rect 39618 6638 39630 6690
rect 43474 6638 43486 6690
rect 43538 6638 43550 6690
rect 46274 6638 46286 6690
rect 46338 6638 46350 6690
rect 47954 6638 47966 6690
rect 48018 6638 48030 6690
rect 35870 6626 35922 6638
rect 47070 6626 47122 6638
rect 36418 6526 36430 6578
rect 36482 6526 36494 6578
rect 39666 6526 39678 6578
rect 39730 6526 39742 6578
rect 44594 6526 44606 6578
rect 44658 6526 44670 6578
rect 45938 6526 45950 6578
rect 46002 6526 46014 6578
rect 35534 6466 35586 6478
rect 35534 6402 35586 6414
rect 37438 6466 37490 6478
rect 37438 6402 37490 6414
rect 40350 6466 40402 6478
rect 40350 6402 40402 6414
rect 47742 6466 47794 6478
rect 47742 6402 47794 6414
rect 1344 6298 48608 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 48608 6298
rect 1344 6212 48608 6246
rect 38894 6130 38946 6142
rect 38894 6066 38946 6078
rect 44158 6130 44210 6142
rect 44158 6066 44210 6078
rect 35086 6018 35138 6030
rect 35086 5954 35138 5966
rect 35422 6018 35474 6030
rect 36754 5966 36766 6018
rect 36818 5966 36830 6018
rect 37314 5966 37326 6018
rect 37378 5966 37390 6018
rect 46834 5966 46846 6018
rect 46898 5966 46910 6018
rect 35422 5954 35474 5966
rect 37550 5906 37602 5918
rect 47506 5854 47518 5906
rect 47570 5854 47582 5906
rect 37550 5842 37602 5854
rect 38446 5794 38498 5806
rect 44706 5742 44718 5794
rect 44770 5742 44782 5794
rect 38446 5730 38498 5742
rect 37886 5682 37938 5694
rect 37886 5618 37938 5630
rect 1344 5514 48608 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 48608 5514
rect 1344 5428 48608 5462
rect 9214 5234 9266 5246
rect 38334 5234 38386 5246
rect 6514 5182 6526 5234
rect 6578 5182 6590 5234
rect 8642 5182 8654 5234
rect 8706 5182 8718 5234
rect 34626 5182 34638 5234
rect 34690 5182 34702 5234
rect 36754 5182 36766 5234
rect 36818 5182 36830 5234
rect 9214 5170 9266 5182
rect 38334 5170 38386 5182
rect 44830 5234 44882 5246
rect 44830 5170 44882 5182
rect 37886 5122 37938 5134
rect 5842 5070 5854 5122
rect 5906 5070 5918 5122
rect 33954 5070 33966 5122
rect 34018 5070 34030 5122
rect 37886 5058 37938 5070
rect 44270 5122 44322 5134
rect 46622 5122 46674 5134
rect 45490 5070 45502 5122
rect 45554 5070 45566 5122
rect 47506 5070 47518 5122
rect 47570 5070 47582 5122
rect 44270 5058 44322 5070
rect 46622 5058 46674 5070
rect 37550 4898 37602 4910
rect 47282 4846 47294 4898
rect 47346 4846 47358 4898
rect 37550 4834 37602 4846
rect 1344 4730 48608 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 48608 4730
rect 1344 4644 48608 4678
rect 38782 4562 38834 4574
rect 38782 4498 38834 4510
rect 44606 4562 44658 4574
rect 44606 4498 44658 4510
rect 46958 4562 47010 4574
rect 46958 4498 47010 4510
rect 36194 4398 36206 4450
rect 36258 4398 36270 4450
rect 44930 4398 44942 4450
rect 44994 4398 45006 4450
rect 35522 4286 35534 4338
rect 35586 4286 35598 4338
rect 1822 4226 1874 4238
rect 38322 4174 38334 4226
rect 38386 4174 38398 4226
rect 1822 4162 1874 4174
rect 1344 3946 48608 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 48608 3946
rect 1344 3860 48608 3894
rect 3266 3614 3278 3666
rect 3330 3614 3342 3666
rect 44270 3554 44322 3566
rect 44930 3502 44942 3554
rect 44994 3502 45006 3554
rect 44270 3490 44322 3502
rect 1922 3390 1934 3442
rect 1986 3390 1998 3442
rect 46050 3390 46062 3442
rect 46114 3390 46126 3442
rect 8654 3330 8706 3342
rect 8654 3266 8706 3278
rect 14142 3330 14194 3342
rect 14142 3266 14194 3278
rect 19630 3330 19682 3342
rect 19630 3266 19682 3278
rect 25342 3330 25394 3342
rect 25342 3266 25394 3278
rect 1344 3162 48608 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 48608 3162
rect 1344 3076 48608 3110
<< via1 >>
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 1822 46062 1874 46114
rect 47854 45950 47906 46002
rect 44942 45838 44994 45890
rect 46734 45838 46786 45890
rect 46062 45726 46114 45778
rect 44158 45614 44210 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 44942 45054 44994 45106
rect 44494 44942 44546 44994
rect 45950 44942 46002 44994
rect 46622 44942 46674 44994
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 44718 44270 44770 44322
rect 45502 44270 45554 44322
rect 46622 44158 46674 44210
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 45502 42702 45554 42754
rect 46622 42590 46674 42642
rect 44718 42478 44770 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 3054 41134 3106 41186
rect 44718 41134 44770 41186
rect 45502 41134 45554 41186
rect 1934 41022 1986 41074
rect 46622 41022 46674 41074
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 3278 40574 3330 40626
rect 3614 40350 3666 40402
rect 4062 40350 4114 40402
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 45502 39566 45554 39618
rect 46622 39454 46674 39506
rect 44718 39342 44770 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 44942 38782 44994 38834
rect 46062 38670 46114 38722
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 45726 37998 45778 38050
rect 46622 37886 46674 37938
rect 47182 37774 47234 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 39454 37438 39506 37490
rect 39902 37438 39954 37490
rect 43374 37438 43426 37490
rect 42366 37326 42418 37378
rect 42814 37326 42866 37378
rect 42030 37214 42082 37266
rect 46174 37214 46226 37266
rect 45278 37102 45330 37154
rect 41694 36990 41746 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 38334 36654 38386 36706
rect 40238 36654 40290 36706
rect 42142 36654 42194 36706
rect 35646 36542 35698 36594
rect 36878 36542 36930 36594
rect 43486 36430 43538 36482
rect 44494 36430 44546 36482
rect 46734 36430 46786 36482
rect 38670 36318 38722 36370
rect 39118 36318 39170 36370
rect 40462 36318 40514 36370
rect 41022 36318 41074 36370
rect 42366 36318 42418 36370
rect 42926 36318 42978 36370
rect 46174 36318 46226 36370
rect 46510 36318 46562 36370
rect 47630 36318 47682 36370
rect 35198 36206 35250 36258
rect 36206 36206 36258 36258
rect 37998 36206 38050 36258
rect 39902 36206 39954 36258
rect 41806 36206 41858 36258
rect 44718 36206 44770 36258
rect 47070 36206 47122 36258
rect 48078 36206 48130 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 42366 35870 42418 35922
rect 34302 35758 34354 35810
rect 34862 35758 34914 35810
rect 40126 35758 40178 35810
rect 40462 35758 40514 35810
rect 41918 35758 41970 35810
rect 45054 35758 45106 35810
rect 47742 35758 47794 35810
rect 35982 35646 36034 35698
rect 41694 35646 41746 35698
rect 44270 35646 44322 35698
rect 47966 35646 48018 35698
rect 32734 35534 32786 35586
rect 36654 35534 36706 35586
rect 38782 35534 38834 35586
rect 39230 35534 39282 35586
rect 43822 35534 43874 35586
rect 47182 35534 47234 35586
rect 33742 35422 33794 35474
rect 34078 35422 34130 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 45950 35086 46002 35138
rect 46286 35086 46338 35138
rect 32510 34974 32562 35026
rect 34862 34974 34914 35026
rect 38334 34974 38386 35026
rect 40126 34974 40178 35026
rect 42254 34974 42306 35026
rect 47630 34974 47682 35026
rect 29710 34862 29762 34914
rect 33518 34862 33570 34914
rect 34302 34862 34354 34914
rect 35870 34862 35922 34914
rect 37886 34862 37938 34914
rect 39454 34862 39506 34914
rect 30382 34750 30434 34802
rect 34078 34750 34130 34802
rect 37550 34750 37602 34802
rect 44382 34750 44434 34802
rect 46510 34750 46562 34802
rect 46958 34750 47010 34802
rect 1822 34638 1874 34690
rect 33182 34638 33234 34690
rect 35646 34638 35698 34690
rect 36766 34638 36818 34690
rect 38782 34638 38834 34690
rect 43822 34638 43874 34690
rect 44718 34638 44770 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 30494 34302 30546 34354
rect 32846 34302 32898 34354
rect 39230 34302 39282 34354
rect 40798 34302 40850 34354
rect 30830 34190 30882 34242
rect 34750 34190 34802 34242
rect 38446 34190 38498 34242
rect 42366 34190 42418 34242
rect 45838 34190 45890 34242
rect 34078 34078 34130 34130
rect 38558 34078 38610 34130
rect 41694 34078 41746 34130
rect 45054 34078 45106 34130
rect 36878 33966 36930 34018
rect 37886 33966 37938 34018
rect 39678 33966 39730 34018
rect 44494 33966 44546 34018
rect 47966 33966 48018 34018
rect 37550 33854 37602 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 45950 33518 46002 33570
rect 34190 33406 34242 33458
rect 40462 33406 40514 33458
rect 44046 33406 44098 33458
rect 47630 33406 47682 33458
rect 31278 33294 31330 33346
rect 35870 33294 35922 33346
rect 36542 33294 36594 33346
rect 37662 33294 37714 33346
rect 44718 33294 44770 33346
rect 46286 33294 46338 33346
rect 32062 33182 32114 33234
rect 36654 33182 36706 33234
rect 38334 33182 38386 33234
rect 46510 33182 46562 33234
rect 46846 33182 46898 33234
rect 34638 33070 34690 33122
rect 35534 33070 35586 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 32286 32734 32338 32786
rect 32622 32622 32674 32674
rect 45390 32622 45442 32674
rect 34862 32510 34914 32562
rect 35534 32510 35586 32562
rect 39118 32510 39170 32562
rect 39678 32510 39730 32562
rect 40798 32510 40850 32562
rect 41470 32510 41522 32562
rect 44046 32510 44098 32562
rect 44606 32510 44658 32562
rect 36206 32398 36258 32450
rect 38334 32398 38386 32450
rect 40350 32398 40402 32450
rect 42254 32398 42306 32450
rect 43262 32398 43314 32450
rect 47518 32398 47570 32450
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 36878 31838 36930 31890
rect 35982 31726 36034 31778
rect 37662 31726 37714 31778
rect 43598 31726 43650 31778
rect 45726 31726 45778 31778
rect 36318 31614 36370 31666
rect 37886 31614 37938 31666
rect 44382 31614 44434 31666
rect 46622 31614 46674 31666
rect 39902 31502 39954 31554
rect 42478 31502 42530 31554
rect 43038 31502 43090 31554
rect 44718 31502 44770 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 43374 31166 43426 31218
rect 44718 31054 44770 31106
rect 43934 30942 43986 30994
rect 46846 30830 46898 30882
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 46174 30382 46226 30434
rect 44046 30270 44098 30322
rect 44718 30158 44770 30210
rect 45838 30158 45890 30210
rect 46398 30046 46450 30098
rect 46734 30046 46786 30098
rect 47518 30046 47570 30098
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 43822 29374 43874 29426
rect 43262 29262 43314 29314
rect 44606 29262 44658 29314
rect 46734 29262 46786 29314
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 45950 28814 46002 28866
rect 3278 28702 3330 28754
rect 43486 28590 43538 28642
rect 45614 28590 45666 28642
rect 1934 28478 1986 28530
rect 38446 28478 38498 28530
rect 42590 28478 42642 28530
rect 44606 28478 44658 28530
rect 46174 28478 46226 28530
rect 46734 28478 46786 28530
rect 38110 28366 38162 28418
rect 42926 28366 42978 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 1822 28030 1874 28082
rect 46286 28030 46338 28082
rect 37550 27918 37602 27970
rect 43598 27918 43650 27970
rect 36878 27806 36930 27858
rect 41582 27806 41634 27858
rect 42814 27806 42866 27858
rect 46622 27806 46674 27858
rect 39678 27694 39730 27746
rect 40126 27694 40178 27746
rect 40798 27694 40850 27746
rect 42030 27694 42082 27746
rect 45726 27694 45778 27746
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 46398 27246 46450 27298
rect 46734 27246 46786 27298
rect 40462 27134 40514 27186
rect 42814 27134 42866 27186
rect 43262 27134 43314 27186
rect 30494 27022 30546 27074
rect 37662 27022 37714 27074
rect 41134 27022 41186 27074
rect 41470 27022 41522 27074
rect 29934 26910 29986 26962
rect 33630 26910 33682 26962
rect 38334 26910 38386 26962
rect 41694 26910 41746 26962
rect 42142 26910 42194 26962
rect 45614 26910 45666 26962
rect 46174 26910 46226 26962
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 38446 26462 38498 26514
rect 39454 26462 39506 26514
rect 38782 26350 38834 26402
rect 40574 26350 40626 26402
rect 46174 26350 46226 26402
rect 39790 26238 39842 26290
rect 40238 26238 40290 26290
rect 41582 26238 41634 26290
rect 45054 26238 45106 26290
rect 42366 26126 42418 26178
rect 44494 26126 44546 26178
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 41246 25566 41298 25618
rect 44494 25454 44546 25506
rect 45502 25454 45554 25506
rect 42590 25342 42642 25394
rect 42926 25342 42978 25394
rect 46622 25342 46674 25394
rect 44718 25230 44770 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 45278 24782 45330 24834
rect 44606 24670 44658 24722
rect 43934 24558 43986 24610
rect 47406 24558 47458 24610
rect 43710 24446 43762 24498
rect 43934 24446 43986 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 43486 24110 43538 24162
rect 43822 24110 43874 24162
rect 45950 24110 46002 24162
rect 46286 24110 46338 24162
rect 44382 23886 44434 23938
rect 44494 23774 44546 23826
rect 46510 23774 46562 23826
rect 46846 23774 46898 23826
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 40462 23326 40514 23378
rect 42254 23326 42306 23378
rect 6414 23214 6466 23266
rect 37662 23214 37714 23266
rect 5742 23102 5794 23154
rect 33742 23102 33794 23154
rect 34302 23102 34354 23154
rect 40126 23102 40178 23154
rect 43934 23102 43986 23154
rect 44606 23102 44658 23154
rect 8542 22990 8594 23042
rect 8990 22990 9042 23042
rect 43374 22990 43426 23042
rect 45390 22990 45442 23042
rect 47518 22990 47570 23042
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 44046 22430 44098 22482
rect 44718 22318 44770 22370
rect 45950 22318 46002 22370
rect 46734 22318 46786 22370
rect 47070 22318 47122 22370
rect 47966 22318 48018 22370
rect 46174 22206 46226 22258
rect 1822 22094 1874 22146
rect 39790 22094 39842 22146
rect 47742 22094 47794 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 43374 21758 43426 21810
rect 43934 21534 43986 21586
rect 44718 21422 44770 21474
rect 46846 21422 46898 21474
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 46174 20974 46226 21026
rect 44494 20750 44546 20802
rect 45838 20750 45890 20802
rect 44718 20638 44770 20690
rect 46398 20638 46450 20690
rect 46734 20638 46786 20690
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 30270 20078 30322 20130
rect 26798 19966 26850 20018
rect 43262 19966 43314 20018
rect 43822 19966 43874 20018
rect 44382 19966 44434 20018
rect 46174 19966 46226 20018
rect 26350 19854 26402 19906
rect 45278 19854 45330 19906
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 45726 19182 45778 19234
rect 44718 19070 44770 19122
rect 46622 19070 46674 19122
rect 44382 18958 44434 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 44494 18510 44546 18562
rect 43150 18398 43202 18450
rect 43710 18398 43762 18450
rect 46622 18286 46674 18338
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 45614 17838 45666 17890
rect 45950 17838 46002 17890
rect 42926 17726 42978 17778
rect 41806 17614 41858 17666
rect 42478 17614 42530 17666
rect 43710 17614 43762 17666
rect 44606 17614 44658 17666
rect 46174 17502 46226 17554
rect 46510 17502 46562 17554
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 38782 17054 38834 17106
rect 46286 16942 46338 16994
rect 47630 16942 47682 16994
rect 37886 16830 37938 16882
rect 38446 16830 38498 16882
rect 43598 16830 43650 16882
rect 47070 16830 47122 16882
rect 47854 16830 47906 16882
rect 42926 16718 42978 16770
rect 44158 16718 44210 16770
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 46398 16270 46450 16322
rect 46734 16270 46786 16322
rect 3278 16158 3330 16210
rect 44046 16158 44098 16210
rect 44494 16158 44546 16210
rect 41246 16046 41298 16098
rect 1934 15934 1986 15986
rect 41918 15934 41970 15986
rect 45614 15934 45666 15986
rect 46174 15934 46226 15986
rect 40574 15822 40626 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 1822 15486 1874 15538
rect 42478 15486 42530 15538
rect 21982 15374 22034 15426
rect 45054 15374 45106 15426
rect 45502 15374 45554 15426
rect 21422 15262 21474 15314
rect 21758 15262 21810 15314
rect 42814 15262 42866 15314
rect 44382 15262 44434 15314
rect 44718 15262 44770 15314
rect 46174 15262 46226 15314
rect 20302 15150 20354 15202
rect 20974 15150 21026 15202
rect 22094 15150 22146 15202
rect 47294 15150 47346 15202
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 22094 14702 22146 14754
rect 45950 14702 46002 14754
rect 19966 14590 20018 14642
rect 44718 14590 44770 14642
rect 17054 14478 17106 14530
rect 20526 14478 20578 14530
rect 20862 14478 20914 14530
rect 41806 14478 41858 14530
rect 17838 14366 17890 14418
rect 20638 14366 20690 14418
rect 22206 14366 22258 14418
rect 42590 14366 42642 14418
rect 46286 14366 46338 14418
rect 46510 14366 46562 14418
rect 41246 14254 41298 14306
rect 45614 14254 45666 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 10446 13918 10498 13970
rect 43486 13918 43538 13970
rect 6862 13806 6914 13858
rect 11790 13806 11842 13858
rect 20190 13806 20242 13858
rect 43822 13806 43874 13858
rect 6190 13694 6242 13746
rect 11006 13694 11058 13746
rect 14366 13694 14418 13746
rect 19406 13694 19458 13746
rect 46174 13694 46226 13746
rect 8990 13582 9042 13634
rect 9662 13582 9714 13634
rect 13918 13582 13970 13634
rect 18846 13582 18898 13634
rect 22318 13582 22370 13634
rect 22766 13582 22818 13634
rect 45278 13582 45330 13634
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 45726 12910 45778 12962
rect 46622 12798 46674 12850
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 16718 12350 16770 12402
rect 33742 12350 33794 12402
rect 14142 12238 14194 12290
rect 39342 12238 39394 12290
rect 43262 12238 43314 12290
rect 13470 12126 13522 12178
rect 24446 12126 24498 12178
rect 24894 12126 24946 12178
rect 34302 12126 34354 12178
rect 43822 12126 43874 12178
rect 16270 12014 16322 12066
rect 21646 12014 21698 12066
rect 44606 12014 44658 12066
rect 46734 12014 46786 12066
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 45950 11566 46002 11618
rect 46734 11342 46786 11394
rect 43822 11230 43874 11282
rect 44382 11230 44434 11282
rect 44718 11230 44770 11282
rect 45614 11230 45666 11282
rect 46510 11230 46562 11282
rect 43486 11118 43538 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 42366 10782 42418 10834
rect 46510 10782 46562 10834
rect 39118 10670 39170 10722
rect 43710 10670 43762 10722
rect 47070 10670 47122 10722
rect 47406 10670 47458 10722
rect 39454 10558 39506 10610
rect 42926 10558 42978 10610
rect 46846 10558 46898 10610
rect 45838 10446 45890 10498
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 39006 9886 39058 9938
rect 41134 9886 41186 9938
rect 43598 9886 43650 9938
rect 44718 9886 44770 9938
rect 46062 9886 46114 9938
rect 38222 9774 38274 9826
rect 46622 9774 46674 9826
rect 1822 9550 1874 9602
rect 37662 9550 37714 9602
rect 44158 9550 44210 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 39118 9214 39170 9266
rect 39678 9214 39730 9266
rect 46734 9102 46786 9154
rect 46062 8990 46114 9042
rect 47070 8990 47122 9042
rect 38670 8878 38722 8930
rect 45278 8878 45330 8930
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 47070 8430 47122 8482
rect 16606 8318 16658 8370
rect 25230 8318 25282 8370
rect 25790 8318 25842 8370
rect 39454 8318 39506 8370
rect 13806 8206 13858 8258
rect 17054 8206 17106 8258
rect 22318 8206 22370 8258
rect 26014 8206 26066 8258
rect 39790 8206 39842 8258
rect 43598 8206 43650 8258
rect 46286 8206 46338 8258
rect 46734 8206 46786 8258
rect 14478 8094 14530 8146
rect 21758 8094 21810 8146
rect 23102 8094 23154 8146
rect 38334 8094 38386 8146
rect 40014 8094 40066 8146
rect 40462 8094 40514 8146
rect 44606 8094 44658 8146
rect 46062 8094 46114 8146
rect 26350 7982 26402 8034
rect 37998 7982 38050 8034
rect 41134 7982 41186 8034
rect 42926 7982 42978 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 21758 7646 21810 7698
rect 25678 7646 25730 7698
rect 37998 7534 38050 7586
rect 45166 7534 45218 7586
rect 37326 7422 37378 7474
rect 40574 7422 40626 7474
rect 43822 7422 43874 7474
rect 44382 7422 44434 7474
rect 40126 7310 40178 7362
rect 47294 7310 47346 7362
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 38558 6862 38610 6914
rect 38894 6862 38946 6914
rect 46734 6750 46786 6802
rect 34862 6638 34914 6690
rect 35870 6638 35922 6690
rect 36654 6638 36706 6690
rect 39566 6638 39618 6690
rect 43486 6638 43538 6690
rect 46286 6638 46338 6690
rect 47070 6638 47122 6690
rect 47966 6638 48018 6690
rect 36430 6526 36482 6578
rect 39678 6526 39730 6578
rect 44606 6526 44658 6578
rect 45950 6526 46002 6578
rect 35534 6414 35586 6466
rect 37438 6414 37490 6466
rect 40350 6414 40402 6466
rect 47742 6414 47794 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 38894 6078 38946 6130
rect 44158 6078 44210 6130
rect 35086 5966 35138 6018
rect 35422 5966 35474 6018
rect 36766 5966 36818 6018
rect 37326 5966 37378 6018
rect 46846 5966 46898 6018
rect 37550 5854 37602 5906
rect 47518 5854 47570 5906
rect 38446 5742 38498 5794
rect 44718 5742 44770 5794
rect 37886 5630 37938 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 6526 5182 6578 5234
rect 8654 5182 8706 5234
rect 9214 5182 9266 5234
rect 34638 5182 34690 5234
rect 36766 5182 36818 5234
rect 38334 5182 38386 5234
rect 44830 5182 44882 5234
rect 5854 5070 5906 5122
rect 33966 5070 34018 5122
rect 37886 5070 37938 5122
rect 44270 5070 44322 5122
rect 45502 5070 45554 5122
rect 46622 5070 46674 5122
rect 47518 5070 47570 5122
rect 37550 4846 37602 4898
rect 47294 4846 47346 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 38782 4510 38834 4562
rect 44606 4510 44658 4562
rect 46958 4510 47010 4562
rect 36206 4398 36258 4450
rect 44942 4398 44994 4450
rect 35534 4286 35586 4338
rect 1822 4174 1874 4226
rect 38334 4174 38386 4226
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 3278 3614 3330 3666
rect 44270 3502 44322 3554
rect 44942 3502 44994 3554
rect 1934 3390 1986 3442
rect 46062 3390 46114 3442
rect 8654 3278 8706 3330
rect 14142 3278 14194 3330
rect 19630 3278 19682 3330
rect 25342 3278 25394 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 47852 48244 47908 48254
rect 45948 46788 46004 46798
rect 1820 46564 1876 46574
rect 1820 46114 1876 46508
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 1820 46062 1822 46114
rect 1874 46062 1876 46114
rect 1820 46050 1876 46062
rect 44940 45892 44996 45902
rect 44156 45890 44996 45892
rect 44156 45838 44942 45890
rect 44994 45838 44996 45890
rect 44156 45836 44996 45838
rect 44156 45666 44212 45836
rect 44940 45826 44996 45836
rect 44156 45614 44158 45666
rect 44210 45614 44212 45666
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 3052 41188 3108 41198
rect 39900 41188 39956 41198
rect 3052 41186 3332 41188
rect 3052 41134 3054 41186
rect 3106 41134 3332 41186
rect 3052 41132 3332 41134
rect 3052 41122 3108 41132
rect 1932 41074 1988 41086
rect 1932 41022 1934 41074
rect 1986 41022 1988 41074
rect 1932 40404 1988 41022
rect 3276 40626 3332 41132
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 3276 40574 3278 40626
rect 3330 40574 3332 40626
rect 3276 40562 3332 40574
rect 1932 40338 1988 40348
rect 3612 40404 3668 40414
rect 4060 40404 4116 40414
rect 3612 40402 4116 40404
rect 3612 40350 3614 40402
rect 3666 40350 4062 40402
rect 4114 40350 4116 40402
rect 3612 40348 4116 40350
rect 3612 40338 3668 40348
rect 1820 34690 1876 34702
rect 1820 34638 1822 34690
rect 1874 34638 1876 34690
rect 1820 34244 1876 34638
rect 1820 34178 1876 34188
rect 4060 34020 4116 40348
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 39452 37492 39508 37502
rect 39900 37492 39956 41132
rect 42028 37492 42084 37502
rect 39452 37490 40292 37492
rect 39452 37438 39454 37490
rect 39506 37438 39902 37490
rect 39954 37438 40292 37490
rect 39452 37436 40292 37438
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35644 36820 35700 36830
rect 35644 36594 35700 36764
rect 35644 36542 35646 36594
rect 35698 36542 35700 36594
rect 35196 36258 35252 36270
rect 35196 36206 35198 36258
rect 35250 36206 35252 36258
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 34300 35810 34356 35822
rect 34300 35758 34302 35810
rect 34354 35758 34356 35810
rect 32732 35588 32788 35598
rect 32732 35494 32788 35532
rect 33964 35588 34020 35598
rect 33740 35474 33796 35486
rect 33740 35422 33742 35474
rect 33794 35422 33796 35474
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 32508 35026 32564 35038
rect 32508 34974 32510 35026
rect 32562 34974 32564 35026
rect 29708 34916 29764 34926
rect 29708 34822 29764 34860
rect 31276 34916 31332 34926
rect 30380 34802 30436 34814
rect 30380 34750 30382 34802
rect 30434 34750 30436 34802
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 30380 34356 30436 34750
rect 30492 34356 30548 34366
rect 30380 34354 30548 34356
rect 30380 34302 30494 34354
rect 30546 34302 30548 34354
rect 30380 34300 30548 34302
rect 30492 34290 30548 34300
rect 30828 34244 30884 34254
rect 30828 34150 30884 34188
rect 4060 33954 4116 33964
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 31276 33348 31332 34860
rect 32508 34356 32564 34974
rect 32508 34020 32564 34300
rect 32508 33954 32564 33964
rect 32620 35028 32676 35038
rect 31276 33216 31332 33292
rect 32060 33236 32116 33246
rect 32060 33234 32340 33236
rect 32060 33182 32062 33234
rect 32114 33182 32340 33234
rect 32060 33180 32340 33182
rect 32060 33170 32116 33180
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 32284 32786 32340 33180
rect 32284 32734 32286 32786
rect 32338 32734 32340 32786
rect 32284 32722 32340 32734
rect 32620 32674 32676 34972
rect 33740 35028 33796 35422
rect 33740 34962 33796 34972
rect 33516 34914 33572 34926
rect 33516 34862 33518 34914
rect 33570 34862 33572 34914
rect 33180 34690 33236 34702
rect 33180 34638 33182 34690
rect 33234 34638 33236 34690
rect 32844 34356 32900 34366
rect 32844 34262 32900 34300
rect 33180 34244 33236 34638
rect 33516 34356 33572 34862
rect 33516 34290 33572 34300
rect 33180 34178 33236 34188
rect 33964 34132 34020 35532
rect 34076 35476 34132 35486
rect 34076 34804 34132 35420
rect 34300 34916 34356 35758
rect 34860 35812 34916 35822
rect 35196 35812 35252 36206
rect 34860 35810 35252 35812
rect 34860 35758 34862 35810
rect 34914 35758 35252 35810
rect 34860 35756 35252 35758
rect 34860 35746 34916 35756
rect 34860 35588 34916 35598
rect 34860 35026 34916 35532
rect 35196 35476 35252 35756
rect 35644 35588 35700 36542
rect 36876 36708 36932 36718
rect 36876 36594 36932 36652
rect 36876 36542 36878 36594
rect 36930 36542 36932 36594
rect 36204 36258 36260 36270
rect 36204 36206 36206 36258
rect 36258 36206 36260 36258
rect 35644 35522 35700 35532
rect 35980 35700 36036 35710
rect 36204 35700 36260 36206
rect 35980 35698 36260 35700
rect 35980 35646 35982 35698
rect 36034 35646 36260 35698
rect 35980 35644 36260 35646
rect 35196 35410 35252 35420
rect 35868 35364 35924 35374
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 34860 34974 34862 35026
rect 34914 34974 34916 35026
rect 34860 34962 34916 34974
rect 34300 34822 34356 34860
rect 35868 34914 35924 35308
rect 35980 35028 36036 35644
rect 35980 34962 36036 34972
rect 36652 35586 36708 35598
rect 36652 35534 36654 35586
rect 36706 35534 36708 35586
rect 35868 34862 35870 34914
rect 35922 34862 35924 34914
rect 35868 34850 35924 34862
rect 36540 34916 36596 34926
rect 34076 34802 34244 34804
rect 34076 34750 34078 34802
rect 34130 34750 34244 34802
rect 34076 34748 34244 34750
rect 34076 34738 34132 34748
rect 34076 34132 34132 34142
rect 33964 34076 34076 34132
rect 34076 34038 34132 34076
rect 34188 33458 34244 34748
rect 35644 34690 35700 34702
rect 35644 34638 35646 34690
rect 35698 34638 35700 34690
rect 34748 34244 34804 34254
rect 34748 34150 34804 34188
rect 35644 34244 35700 34638
rect 35644 34178 35700 34188
rect 34188 33406 34190 33458
rect 34242 33406 34244 33458
rect 34188 33394 34244 33406
rect 34636 34132 34692 34142
rect 32620 32622 32622 32674
rect 32674 32622 32676 32674
rect 32620 32610 32676 32622
rect 34636 33348 34692 34076
rect 36540 34132 36596 34860
rect 36652 34804 36708 35534
rect 36652 34738 36708 34748
rect 36764 35028 36820 35038
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35644 33684 35700 33694
rect 34636 33122 34692 33292
rect 35532 33124 35588 33134
rect 34636 33070 34638 33122
rect 34690 33070 34692 33122
rect 34636 32564 34692 33070
rect 35420 33122 35588 33124
rect 35420 33070 35534 33122
rect 35586 33070 35588 33122
rect 35420 33068 35588 33070
rect 34860 32564 34916 32574
rect 34636 32508 34860 32564
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 3276 28756 3332 28766
rect 3276 28754 3444 28756
rect 3276 28702 3278 28754
rect 3330 28702 3444 28754
rect 3276 28700 3444 28702
rect 3276 28690 3332 28700
rect 1932 28532 1988 28542
rect 1820 28530 1988 28532
rect 1820 28478 1934 28530
rect 1986 28478 1988 28530
rect 1820 28476 1988 28478
rect 1820 28084 1876 28476
rect 1932 28466 1988 28476
rect 1820 27990 1876 28028
rect 3388 26964 3444 28700
rect 34860 28532 34916 32508
rect 35420 32340 35476 33068
rect 35532 33058 35588 33068
rect 35532 32564 35588 32574
rect 35644 32564 35700 33628
rect 35588 32508 35700 32564
rect 35868 33346 35924 33358
rect 35868 33294 35870 33346
rect 35922 33294 35924 33346
rect 35868 32564 35924 33294
rect 36540 33346 36596 34076
rect 36764 34690 36820 34972
rect 36764 34638 36766 34690
rect 36818 34638 36820 34690
rect 36764 33684 36820 34638
rect 36876 34018 36932 36542
rect 38332 36708 38388 36718
rect 37884 36260 37940 36270
rect 37884 34914 37940 36204
rect 37996 36258 38052 36270
rect 37996 36206 37998 36258
rect 38050 36206 38052 36258
rect 37996 35364 38052 36206
rect 37996 35298 38052 35308
rect 37884 34862 37886 34914
rect 37938 34862 37940 34914
rect 37884 34850 37940 34862
rect 38332 35026 38388 36652
rect 38668 36372 38724 36382
rect 39116 36372 39172 36382
rect 39452 36372 39508 37436
rect 39900 37426 39956 37436
rect 40236 36706 40292 37436
rect 42028 37266 42084 37436
rect 42476 37492 42532 37502
rect 42028 37214 42030 37266
rect 42082 37214 42084 37266
rect 42028 37202 42084 37214
rect 42364 37378 42420 37390
rect 42364 37326 42366 37378
rect 42418 37326 42420 37378
rect 41692 37044 41748 37054
rect 40236 36654 40238 36706
rect 40290 36654 40292 36706
rect 40236 36642 40292 36654
rect 40572 37042 41748 37044
rect 40572 36990 41694 37042
rect 41746 36990 41748 37042
rect 40572 36988 41748 36990
rect 38668 36278 38724 36316
rect 38780 36370 39508 36372
rect 38780 36318 39118 36370
rect 39170 36318 39508 36370
rect 38780 36316 39508 36318
rect 40348 36372 40404 36382
rect 40460 36372 40516 36382
rect 40404 36370 40516 36372
rect 40404 36318 40462 36370
rect 40514 36318 40516 36370
rect 40404 36316 40516 36318
rect 38780 35586 38836 36316
rect 39116 36306 39172 36316
rect 39900 36260 39956 36270
rect 39900 36166 39956 36204
rect 40124 35810 40180 35822
rect 40124 35758 40126 35810
rect 40178 35758 40180 35810
rect 38780 35534 38782 35586
rect 38834 35534 38836 35586
rect 38780 35522 38836 35534
rect 39228 35586 39284 35598
rect 39228 35534 39230 35586
rect 39282 35534 39284 35586
rect 38332 34974 38334 35026
rect 38386 34974 38388 35026
rect 37548 34804 37604 34814
rect 37548 34710 37604 34748
rect 38332 34244 38388 34974
rect 38780 34692 38836 34702
rect 38444 34244 38500 34254
rect 38332 34242 38500 34244
rect 38332 34190 38446 34242
rect 38498 34190 38500 34242
rect 38332 34188 38500 34190
rect 38444 34178 38500 34188
rect 38556 34132 38612 34142
rect 38556 34038 38612 34076
rect 36876 33966 36878 34018
rect 36930 33966 36932 34018
rect 36876 33954 36932 33966
rect 37884 34020 37940 34030
rect 36764 33618 36820 33628
rect 37548 33906 37604 33918
rect 37548 33854 37550 33906
rect 37602 33854 37604 33906
rect 36540 33294 36542 33346
rect 36594 33294 36596 33346
rect 36540 33282 36596 33294
rect 36652 33460 36708 33470
rect 35532 32432 35588 32508
rect 35868 32498 35924 32508
rect 36652 33234 36708 33404
rect 36652 33182 36654 33234
rect 36706 33182 36708 33234
rect 36204 32450 36260 32462
rect 36204 32398 36206 32450
rect 36258 32398 36260 32450
rect 35420 32284 36036 32340
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35980 31778 36036 32284
rect 35980 31726 35982 31778
rect 36034 31726 36036 31778
rect 35980 31714 36036 31726
rect 36204 31668 36260 32398
rect 36652 31948 36708 33182
rect 37548 31948 37604 33854
rect 37660 33572 37716 33582
rect 37660 33346 37716 33516
rect 37884 33460 37940 33964
rect 38780 33684 38836 34636
rect 39228 34692 39284 35534
rect 40124 35026 40180 35758
rect 40124 34974 40126 35026
rect 40178 34974 40180 35026
rect 40124 34962 40180 34974
rect 39228 34626 39284 34636
rect 39452 34914 39508 34926
rect 39452 34862 39454 34914
rect 39506 34862 39508 34914
rect 39452 34692 39508 34862
rect 39452 34626 39508 34636
rect 39228 34468 39284 34478
rect 39228 34354 39284 34412
rect 39228 34302 39230 34354
rect 39282 34302 39284 34354
rect 38780 33618 38836 33628
rect 39116 34132 39172 34142
rect 37884 33394 37940 33404
rect 37660 33294 37662 33346
rect 37714 33294 37716 33346
rect 37660 33282 37716 33294
rect 38332 33236 38388 33246
rect 37884 33234 38388 33236
rect 37884 33182 38334 33234
rect 38386 33182 38388 33234
rect 37884 33180 38388 33182
rect 36652 31892 36932 31948
rect 37548 31892 37716 31948
rect 36876 31890 36932 31892
rect 36876 31838 36878 31890
rect 36930 31838 36932 31890
rect 36876 31826 36932 31838
rect 37660 31778 37716 31892
rect 37660 31726 37662 31778
rect 37714 31726 37716 31778
rect 37660 31714 37716 31726
rect 36316 31668 36372 31678
rect 36204 31666 36372 31668
rect 36204 31614 36318 31666
rect 36370 31614 36372 31666
rect 36204 31612 36372 31614
rect 36316 31602 36372 31612
rect 37884 31666 37940 33180
rect 38332 33170 38388 33180
rect 39116 32562 39172 34076
rect 39116 32510 39118 32562
rect 39170 32510 39172 32562
rect 39116 32498 39172 32510
rect 38332 32452 38388 32462
rect 38332 32358 38388 32396
rect 39228 32452 39284 34302
rect 39676 34020 39732 34030
rect 39676 33926 39732 33964
rect 39228 32386 39284 32396
rect 39676 32562 39732 32574
rect 39676 32510 39678 32562
rect 39730 32510 39732 32562
rect 39676 31948 39732 32510
rect 40348 32450 40404 36316
rect 40460 36306 40516 36316
rect 40460 35812 40516 35822
rect 40572 35812 40628 36988
rect 41692 36978 41748 36988
rect 42140 36932 42196 36942
rect 42140 36706 42196 36876
rect 42140 36654 42142 36706
rect 42194 36654 42196 36706
rect 42140 36642 42196 36654
rect 42364 36484 42420 37326
rect 41020 36372 41076 36382
rect 41020 36278 41076 36316
rect 42364 36370 42420 36428
rect 42364 36318 42366 36370
rect 42418 36318 42420 36370
rect 42364 36306 42420 36318
rect 42476 36372 42532 37436
rect 43372 37492 43428 37502
rect 43372 37398 43428 37436
rect 42812 37378 42868 37390
rect 42812 37326 42814 37378
rect 42866 37326 42868 37378
rect 42812 36932 42868 37326
rect 42812 36866 42868 36876
rect 40460 35810 40628 35812
rect 40460 35758 40462 35810
rect 40514 35758 40628 35810
rect 40460 35756 40628 35758
rect 41804 36258 41860 36270
rect 41804 36206 41806 36258
rect 41858 36206 41860 36258
rect 40460 35746 40516 35756
rect 41692 35700 41748 35710
rect 41804 35700 41860 36206
rect 42364 35924 42420 35934
rect 42476 35924 42532 36316
rect 42924 36484 42980 36494
rect 42924 36370 42980 36428
rect 43484 36484 43540 36494
rect 43484 36390 43540 36428
rect 42924 36318 42926 36370
rect 42978 36318 42980 36370
rect 42924 36306 42980 36318
rect 42252 35922 42532 35924
rect 42252 35870 42366 35922
rect 42418 35870 42532 35922
rect 42252 35868 42532 35870
rect 43708 35924 43764 35934
rect 41692 35698 41860 35700
rect 41692 35646 41694 35698
rect 41746 35646 41860 35698
rect 41692 35644 41860 35646
rect 41916 35810 41972 35822
rect 41916 35758 41918 35810
rect 41970 35758 41972 35810
rect 41692 35634 41748 35644
rect 40796 34692 40852 34702
rect 40796 34354 40852 34636
rect 40796 34302 40798 34354
rect 40850 34302 40852 34354
rect 40796 34290 40852 34302
rect 41692 34692 41748 34702
rect 41692 34130 41748 34636
rect 41916 34244 41972 35758
rect 42252 35026 42308 35868
rect 42364 35858 42420 35868
rect 42252 34974 42254 35026
rect 42306 34974 42308 35026
rect 42252 34962 42308 34974
rect 43708 34468 43764 35868
rect 44156 35924 44212 45614
rect 44940 45108 44996 45118
rect 44492 45106 44996 45108
rect 44492 45054 44942 45106
rect 44994 45054 44996 45106
rect 44492 45052 44996 45054
rect 44492 44996 44548 45052
rect 44940 45042 44996 45052
rect 44380 44994 44548 44996
rect 44380 44942 44494 44994
rect 44546 44942 44548 44994
rect 44380 44940 44548 44942
rect 44268 36932 44324 36942
rect 44268 35924 44324 36876
rect 44380 36820 44436 44940
rect 44492 44930 44548 44940
rect 45948 44994 46004 46732
rect 47852 46002 47908 48188
rect 47852 45950 47854 46002
rect 47906 45950 47908 46002
rect 47852 45938 47908 45950
rect 46732 45892 46788 45902
rect 46620 45890 46788 45892
rect 46620 45838 46734 45890
rect 46786 45838 46788 45890
rect 46620 45836 46788 45838
rect 46060 45778 46116 45790
rect 46060 45726 46062 45778
rect 46114 45726 46116 45778
rect 46060 45332 46116 45726
rect 46060 45266 46116 45276
rect 46620 44996 46676 45836
rect 46732 45826 46788 45836
rect 45948 44942 45950 44994
rect 46002 44942 46004 44994
rect 45948 44930 46004 44942
rect 46396 44994 46676 44996
rect 46396 44942 46622 44994
rect 46674 44942 46676 44994
rect 46396 44940 46676 44942
rect 44716 44324 44772 44334
rect 44604 44268 44716 44324
rect 44604 43708 44660 44268
rect 44716 44230 44772 44268
rect 45500 44324 45556 44334
rect 45500 44230 45556 44268
rect 44604 43652 45220 43708
rect 44716 42756 44772 42766
rect 44716 42532 44772 42700
rect 44380 36754 44436 36764
rect 44604 42530 44772 42532
rect 44604 42478 44718 42530
rect 44770 42478 44772 42530
rect 44604 42476 44772 42478
rect 44604 36708 44660 42476
rect 44716 42466 44772 42476
rect 44716 41188 44772 41198
rect 44716 41094 44772 41132
rect 44716 39394 44772 39406
rect 44716 39342 44718 39394
rect 44770 39342 44772 39394
rect 44716 38612 44772 39342
rect 44716 37492 44772 38556
rect 44716 37426 44772 37436
rect 44940 38834 44996 38846
rect 44940 38782 44942 38834
rect 44994 38782 44996 38834
rect 44940 36932 44996 38782
rect 44940 36866 44996 36876
rect 44604 36642 44660 36652
rect 44492 36482 44548 36494
rect 44492 36430 44494 36482
rect 44546 36430 44548 36482
rect 44268 35868 44436 35924
rect 44156 35858 44212 35868
rect 44268 35698 44324 35710
rect 44268 35646 44270 35698
rect 44322 35646 44324 35698
rect 43820 35588 43876 35598
rect 44268 35588 44324 35646
rect 43820 35586 44324 35588
rect 43820 35534 43822 35586
rect 43874 35534 44324 35586
rect 43820 35532 44324 35534
rect 44380 35588 44436 35868
rect 44492 35812 44548 36430
rect 44716 36258 44772 36270
rect 44716 36206 44718 36258
rect 44770 36206 44772 36258
rect 44716 36036 44772 36206
rect 44716 35980 45108 36036
rect 44492 35756 44772 35812
rect 44380 35532 44548 35588
rect 43820 35522 43876 35532
rect 43708 34402 43764 34412
rect 43820 34692 43876 34702
rect 41916 34178 41972 34188
rect 42364 34244 42420 34254
rect 42364 34150 42420 34188
rect 41692 34078 41694 34130
rect 41746 34078 41748 34130
rect 41692 34066 41748 34078
rect 43820 34132 43876 34636
rect 43820 34066 43876 34076
rect 40460 34020 40516 34030
rect 40460 33460 40516 33964
rect 40460 33366 40516 33404
rect 44044 33684 44100 33694
rect 44044 33458 44100 33628
rect 44044 33406 44046 33458
rect 44098 33406 44100 33458
rect 44044 33394 44100 33406
rect 44044 33236 44100 33246
rect 40348 32398 40350 32450
rect 40402 32398 40404 32450
rect 40348 32386 40404 32398
rect 40796 32564 40852 32574
rect 41468 32564 41524 32574
rect 40796 32562 41524 32564
rect 40796 32510 40798 32562
rect 40850 32510 41470 32562
rect 41522 32510 41524 32562
rect 40796 32508 41524 32510
rect 39676 31892 39956 31948
rect 37884 31614 37886 31666
rect 37938 31614 37940 31666
rect 37884 31602 37940 31614
rect 39900 31556 39956 31892
rect 39900 31462 39956 31500
rect 40796 31556 40852 32508
rect 41468 32498 41524 32508
rect 44044 32562 44100 33180
rect 44044 32510 44046 32562
rect 44098 32510 44100 32562
rect 44044 32498 44100 32510
rect 44268 32564 44324 35532
rect 44380 34802 44436 34814
rect 44380 34750 44382 34802
rect 44434 34750 44436 34802
rect 44380 33572 44436 34750
rect 44492 34018 44548 35532
rect 44716 35140 44772 35756
rect 45052 35810 45108 35980
rect 45052 35758 45054 35810
rect 45106 35758 45108 35810
rect 45052 35746 45108 35758
rect 44716 35074 44772 35084
rect 44716 34690 44772 34702
rect 44716 34638 44718 34690
rect 44770 34638 44772 34690
rect 44716 34244 44772 34638
rect 44716 34178 44772 34188
rect 45052 34132 45108 34142
rect 45052 34038 45108 34076
rect 44492 33966 44494 34018
rect 44546 33966 44548 34018
rect 44492 33954 44548 33966
rect 44380 33506 44436 33516
rect 45164 33460 45220 43652
rect 45500 42756 45556 42766
rect 45500 42662 45556 42700
rect 45500 41188 45556 41198
rect 45500 41094 45556 41132
rect 45500 39618 45556 39630
rect 45500 39566 45502 39618
rect 45554 39566 45556 39618
rect 45500 38612 45556 39566
rect 45500 38546 45556 38556
rect 46060 38722 46116 38734
rect 46060 38670 46062 38722
rect 46114 38670 46116 38722
rect 45724 38050 45780 38062
rect 45724 37998 45726 38050
rect 45778 37998 45780 38050
rect 45276 37154 45332 37166
rect 45276 37102 45278 37154
rect 45330 37102 45332 37154
rect 45276 35252 45332 37102
rect 45724 36932 45780 37998
rect 46060 38052 46116 38670
rect 46060 37986 46116 37996
rect 45724 36484 45780 36876
rect 45724 36418 45780 36428
rect 46172 37266 46228 37278
rect 46172 37214 46174 37266
rect 46226 37214 46228 37266
rect 45276 35186 45332 35196
rect 46172 36370 46228 37214
rect 46172 36318 46174 36370
rect 46226 36318 46228 36370
rect 46172 35588 46228 36318
rect 45948 35140 46004 35150
rect 46172 35140 46228 35532
rect 46284 35140 46340 35150
rect 46172 35138 46340 35140
rect 46172 35086 46286 35138
rect 46338 35086 46340 35138
rect 46172 35084 46340 35086
rect 45948 35046 46004 35084
rect 46284 35074 46340 35084
rect 46396 34356 46452 44940
rect 46620 44930 46676 44940
rect 46620 44210 46676 44222
rect 46620 44158 46622 44210
rect 46674 44158 46676 44210
rect 46620 43876 46676 44158
rect 46620 43810 46676 43820
rect 46620 42642 46676 42654
rect 46620 42590 46622 42642
rect 46674 42590 46676 42642
rect 46620 42420 46676 42590
rect 46620 42354 46676 42364
rect 46620 41074 46676 41086
rect 46620 41022 46622 41074
rect 46674 41022 46676 41074
rect 46620 40964 46676 41022
rect 46620 40898 46676 40908
rect 46620 39508 46676 39518
rect 46620 39414 46676 39452
rect 46620 37938 46676 37950
rect 46620 37886 46622 37938
rect 46674 37886 46676 37938
rect 46620 36596 46676 37886
rect 46620 36530 46676 36540
rect 47180 37826 47236 37838
rect 47180 37774 47182 37826
rect 47234 37774 47236 37826
rect 47180 36932 47236 37774
rect 46732 36484 46788 36494
rect 47180 36484 47236 36876
rect 46732 36482 47236 36484
rect 46732 36430 46734 36482
rect 46786 36430 47236 36482
rect 46732 36428 47236 36430
rect 46396 34290 46452 34300
rect 46508 36372 46564 36382
rect 46508 34802 46564 36316
rect 46732 35812 46788 36428
rect 47628 36372 47684 36382
rect 46732 35746 46788 35756
rect 47068 36258 47124 36270
rect 47068 36206 47070 36258
rect 47122 36206 47124 36258
rect 47068 35700 47124 36206
rect 47068 35634 47124 35644
rect 47516 35812 47572 35822
rect 47180 35588 47236 35598
rect 47180 35494 47236 35532
rect 46508 34750 46510 34802
rect 46562 34750 46564 34802
rect 45836 34244 45892 34254
rect 45836 34150 45892 34188
rect 45164 33394 45220 33404
rect 45388 34132 45444 34142
rect 44716 33348 44772 33358
rect 44716 33254 44772 33292
rect 45388 32674 45444 34076
rect 45948 33572 46004 33582
rect 45948 33478 46004 33516
rect 46284 33348 46340 33358
rect 46284 33254 46340 33292
rect 46508 33234 46564 34750
rect 46956 34802 47012 34814
rect 46956 34750 46958 34802
rect 47010 34750 47012 34802
rect 46956 34020 47012 34750
rect 46956 33348 47012 33964
rect 46956 33282 47012 33292
rect 46508 33182 46510 33234
rect 46562 33182 46564 33234
rect 46508 33170 46564 33182
rect 46844 33236 46900 33246
rect 45388 32622 45390 32674
rect 45442 32622 45444 32674
rect 45388 32610 45444 32622
rect 44604 32564 44660 32574
rect 44268 32562 44660 32564
rect 44268 32510 44606 32562
rect 44658 32510 44660 32562
rect 44268 32508 44660 32510
rect 42252 32452 42308 32462
rect 42252 32358 42308 32396
rect 42812 32452 42868 32462
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 30492 27076 30548 27086
rect 30268 27074 30548 27076
rect 30268 27022 30494 27074
rect 30546 27022 30548 27074
rect 30268 27020 30548 27022
rect 3388 26898 3444 26908
rect 6412 26964 6468 26974
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 6412 23266 6468 26908
rect 29932 26964 29988 26974
rect 30268 26964 30324 27020
rect 30492 27010 30548 27020
rect 29932 26962 30324 26964
rect 29932 26910 29934 26962
rect 29986 26910 30324 26962
rect 29932 26908 30324 26910
rect 29932 26898 29988 26908
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 6412 23214 6414 23266
rect 6466 23214 6468 23266
rect 6412 23202 6468 23214
rect 5740 23154 5796 23166
rect 5740 23102 5742 23154
rect 5794 23102 5796 23154
rect 5740 23044 5796 23102
rect 5740 22978 5796 22988
rect 8540 23042 8596 23054
rect 8540 22990 8542 23042
rect 8594 22990 8596 23042
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 8540 22484 8596 22990
rect 8988 23044 9044 23054
rect 8988 22950 9044 22988
rect 8540 22418 8596 22428
rect 10444 22484 10500 22494
rect 1820 22146 1876 22158
rect 1820 22094 1822 22146
rect 1874 22094 1876 22146
rect 1820 21924 1876 22094
rect 1820 21858 1876 21868
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 3276 16212 3332 16222
rect 3276 16210 3444 16212
rect 3276 16158 3278 16210
rect 3330 16158 3444 16210
rect 3276 16156 3444 16158
rect 3276 16146 3332 16156
rect 1932 15986 1988 15998
rect 1932 15934 1934 15986
rect 1986 15934 1988 15986
rect 1820 15764 1876 15774
rect 1932 15764 1988 15934
rect 1876 15708 1988 15764
rect 1820 15538 1876 15708
rect 1820 15486 1822 15538
rect 1874 15486 1876 15538
rect 1820 15474 1876 15486
rect 3388 13860 3444 16156
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 10444 13970 10500 22428
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 30268 20130 30324 26908
rect 33628 26964 33684 26974
rect 33628 23044 33684 26908
rect 34860 26964 34916 28476
rect 38444 28530 38500 28542
rect 38444 28478 38446 28530
rect 38498 28478 38500 28530
rect 38108 28420 38164 28430
rect 37548 28418 38164 28420
rect 37548 28366 38110 28418
rect 38162 28366 38164 28418
rect 37548 28364 38164 28366
rect 37548 27970 37604 28364
rect 38108 28354 38164 28364
rect 37548 27918 37550 27970
rect 37602 27918 37604 27970
rect 37548 27906 37604 27918
rect 36876 27860 36932 27870
rect 36876 27766 36932 27804
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 34860 26898 34916 26908
rect 37660 27074 37716 27086
rect 37660 27022 37662 27074
rect 37714 27022 37716 27074
rect 37660 26964 37716 27022
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 37660 23266 37716 26908
rect 38332 26962 38388 26974
rect 38332 26910 38334 26962
rect 38386 26910 38388 26962
rect 38332 26516 38388 26910
rect 38444 26740 38500 28478
rect 39788 28420 39844 28430
rect 39676 27748 39732 27758
rect 39788 27748 39844 28364
rect 39676 27746 39844 27748
rect 39676 27694 39678 27746
rect 39730 27694 39844 27746
rect 39676 27692 39844 27694
rect 39676 27682 39732 27692
rect 38444 26674 38500 26684
rect 38780 27076 38836 27086
rect 38444 26516 38500 26526
rect 38332 26514 38500 26516
rect 38332 26462 38446 26514
rect 38498 26462 38500 26514
rect 38332 26460 38500 26462
rect 38444 26450 38500 26460
rect 38780 26402 38836 27020
rect 39452 26740 39508 26750
rect 39452 26514 39508 26684
rect 39452 26462 39454 26514
rect 39506 26462 39508 26514
rect 39452 26450 39508 26462
rect 38780 26350 38782 26402
rect 38834 26350 38836 26402
rect 38780 26338 38836 26350
rect 39788 26290 39844 27692
rect 40124 27860 40180 27870
rect 40124 27746 40180 27804
rect 40124 27694 40126 27746
rect 40178 27694 40180 27746
rect 40124 27188 40180 27694
rect 40796 27748 40852 31500
rect 42476 31556 42532 31566
rect 42476 31462 42532 31500
rect 42588 28644 42644 28654
rect 42588 28530 42644 28588
rect 42588 28478 42590 28530
rect 42642 28478 42644 28530
rect 42588 28466 42644 28478
rect 41580 27858 41636 27870
rect 41580 27806 41582 27858
rect 41634 27806 41636 27858
rect 41580 27748 41636 27806
rect 42812 27858 42868 32396
rect 43260 32450 43316 32462
rect 43260 32398 43262 32450
rect 43314 32398 43316 32450
rect 43260 32228 43316 32398
rect 43260 32162 43316 32172
rect 43372 32452 43428 32462
rect 43372 32004 43428 32396
rect 43036 31556 43092 31566
rect 43036 31462 43092 31500
rect 43372 31218 43428 31948
rect 43932 32004 43988 32014
rect 44268 31948 44324 32508
rect 44604 32498 44660 32508
rect 43932 31892 44324 31948
rect 43372 31166 43374 31218
rect 43426 31166 43428 31218
rect 43372 31154 43428 31166
rect 43596 31778 43652 31790
rect 43596 31726 43598 31778
rect 43650 31726 43652 31778
rect 43596 30100 43652 31726
rect 43932 30994 43988 31892
rect 45724 31780 45780 31790
rect 45724 31778 46116 31780
rect 45724 31726 45726 31778
rect 45778 31726 46116 31778
rect 45724 31724 46116 31726
rect 45724 31714 45780 31724
rect 43932 30942 43934 30994
rect 43986 30942 43988 30994
rect 43932 30930 43988 30942
rect 44380 31666 44436 31678
rect 44380 31614 44382 31666
rect 44434 31614 44436 31666
rect 43596 30034 43652 30044
rect 44044 30322 44100 30334
rect 44044 30270 44046 30322
rect 44098 30270 44100 30322
rect 43260 29428 43316 29438
rect 43260 29314 43316 29372
rect 43820 29428 43876 29438
rect 43820 29334 43876 29372
rect 43260 29262 43262 29314
rect 43314 29262 43316 29314
rect 43260 28532 43316 29262
rect 44044 29316 44100 30270
rect 44380 30212 44436 31614
rect 44716 31554 44772 31566
rect 44716 31502 44718 31554
rect 44770 31502 44772 31554
rect 44716 31106 44772 31502
rect 44716 31054 44718 31106
rect 44770 31054 44772 31106
rect 44716 31042 44772 31054
rect 44380 30146 44436 30156
rect 44716 30210 44772 30222
rect 44716 30158 44718 30210
rect 44770 30158 44772 30210
rect 44716 29540 44772 30158
rect 45836 30212 45892 30222
rect 45836 30118 45892 30156
rect 46060 30212 46116 31724
rect 46620 31666 46676 31678
rect 46620 31614 46622 31666
rect 46674 31614 46676 31666
rect 46620 30772 46676 31614
rect 46844 30884 46900 33180
rect 47516 32450 47572 35756
rect 47516 32398 47518 32450
rect 47570 32398 47572 32450
rect 47516 32386 47572 32398
rect 47628 35026 47684 36316
rect 48076 36258 48132 36270
rect 48076 36206 48078 36258
rect 48130 36206 48132 36258
rect 47628 34974 47630 35026
rect 47682 34974 47684 35026
rect 47628 33458 47684 34974
rect 47740 35810 47796 35822
rect 47740 35758 47742 35810
rect 47794 35758 47796 35810
rect 47740 34132 47796 35758
rect 48076 35812 48132 36206
rect 48076 35746 48132 35756
rect 47964 35700 48020 35710
rect 47964 35606 48020 35644
rect 47740 34066 47796 34076
rect 47964 34020 48020 34030
rect 47964 33926 48020 33964
rect 47628 33406 47630 33458
rect 47682 33406 47684 33458
rect 47628 31948 47684 33406
rect 46620 30706 46676 30716
rect 46732 30882 46900 30884
rect 46732 30830 46846 30882
rect 46898 30830 46900 30882
rect 46732 30828 46900 30830
rect 46732 30548 46788 30828
rect 46844 30818 46900 30828
rect 47516 31892 47684 31948
rect 46172 30492 46788 30548
rect 46172 30434 46228 30492
rect 46172 30382 46174 30434
rect 46226 30382 46228 30434
rect 46172 30370 46228 30382
rect 46284 30268 46788 30324
rect 46284 30212 46340 30268
rect 46060 30156 46340 30212
rect 44716 29474 44772 29484
rect 44044 29250 44100 29260
rect 44604 29316 44660 29326
rect 44604 29314 44772 29316
rect 44604 29262 44606 29314
rect 44658 29262 44772 29314
rect 44604 29260 44772 29262
rect 44604 29250 44660 29260
rect 43260 28466 43316 28476
rect 43484 28642 43540 28654
rect 43484 28590 43486 28642
rect 43538 28590 43540 28642
rect 42924 28420 42980 28430
rect 43484 28420 43540 28590
rect 42924 28418 43204 28420
rect 42924 28366 42926 28418
rect 42978 28366 43204 28418
rect 42924 28364 43204 28366
rect 42924 28354 42980 28364
rect 43148 28084 43204 28364
rect 43484 28354 43540 28364
rect 44604 28530 44660 28542
rect 44604 28478 44606 28530
rect 44658 28478 44660 28530
rect 43148 28028 43652 28084
rect 43596 27970 43652 28028
rect 43596 27918 43598 27970
rect 43650 27918 43652 27970
rect 43596 27906 43652 27918
rect 42812 27806 42814 27858
rect 42866 27806 42868 27858
rect 40796 27746 41636 27748
rect 40796 27694 40798 27746
rect 40850 27694 41636 27746
rect 40796 27692 41636 27694
rect 42028 27746 42084 27758
rect 42028 27694 42030 27746
rect 42082 27694 42084 27746
rect 40124 27122 40180 27132
rect 40236 27300 40292 27310
rect 39788 26238 39790 26290
rect 39842 26238 39844 26290
rect 39788 26226 39844 26238
rect 40236 26290 40292 27244
rect 40460 27186 40516 27198
rect 40460 27134 40462 27186
rect 40514 27134 40516 27186
rect 40460 26852 40516 27134
rect 40516 26796 40628 26852
rect 40460 26786 40516 26796
rect 40572 26402 40628 26796
rect 40572 26350 40574 26402
rect 40626 26350 40628 26402
rect 40572 26338 40628 26350
rect 40236 26238 40238 26290
rect 40290 26238 40292 26290
rect 40236 26226 40292 26238
rect 40460 23380 40516 23390
rect 40796 23380 40852 27692
rect 41692 27300 41748 27310
rect 41580 27188 41636 27198
rect 41132 27076 41188 27086
rect 41132 26982 41188 27020
rect 41468 27074 41524 27086
rect 41468 27022 41470 27074
rect 41522 27022 41524 27074
rect 41468 26852 41524 27022
rect 41468 26786 41524 26796
rect 41580 26292 41636 27132
rect 41692 26962 41748 27244
rect 42028 27300 42084 27694
rect 42028 27234 42084 27244
rect 42812 27188 42868 27806
rect 44604 27860 44660 28478
rect 44716 28084 44772 29260
rect 45948 28868 46004 28878
rect 46060 28868 46116 30156
rect 46396 30100 46452 30110
rect 46396 30006 46452 30044
rect 46732 30098 46788 30268
rect 46732 30046 46734 30098
rect 46786 30046 46788 30098
rect 46732 30034 46788 30046
rect 47516 30100 47572 31892
rect 47516 30006 47572 30044
rect 45724 28866 46116 28868
rect 45724 28814 45950 28866
rect 46002 28814 46116 28866
rect 45724 28812 46116 28814
rect 46732 29540 46788 29550
rect 46732 29314 46788 29484
rect 46732 29262 46734 29314
rect 46786 29262 46788 29314
rect 45612 28644 45668 28654
rect 45612 28550 45668 28588
rect 44716 28018 44772 28028
rect 45612 28308 45668 28318
rect 44604 27794 44660 27804
rect 43260 27188 43316 27198
rect 42868 27186 43316 27188
rect 42868 27134 43262 27186
rect 43314 27134 43316 27186
rect 42868 27132 43316 27134
rect 41692 26910 41694 26962
rect 41746 26910 41748 26962
rect 41692 26898 41748 26910
rect 42140 27076 42196 27086
rect 42812 27056 42868 27132
rect 42140 26962 42196 27020
rect 42140 26910 42142 26962
rect 42194 26910 42196 26962
rect 42140 26898 42196 26910
rect 42252 26964 42308 26974
rect 41244 26290 41636 26292
rect 41244 26238 41582 26290
rect 41634 26238 41636 26290
rect 41244 26236 41636 26238
rect 41244 25618 41300 26236
rect 41580 26226 41636 26236
rect 41244 25566 41246 25618
rect 41298 25566 41300 25618
rect 41244 25554 41300 25566
rect 40460 23378 40852 23380
rect 40460 23326 40462 23378
rect 40514 23326 40852 23378
rect 40460 23324 40852 23326
rect 42252 23378 42308 26908
rect 42364 26180 42420 26190
rect 42364 26178 42644 26180
rect 42364 26126 42366 26178
rect 42418 26126 42644 26178
rect 42364 26124 42644 26126
rect 42364 26114 42420 26124
rect 42588 25394 42644 26124
rect 42588 25342 42590 25394
rect 42642 25342 42644 25394
rect 42588 25330 42644 25342
rect 42924 25396 42980 25406
rect 42924 25394 43204 25396
rect 42924 25342 42926 25394
rect 42978 25342 43204 25394
rect 42924 25340 43204 25342
rect 42924 25330 42980 25340
rect 43148 24500 43204 25340
rect 43260 24836 43316 27132
rect 43820 26964 43876 26974
rect 43260 24780 43764 24836
rect 43148 24444 43540 24500
rect 43484 24162 43540 24444
rect 43708 24498 43764 24780
rect 43708 24446 43710 24498
rect 43762 24446 43764 24498
rect 43708 24434 43764 24446
rect 43484 24110 43486 24162
rect 43538 24110 43540 24162
rect 43484 24098 43540 24110
rect 43820 24162 43876 26908
rect 44492 26964 44548 26974
rect 44492 26178 44548 26908
rect 45500 26964 45556 26974
rect 45052 26852 45108 26862
rect 45052 26290 45108 26796
rect 45052 26238 45054 26290
rect 45106 26238 45108 26290
rect 45052 26226 45108 26238
rect 44492 26126 44494 26178
rect 44546 26126 44548 26178
rect 44492 26114 44548 26126
rect 44492 25506 44548 25518
rect 44492 25454 44494 25506
rect 44546 25454 44548 25506
rect 44492 24836 44548 25454
rect 45500 25506 45556 26908
rect 45612 26962 45668 28252
rect 45724 27746 45780 28812
rect 45948 28802 46004 28812
rect 45724 27694 45726 27746
rect 45778 27694 45780 27746
rect 45724 27682 45780 27694
rect 46172 28530 46228 28542
rect 46732 28532 46788 29262
rect 46172 28478 46174 28530
rect 46226 28478 46228 28530
rect 45612 26910 45614 26962
rect 45666 26910 45668 26962
rect 45612 26898 45668 26910
rect 46172 27300 46228 28478
rect 46396 28530 46788 28532
rect 46396 28478 46734 28530
rect 46786 28478 46788 28530
rect 46396 28476 46788 28478
rect 46284 28084 46340 28094
rect 46284 27990 46340 28028
rect 46172 26962 46228 27244
rect 46396 27298 46452 28476
rect 46732 28466 46788 28476
rect 46396 27246 46398 27298
rect 46450 27246 46452 27298
rect 46396 27234 46452 27246
rect 46620 27858 46676 27870
rect 46620 27806 46622 27858
rect 46674 27806 46676 27858
rect 46620 27300 46676 27806
rect 46732 27300 46788 27310
rect 46620 27298 46788 27300
rect 46620 27246 46734 27298
rect 46786 27246 46788 27298
rect 46620 27244 46788 27246
rect 46732 27234 46788 27244
rect 46172 26910 46174 26962
rect 46226 26910 46228 26962
rect 46172 26898 46228 26910
rect 46172 26404 46228 26414
rect 46172 26310 46228 26348
rect 45500 25454 45502 25506
rect 45554 25454 45556 25506
rect 45500 25442 45556 25454
rect 46620 25394 46676 25406
rect 46620 25342 46622 25394
rect 46674 25342 46676 25394
rect 44716 25284 44772 25294
rect 44716 25282 45332 25284
rect 44716 25230 44718 25282
rect 44770 25230 45332 25282
rect 44716 25228 45332 25230
rect 44716 25218 44772 25228
rect 44492 24770 44548 24780
rect 45276 24834 45332 25228
rect 46620 24948 46676 25342
rect 46620 24882 46676 24892
rect 45276 24782 45278 24834
rect 45330 24782 45332 24834
rect 45276 24770 45332 24782
rect 45948 24836 46004 24846
rect 44604 24722 44660 24734
rect 44604 24670 44606 24722
rect 44658 24670 44660 24722
rect 43932 24612 43988 24622
rect 44604 24612 44660 24670
rect 43932 24610 44660 24612
rect 43932 24558 43934 24610
rect 43986 24558 44660 24610
rect 43932 24556 44660 24558
rect 43932 24498 43988 24556
rect 43932 24446 43934 24498
rect 43986 24446 43988 24498
rect 43932 24434 43988 24446
rect 43820 24110 43822 24162
rect 43874 24110 43876 24162
rect 43820 24098 43876 24110
rect 44380 23938 44436 23950
rect 44380 23886 44382 23938
rect 44434 23886 44436 23938
rect 42252 23326 42254 23378
rect 42306 23326 42308 23378
rect 40460 23314 40516 23324
rect 37660 23214 37662 23266
rect 37714 23214 37716 23266
rect 37660 23202 37716 23214
rect 42252 23268 42308 23326
rect 43932 23828 43988 23838
rect 42252 23202 42308 23212
rect 43596 23268 43652 23278
rect 33628 22978 33684 22988
rect 33740 23156 33796 23166
rect 34300 23156 34356 23166
rect 33740 23154 34356 23156
rect 33740 23102 33742 23154
rect 33794 23102 34302 23154
rect 34354 23102 34356 23154
rect 33740 23100 34356 23102
rect 30268 20078 30270 20130
rect 30322 20078 30324 20130
rect 26796 20020 26852 20030
rect 26348 20018 26852 20020
rect 26348 19966 26798 20018
rect 26850 19966 26852 20018
rect 26348 19964 26852 19966
rect 26348 19908 26404 19964
rect 26796 19954 26852 19964
rect 26236 19906 26404 19908
rect 26236 19854 26350 19906
rect 26402 19854 26404 19906
rect 26236 19852 26404 19854
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 21980 15426 22036 15438
rect 21980 15374 21982 15426
rect 22034 15374 22036 15426
rect 21420 15316 21476 15326
rect 21084 15314 21476 15316
rect 21084 15262 21422 15314
rect 21474 15262 21476 15314
rect 21084 15260 21476 15262
rect 20300 15202 20356 15214
rect 20300 15150 20302 15202
rect 20354 15150 20356 15202
rect 20188 15092 20244 15102
rect 19964 14642 20020 14654
rect 19964 14590 19966 14642
rect 20018 14590 20020 14642
rect 10444 13918 10446 13970
rect 10498 13918 10500 13970
rect 3388 13794 3444 13804
rect 6860 13860 6916 13870
rect 6860 13766 6916 13804
rect 10444 13860 10500 13918
rect 17052 14530 17108 14542
rect 17052 14478 17054 14530
rect 17106 14478 17108 14530
rect 10444 13794 10500 13804
rect 11788 13860 11844 13870
rect 11788 13766 11844 13804
rect 6188 13748 6244 13758
rect 6188 13654 6244 13692
rect 9660 13748 9716 13758
rect 8988 13634 9044 13646
rect 8988 13582 8990 13634
rect 9042 13582 9044 13634
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 8988 12292 9044 13582
rect 8988 12226 9044 12236
rect 9660 13634 9716 13692
rect 11004 13748 11060 13758
rect 11004 13654 11060 13692
rect 13468 13748 13524 13758
rect 9660 13582 9662 13634
rect 9714 13582 9716 13634
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 1820 9604 1876 9614
rect 1820 9510 1876 9548
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 9660 8428 9716 13582
rect 13468 12178 13524 13692
rect 14364 13748 14420 13758
rect 14364 13654 14420 13692
rect 16716 13748 16772 13758
rect 13916 13636 13972 13646
rect 13916 13542 13972 13580
rect 16716 12402 16772 13692
rect 17052 13748 17108 14478
rect 17052 13682 17108 13692
rect 17836 14532 17892 14542
rect 17836 14418 17892 14476
rect 17836 14366 17838 14418
rect 17890 14366 17892 14418
rect 17836 13636 17892 14366
rect 19964 14420 20020 14590
rect 19964 14354 20020 14364
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 20188 13858 20244 15036
rect 20188 13806 20190 13858
rect 20242 13806 20244 13858
rect 19404 13748 19460 13758
rect 19404 13654 19460 13692
rect 17836 13570 17892 13580
rect 18844 13636 18900 13646
rect 16716 12350 16718 12402
rect 16770 12350 16772 12402
rect 16716 12338 16772 12350
rect 14140 12292 14196 12302
rect 14140 12198 14196 12236
rect 13468 12126 13470 12178
rect 13522 12126 13524 12178
rect 13468 12114 13524 12126
rect 16268 12068 16324 12078
rect 16268 11974 16324 12012
rect 9212 8372 9716 8428
rect 16604 8372 16660 8382
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 3388 5236 3444 5246
rect 1820 4228 1876 4238
rect 2940 4228 2996 4238
rect 1820 4226 1988 4228
rect 1820 4174 1822 4226
rect 1874 4174 1988 4226
rect 1820 4172 1988 4174
rect 1820 4162 1876 4172
rect 1932 3444 1988 4172
rect 1932 3350 1988 3388
rect 2940 800 2996 4172
rect 3276 3668 3332 3678
rect 3388 3668 3444 5180
rect 6524 5236 6580 5246
rect 6524 5142 6580 5180
rect 8652 5234 8708 5246
rect 8652 5182 8654 5234
rect 8706 5182 8708 5234
rect 5852 5124 5908 5134
rect 5852 5030 5908 5068
rect 8652 5012 8708 5182
rect 9212 5234 9268 8372
rect 16604 8278 16660 8316
rect 18844 8372 18900 13580
rect 20188 13636 20244 13806
rect 20300 13748 20356 15150
rect 20972 15202 21028 15214
rect 20972 15150 20974 15202
rect 21026 15150 21028 15202
rect 20972 15092 21028 15150
rect 20972 15026 21028 15036
rect 20524 14532 20580 14542
rect 20524 14438 20580 14476
rect 20860 14532 20916 14542
rect 21084 14532 21140 15260
rect 21420 15250 21476 15260
rect 21756 15314 21812 15326
rect 21756 15262 21758 15314
rect 21810 15262 21812 15314
rect 21756 15092 21812 15262
rect 21756 15026 21812 15036
rect 21980 14756 22036 15374
rect 22092 15204 22148 15214
rect 22092 15110 22148 15148
rect 22092 14756 22148 14766
rect 21980 14754 22148 14756
rect 21980 14702 22094 14754
rect 22146 14702 22148 14754
rect 21980 14700 22148 14702
rect 22092 14690 22148 14700
rect 20860 14530 21140 14532
rect 20860 14478 20862 14530
rect 20914 14478 21140 14530
rect 20860 14476 21140 14478
rect 20860 14466 20916 14476
rect 20636 14420 20692 14430
rect 20636 14326 20692 14364
rect 22204 14418 22260 14430
rect 22204 14366 22206 14418
rect 22258 14366 22260 14418
rect 20300 13682 20356 13692
rect 20188 13570 20244 13580
rect 21644 13636 21700 13646
rect 22204 13636 22260 14366
rect 22316 13636 22372 13646
rect 22204 13634 22372 13636
rect 22204 13582 22318 13634
rect 22370 13582 22372 13634
rect 22204 13580 22372 13582
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 21532 12068 21588 12078
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 18844 8306 18900 8316
rect 13804 8260 13860 8270
rect 13804 8166 13860 8204
rect 17052 8260 17108 8270
rect 17052 8166 17108 8204
rect 9212 5182 9214 5234
rect 9266 5182 9268 5234
rect 9212 5124 9268 5182
rect 9212 5058 9268 5068
rect 14476 8146 14532 8158
rect 14476 8094 14478 8146
rect 14530 8094 14532 8146
rect 8652 4946 8708 4956
rect 14476 5012 14532 8094
rect 21532 8148 21588 12012
rect 21532 8082 21588 8092
rect 21644 12066 21700 13580
rect 22316 13570 22372 13580
rect 22764 13636 22820 13646
rect 22764 13542 22820 13580
rect 24444 12180 24500 12190
rect 24444 12086 24500 12124
rect 24892 12180 24948 12190
rect 24892 12086 24948 12124
rect 21644 12014 21646 12066
rect 21698 12014 21700 12066
rect 21644 8260 21700 12014
rect 25228 8372 25284 8382
rect 25788 8372 25844 8382
rect 25228 8370 25844 8372
rect 25228 8318 25230 8370
rect 25282 8318 25790 8370
rect 25842 8318 25844 8370
rect 25228 8316 25844 8318
rect 25228 8306 25284 8316
rect 25788 8306 25844 8316
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 21644 7700 21700 8204
rect 22316 8260 22372 8270
rect 22316 8166 22372 8204
rect 26012 8258 26068 8270
rect 26012 8206 26014 8258
rect 26066 8206 26068 8258
rect 21756 8148 21812 8158
rect 21756 8054 21812 8092
rect 23100 8148 23156 8158
rect 23100 8054 23156 8092
rect 26012 8148 26068 8206
rect 21756 7700 21812 7710
rect 21644 7698 21812 7700
rect 21644 7646 21758 7698
rect 21810 7646 21812 7698
rect 21644 7644 21812 7646
rect 21756 7634 21812 7644
rect 25676 7700 25732 7710
rect 26012 7700 26068 8092
rect 25676 7698 26068 7700
rect 25676 7646 25678 7698
rect 25730 7646 26068 7698
rect 25676 7644 26068 7646
rect 25676 7634 25732 7644
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 14476 4946 14532 4956
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 26236 4228 26292 19852
rect 26348 19842 26404 19852
rect 30268 19908 30324 20078
rect 30268 19842 30324 19852
rect 33740 19908 33796 23100
rect 34300 23090 34356 23100
rect 40124 23154 40180 23166
rect 40124 23102 40126 23154
rect 40178 23102 40180 23154
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 39788 22148 39844 22158
rect 40124 22148 40180 23102
rect 43372 23042 43428 23054
rect 43372 22990 43374 23042
rect 43426 22990 43428 23042
rect 43372 22932 43428 22990
rect 43372 22866 43428 22876
rect 39788 22146 40180 22148
rect 39788 22094 39790 22146
rect 39842 22094 40180 22146
rect 39788 22092 40180 22094
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 33740 12402 33796 19852
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 38780 17668 38836 17678
rect 38780 17106 38836 17612
rect 38780 17054 38782 17106
rect 38834 17054 38836 17106
rect 38780 17042 38836 17054
rect 37884 16884 37940 16894
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 37884 15204 37940 16828
rect 38444 16884 38500 16894
rect 38444 16790 38500 16828
rect 39788 16884 39844 22092
rect 43596 21924 43652 23212
rect 43932 23154 43988 23772
rect 43932 23102 43934 23154
rect 43986 23102 43988 23154
rect 43932 23090 43988 23102
rect 44044 22482 44100 22494
rect 44044 22430 44046 22482
rect 44098 22430 44100 22482
rect 44044 22036 44100 22430
rect 44044 21970 44100 21980
rect 43372 21868 43596 21924
rect 43372 21810 43428 21868
rect 43596 21858 43652 21868
rect 43932 21924 43988 21934
rect 43372 21758 43374 21810
rect 43426 21758 43428 21810
rect 42476 20020 42532 20030
rect 39788 16818 39844 16828
rect 40236 17668 40292 17678
rect 37884 15138 37940 15148
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 33740 12350 33742 12402
rect 33794 12350 33796 12402
rect 33740 12180 33796 12350
rect 39340 12292 39396 12302
rect 39340 12198 39396 12236
rect 33740 12114 33796 12124
rect 34300 12180 34356 12190
rect 34300 12086 34356 12124
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 39116 10722 39172 10734
rect 39116 10670 39118 10722
rect 39170 10670 39172 10722
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 39004 9940 39060 9950
rect 39116 9940 39172 10670
rect 39004 9938 39172 9940
rect 39004 9886 39006 9938
rect 39058 9886 39172 9938
rect 39004 9884 39172 9886
rect 39452 10610 39508 10622
rect 39452 10558 39454 10610
rect 39506 10558 39508 10610
rect 39004 9874 39060 9884
rect 38220 9826 38276 9838
rect 38220 9774 38222 9826
rect 38274 9774 38276 9826
rect 37660 9604 37716 9614
rect 38220 9604 38276 9774
rect 37660 9602 38276 9604
rect 37660 9550 37662 9602
rect 37714 9550 38276 9602
rect 37660 9548 38276 9550
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 26348 8036 26404 8046
rect 26348 7942 26404 7980
rect 34860 8036 34916 8046
rect 34860 6690 34916 7980
rect 37324 7476 37380 7486
rect 37324 7382 37380 7420
rect 37660 7476 37716 9548
rect 39116 9268 39172 9278
rect 39116 9174 39172 9212
rect 38668 8930 38724 8942
rect 38668 8878 38670 8930
rect 38722 8878 38724 8930
rect 38332 8148 38388 8158
rect 38332 8146 38612 8148
rect 38332 8094 38334 8146
rect 38386 8094 38612 8146
rect 38332 8092 38612 8094
rect 38332 8082 38388 8092
rect 37996 8034 38052 8046
rect 37996 7982 37998 8034
rect 38050 7982 38052 8034
rect 37996 7586 38052 7982
rect 37996 7534 37998 7586
rect 38050 7534 38052 7586
rect 37996 7522 38052 7534
rect 37660 7410 37716 7420
rect 38332 7476 38388 7486
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 34860 6638 34862 6690
rect 34914 6638 34916 6690
rect 34860 6580 34916 6638
rect 34860 6514 34916 6524
rect 35868 6690 35924 6702
rect 35868 6638 35870 6690
rect 35922 6638 35924 6690
rect 35532 6466 35588 6478
rect 35532 6414 35534 6466
rect 35586 6414 35588 6466
rect 35084 6020 35140 6030
rect 34636 6018 35140 6020
rect 34636 5966 35086 6018
rect 35138 5966 35140 6018
rect 34636 5964 35140 5966
rect 33964 5236 34020 5246
rect 33964 5122 34020 5180
rect 34636 5234 34692 5964
rect 35084 5954 35140 5964
rect 35420 6020 35476 6030
rect 35532 6020 35588 6414
rect 35420 6018 35588 6020
rect 35420 5966 35422 6018
rect 35474 5966 35588 6018
rect 35420 5964 35588 5966
rect 35420 5954 35476 5964
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 34636 5182 34638 5234
rect 34690 5182 34692 5234
rect 34636 5170 34692 5182
rect 35532 5236 35588 5246
rect 33964 5070 33966 5122
rect 34018 5070 34020 5122
rect 33964 5058 34020 5070
rect 35532 4338 35588 5180
rect 35868 5012 35924 6638
rect 36652 6692 36708 6702
rect 36652 6598 36708 6636
rect 37324 6692 37380 6702
rect 36428 6580 36484 6590
rect 36428 6486 36484 6524
rect 35868 4946 35924 4956
rect 36764 6018 36820 6030
rect 36764 5966 36766 6018
rect 36818 5966 36820 6018
rect 36764 5234 36820 5966
rect 37324 6018 37380 6636
rect 37324 5966 37326 6018
rect 37378 5966 37380 6018
rect 37324 5954 37380 5966
rect 37436 6466 37492 6478
rect 37436 6414 37438 6466
rect 37490 6414 37492 6466
rect 36764 5182 36766 5234
rect 36818 5182 36820 5234
rect 36764 5012 36820 5182
rect 36764 4946 36820 4956
rect 37436 5012 37492 6414
rect 37548 5908 37604 5918
rect 37548 5814 37604 5852
rect 38220 5908 38276 5918
rect 37884 5682 37940 5694
rect 37884 5630 37886 5682
rect 37938 5630 37940 5682
rect 37884 5122 37940 5630
rect 37884 5070 37886 5122
rect 37938 5070 37940 5122
rect 37884 5058 37940 5070
rect 37436 4946 37492 4956
rect 37548 4898 37604 4910
rect 37548 4846 37550 4898
rect 37602 4846 37604 4898
rect 36204 4452 36260 4462
rect 36204 4358 36260 4396
rect 37548 4452 37604 4846
rect 37548 4386 37604 4396
rect 35532 4286 35534 4338
rect 35586 4286 35588 4338
rect 35532 4274 35588 4286
rect 38220 4228 38276 5852
rect 38332 5236 38388 7420
rect 38556 6914 38612 8092
rect 38556 6862 38558 6914
rect 38610 6862 38612 6914
rect 38556 6850 38612 6862
rect 38668 6692 38724 8878
rect 39452 8370 39508 10558
rect 39676 9940 39732 9950
rect 39676 9268 39732 9884
rect 40236 9940 40292 17612
rect 41804 17668 41860 17678
rect 41804 17574 41860 17612
rect 42476 17668 42532 19964
rect 43260 20020 43316 20030
rect 43260 19926 43316 19964
rect 43148 18452 43204 18462
rect 43148 18358 43204 18396
rect 43372 18452 43428 21758
rect 43932 21586 43988 21868
rect 43932 21534 43934 21586
rect 43986 21534 43988 21586
rect 43932 21522 43988 21534
rect 44380 20692 44436 23886
rect 44492 23828 44548 23838
rect 44492 23734 44548 23772
rect 44604 23268 44660 24556
rect 45948 24162 46004 24780
rect 45948 24110 45950 24162
rect 46002 24110 46004 24162
rect 45948 24098 46004 24110
rect 46284 24612 46340 24622
rect 46284 24162 46340 24556
rect 47404 24612 47460 24622
rect 47404 24518 47460 24556
rect 46284 24110 46286 24162
rect 46338 24110 46340 24162
rect 46284 23828 46340 24110
rect 46284 23762 46340 23772
rect 46508 23826 46564 23838
rect 46508 23774 46510 23826
rect 46562 23774 46564 23826
rect 44604 23154 44660 23212
rect 44604 23102 44606 23154
rect 44658 23102 44660 23154
rect 44604 23090 44660 23102
rect 45948 23604 46004 23614
rect 45388 23042 45444 23054
rect 45388 22990 45390 23042
rect 45442 22990 45444 23042
rect 44716 22372 44772 22382
rect 44716 22278 44772 22316
rect 45388 22148 45444 22990
rect 45388 22082 45444 22092
rect 45948 22370 46004 23548
rect 46508 23604 46564 23774
rect 46508 23538 46564 23548
rect 46844 23826 46900 23838
rect 46844 23774 46846 23826
rect 46898 23774 46900 23826
rect 45948 22318 45950 22370
rect 46002 22318 46004 22370
rect 44716 21474 44772 21486
rect 44716 21422 44718 21474
rect 44770 21422 44772 21474
rect 44492 20804 44548 20814
rect 44492 20710 44548 20748
rect 43820 20020 43876 20030
rect 43820 19926 43876 19964
rect 44380 20018 44436 20636
rect 44716 20690 44772 21422
rect 45836 20804 45892 20814
rect 45836 20710 45892 20748
rect 44716 20638 44718 20690
rect 44770 20638 44772 20690
rect 44716 20626 44772 20638
rect 45948 20692 46004 22318
rect 46732 23044 46788 23054
rect 46844 23044 46900 23774
rect 46788 22988 46900 23044
rect 47516 23044 47572 23054
rect 46732 22372 46788 22988
rect 47516 22950 47572 22988
rect 46732 22278 46788 22316
rect 47068 22372 47124 22382
rect 47964 22372 48020 22382
rect 47068 22370 48020 22372
rect 47068 22318 47070 22370
rect 47122 22318 47966 22370
rect 48018 22318 48020 22370
rect 47068 22316 48020 22318
rect 47068 22306 47124 22316
rect 47964 22306 48020 22316
rect 45948 20626 46004 20636
rect 46172 22258 46228 22270
rect 46172 22206 46174 22258
rect 46226 22206 46228 22258
rect 46172 21476 46228 22206
rect 47740 22148 47796 22158
rect 47740 22054 47796 22092
rect 46844 21476 46900 21486
rect 46172 21474 46900 21476
rect 46172 21422 46846 21474
rect 46898 21422 46900 21474
rect 46172 21420 46900 21422
rect 46172 21026 46228 21420
rect 46844 21410 46900 21420
rect 46172 20974 46174 21026
rect 46226 20974 46228 21026
rect 44380 19966 44382 20018
rect 44434 19966 44436 20018
rect 44380 19954 44436 19966
rect 45276 20580 45332 20590
rect 45276 19906 45332 20524
rect 46172 20018 46228 20974
rect 46396 20692 46452 20702
rect 46396 20598 46452 20636
rect 46732 20690 46788 20702
rect 46732 20638 46734 20690
rect 46786 20638 46788 20690
rect 46732 20188 46788 20638
rect 46172 19966 46174 20018
rect 46226 19966 46228 20018
rect 46172 19954 46228 19966
rect 46284 20132 46788 20188
rect 45276 19854 45278 19906
rect 45330 19854 45332 19906
rect 45276 19842 45332 19854
rect 45724 19236 45780 19246
rect 46284 19236 46340 20132
rect 45724 19234 46564 19236
rect 45724 19182 45726 19234
rect 45778 19182 46564 19234
rect 45724 19180 46564 19182
rect 45724 19170 45780 19180
rect 44716 19122 44772 19134
rect 44716 19070 44718 19122
rect 44770 19070 44772 19122
rect 44380 19010 44436 19022
rect 44380 18958 44382 19010
rect 44434 18958 44436 19010
rect 44380 18564 44436 18958
rect 44492 18564 44548 18574
rect 44380 18562 44548 18564
rect 44380 18510 44494 18562
rect 44546 18510 44548 18562
rect 44380 18508 44548 18510
rect 44492 18498 44548 18508
rect 43372 18386 43428 18396
rect 43708 18452 43764 18462
rect 43708 18358 43764 18396
rect 44716 17892 44772 19070
rect 44716 17826 44772 17836
rect 45612 17892 45668 17902
rect 45612 17798 45668 17836
rect 45948 17890 46004 19180
rect 46508 18340 46564 19180
rect 46620 19124 46676 19134
rect 46620 19030 46676 19068
rect 46620 18340 46676 18350
rect 46508 18338 46676 18340
rect 46508 18286 46622 18338
rect 46674 18286 46676 18338
rect 46508 18284 46676 18286
rect 46620 18274 46676 18284
rect 45948 17838 45950 17890
rect 46002 17838 46004 17890
rect 45948 17826 46004 17838
rect 42924 17780 42980 17790
rect 42924 17686 42980 17724
rect 45052 17780 45108 17790
rect 42476 17536 42532 17612
rect 43708 17668 43764 17678
rect 44604 17668 44660 17678
rect 43708 17666 44212 17668
rect 43708 17614 43710 17666
rect 43762 17614 44212 17666
rect 43708 17612 44212 17614
rect 43708 17602 43764 17612
rect 44156 17556 44212 17612
rect 44604 17574 44660 17612
rect 41244 16884 41300 16894
rect 41244 16098 41300 16828
rect 43596 16882 43652 16894
rect 43596 16830 43598 16882
rect 43650 16830 43652 16882
rect 41244 16046 41246 16098
rect 41298 16046 41300 16098
rect 40572 15876 40628 15886
rect 41244 15876 41300 16046
rect 42924 16770 42980 16782
rect 42924 16718 42926 16770
rect 42978 16718 42980 16770
rect 40572 15874 41300 15876
rect 40572 15822 40574 15874
rect 40626 15822 41300 15874
rect 40572 15820 41300 15822
rect 40572 15810 40628 15820
rect 41244 14308 41300 15820
rect 41916 15986 41972 15998
rect 41916 15934 41918 15986
rect 41970 15934 41972 15986
rect 41916 15540 41972 15934
rect 41916 15474 41972 15484
rect 42476 15540 42532 15550
rect 42476 15446 42532 15484
rect 42924 15540 42980 16718
rect 43596 16324 43652 16830
rect 44156 16770 44212 17500
rect 44156 16718 44158 16770
rect 44210 16718 44212 16770
rect 44156 16706 44212 16718
rect 44492 16884 44548 16894
rect 43596 16268 44100 16324
rect 42924 15474 42980 15484
rect 44044 16210 44100 16268
rect 44044 16158 44046 16210
rect 44098 16158 44100 16210
rect 44044 15428 44100 16158
rect 44492 16210 44548 16828
rect 44492 16158 44494 16210
rect 44546 16158 44548 16210
rect 44492 16146 44548 16158
rect 44044 15362 44100 15372
rect 44716 15988 44772 15998
rect 44716 15428 44772 15932
rect 42812 15316 42868 15326
rect 42812 15222 42868 15260
rect 44380 15316 44436 15326
rect 44380 15222 44436 15260
rect 44716 15314 44772 15372
rect 45052 15426 45108 17724
rect 46172 17780 46228 17790
rect 46172 17554 46228 17724
rect 46172 17502 46174 17554
rect 46226 17502 46228 17554
rect 45612 15988 45668 15998
rect 45612 15894 45668 15932
rect 46172 15988 46228 17502
rect 46508 17556 46564 17566
rect 46284 16996 46340 17006
rect 46284 16902 46340 16940
rect 46396 16324 46452 16334
rect 46508 16324 46564 17500
rect 46396 16322 46564 16324
rect 46396 16270 46398 16322
rect 46450 16270 46564 16322
rect 46396 16268 46564 16270
rect 46732 17108 46788 17118
rect 46732 16322 46788 17052
rect 47852 17108 47908 17118
rect 47628 16996 47684 17006
rect 47628 16902 47684 16940
rect 47068 16884 47124 16894
rect 47068 16790 47124 16828
rect 47852 16882 47908 17052
rect 47852 16830 47854 16882
rect 47906 16830 47908 16882
rect 47852 16818 47908 16830
rect 46732 16270 46734 16322
rect 46786 16270 46788 16322
rect 46396 16258 46452 16268
rect 46732 16258 46788 16270
rect 46172 15986 46340 15988
rect 46172 15934 46174 15986
rect 46226 15934 46340 15986
rect 46172 15932 46340 15934
rect 46172 15922 46228 15932
rect 45052 15374 45054 15426
rect 45106 15374 45108 15426
rect 45052 15362 45108 15374
rect 45500 15428 45556 15438
rect 45500 15426 46228 15428
rect 45500 15374 45502 15426
rect 45554 15374 46228 15426
rect 45500 15372 46228 15374
rect 45500 15362 45556 15372
rect 44716 15262 44718 15314
rect 44770 15262 44772 15314
rect 44716 15250 44772 15262
rect 45948 14754 46004 15372
rect 46172 15314 46228 15372
rect 46172 15262 46174 15314
rect 46226 15262 46228 15314
rect 46172 15250 46228 15262
rect 45948 14702 45950 14754
rect 46002 14702 46004 14754
rect 44716 14644 44772 14654
rect 44716 14550 44772 14588
rect 45948 14644 46004 14702
rect 45948 14578 46004 14588
rect 41804 14530 41860 14542
rect 41804 14478 41806 14530
rect 41858 14478 41860 14530
rect 41804 14308 41860 14478
rect 42588 14420 42644 14430
rect 42588 14418 43540 14420
rect 42588 14366 42590 14418
rect 42642 14366 43540 14418
rect 42588 14364 43540 14366
rect 42588 14354 42644 14364
rect 41244 14306 41860 14308
rect 41244 14254 41246 14306
rect 41298 14254 41860 14306
rect 41244 14252 41860 14254
rect 41244 12292 41300 14252
rect 43484 13970 43540 14364
rect 46284 14418 46340 15932
rect 47292 15202 47348 15214
rect 47292 15150 47294 15202
rect 47346 15150 47348 15202
rect 47292 14756 47348 15150
rect 47292 14690 47348 14700
rect 46284 14366 46286 14418
rect 46338 14366 46340 14418
rect 46284 14354 46340 14366
rect 46508 14418 46564 14430
rect 46508 14366 46510 14418
rect 46562 14366 46564 14418
rect 43484 13918 43486 13970
rect 43538 13918 43540 13970
rect 43484 13906 43540 13918
rect 45612 14306 45668 14318
rect 45612 14254 45614 14306
rect 45666 14254 45668 14306
rect 43820 13860 43876 13870
rect 43820 13766 43876 13804
rect 45612 13860 45668 14254
rect 45612 13794 45668 13804
rect 46172 13748 46228 13758
rect 46508 13748 46564 14366
rect 45948 13746 46788 13748
rect 45948 13694 46174 13746
rect 46226 13694 46788 13746
rect 45948 13692 46788 13694
rect 45276 13634 45332 13646
rect 45276 13582 45278 13634
rect 45330 13582 45332 13634
rect 45276 13300 45332 13582
rect 45276 13234 45332 13244
rect 45724 12962 45780 12974
rect 45724 12910 45726 12962
rect 45778 12910 45780 12962
rect 43820 12404 43876 12414
rect 41244 12226 41300 12236
rect 42364 12292 42420 12302
rect 42364 10836 42420 12236
rect 43260 12292 43316 12302
rect 43260 12198 43316 12236
rect 43820 12178 43876 12348
rect 43820 12126 43822 12178
rect 43874 12126 43876 12178
rect 43820 12114 43876 12126
rect 44604 12068 44660 12078
rect 44380 12066 44660 12068
rect 44380 12014 44606 12066
rect 44658 12014 44660 12066
rect 44380 12012 44660 12014
rect 43820 11282 43876 11294
rect 43820 11230 43822 11282
rect 43874 11230 43876 11282
rect 43484 11172 43540 11182
rect 43484 11170 43764 11172
rect 43484 11118 43486 11170
rect 43538 11118 43764 11170
rect 43484 11116 43764 11118
rect 43484 11106 43540 11116
rect 42364 10834 42980 10836
rect 42364 10782 42366 10834
rect 42418 10782 42980 10834
rect 42364 10780 42980 10782
rect 40236 9874 40292 9884
rect 41132 9938 41188 9950
rect 41132 9886 41134 9938
rect 41186 9886 41188 9938
rect 39676 9136 39732 9212
rect 39452 8318 39454 8370
rect 39506 8318 39508 8370
rect 39452 8306 39508 8318
rect 39788 8258 39844 8270
rect 39788 8206 39790 8258
rect 39842 8206 39844 8258
rect 39788 8036 39844 8206
rect 39788 7970 39844 7980
rect 40012 8146 40068 8158
rect 40012 8094 40014 8146
rect 40066 8094 40068 8146
rect 38892 7364 38948 7374
rect 38892 6914 38948 7308
rect 38892 6862 38894 6914
rect 38946 6862 38948 6914
rect 38892 6850 38948 6862
rect 38668 6626 38724 6636
rect 39564 6692 39620 6702
rect 39564 6598 39620 6636
rect 40012 6692 40068 8094
rect 40460 8146 40516 8158
rect 40460 8094 40462 8146
rect 40514 8094 40516 8146
rect 40124 7364 40180 7374
rect 40124 7270 40180 7308
rect 40460 7364 40516 8094
rect 41132 8036 41188 9886
rect 41132 7942 41188 7980
rect 40572 7476 40628 7486
rect 40572 7382 40628 7420
rect 42364 7476 42420 10780
rect 42924 10610 42980 10780
rect 43708 10722 43764 11116
rect 43820 10836 43876 11230
rect 44380 11282 44436 12012
rect 44604 12002 44660 12012
rect 44380 11230 44382 11282
rect 44434 11230 44436 11282
rect 44380 11218 44436 11230
rect 44716 11284 44772 11294
rect 44716 11190 44772 11228
rect 45612 11284 45668 11294
rect 45612 11190 45668 11228
rect 43820 10770 43876 10780
rect 45724 11060 45780 12910
rect 45948 11618 46004 13692
rect 46172 13682 46228 13692
rect 46620 12850 46676 12862
rect 46620 12798 46622 12850
rect 46674 12798 46676 12850
rect 46620 11844 46676 12798
rect 46732 12066 46788 13692
rect 46732 12014 46734 12066
rect 46786 12014 46788 12066
rect 46732 12002 46788 12014
rect 46620 11778 46676 11788
rect 45948 11566 45950 11618
rect 46002 11566 46004 11618
rect 45948 11554 46004 11566
rect 46732 11396 46788 11406
rect 46732 11394 47124 11396
rect 46732 11342 46734 11394
rect 46786 11342 47124 11394
rect 46732 11340 47124 11342
rect 46732 11330 46788 11340
rect 46508 11282 46564 11294
rect 46508 11230 46510 11282
rect 46562 11230 46564 11282
rect 46508 11060 46564 11230
rect 45724 11004 46900 11060
rect 43708 10670 43710 10722
rect 43762 10670 43764 10722
rect 43708 10658 43764 10670
rect 42924 10558 42926 10610
rect 42978 10558 42980 10610
rect 42924 10546 42980 10558
rect 45724 10500 45780 11004
rect 46508 10836 46564 10846
rect 46508 10742 46564 10780
rect 46284 10724 46340 10734
rect 45836 10500 45892 10510
rect 45724 10498 45892 10500
rect 45724 10446 45838 10498
rect 45890 10446 45892 10498
rect 45724 10444 45892 10446
rect 45836 10434 45892 10444
rect 46060 10388 46116 10398
rect 43596 9940 43652 9950
rect 43596 9268 43652 9884
rect 44716 9940 44772 9950
rect 44716 9846 44772 9884
rect 46060 9938 46116 10332
rect 46060 9886 46062 9938
rect 46114 9886 46116 9938
rect 46060 9874 46116 9886
rect 46284 9940 46340 10668
rect 46844 10610 46900 11004
rect 46844 10558 46846 10610
rect 46898 10558 46900 10610
rect 47068 10724 47124 11340
rect 47068 10592 47124 10668
rect 47404 10722 47460 10734
rect 47404 10670 47406 10722
rect 47458 10670 47460 10722
rect 46844 10546 46900 10558
rect 43596 9202 43652 9212
rect 44156 9602 44212 9614
rect 44156 9550 44158 9602
rect 44210 9550 44212 9602
rect 44156 9268 44212 9550
rect 44156 9202 44212 9212
rect 45164 9156 45220 9166
rect 43596 8258 43652 8270
rect 43596 8206 43598 8258
rect 43650 8206 43652 8258
rect 42924 8036 42980 8046
rect 42924 7942 42980 7980
rect 43596 8036 43652 8206
rect 42364 7410 42420 7420
rect 40460 7298 40516 7308
rect 43484 7364 43540 7374
rect 40012 6626 40068 6636
rect 43484 6690 43540 7308
rect 43596 6916 43652 7980
rect 44604 8146 44660 8158
rect 44604 8094 44606 8146
rect 44658 8094 44660 8146
rect 43820 7476 43876 7486
rect 43820 7382 43876 7420
rect 44156 7476 44212 7486
rect 43596 6850 43652 6860
rect 43484 6638 43486 6690
rect 43538 6638 43540 6690
rect 43484 6626 43540 6638
rect 38892 6580 38948 6590
rect 38892 6130 38948 6524
rect 39676 6580 39732 6590
rect 39676 6486 39732 6524
rect 40348 6580 40404 6590
rect 38892 6078 38894 6130
rect 38946 6078 38948 6130
rect 38892 5908 38948 6078
rect 38892 5842 38948 5852
rect 40348 6466 40404 6524
rect 40348 6414 40350 6466
rect 40402 6414 40404 6466
rect 38332 5104 38388 5180
rect 38444 5794 38500 5806
rect 38444 5742 38446 5794
rect 38498 5742 38500 5794
rect 38444 5012 38500 5742
rect 38332 4228 38388 4238
rect 38220 4226 38388 4228
rect 38220 4174 38334 4226
rect 38386 4174 38388 4226
rect 38220 4172 38388 4174
rect 26236 4162 26292 4172
rect 38332 4162 38388 4172
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 3276 3666 3444 3668
rect 3276 3614 3278 3666
rect 3330 3614 3444 3666
rect 3276 3612 3444 3614
rect 3276 3602 3332 3612
rect 38444 3556 38500 4956
rect 38780 5236 38836 5246
rect 38780 4562 38836 5180
rect 40348 5124 40404 6414
rect 40348 5058 40404 5068
rect 44156 6130 44212 7420
rect 44380 7476 44436 7486
rect 44380 7382 44436 7420
rect 44604 7476 44660 8094
rect 45164 7586 45220 9100
rect 46060 9042 46116 9054
rect 46060 8990 46062 9042
rect 46114 8990 46116 9042
rect 45276 8932 45332 8942
rect 45276 8838 45332 8876
rect 45164 7534 45166 7586
rect 45218 7534 45220 7586
rect 45164 7522 45220 7534
rect 46060 8146 46116 8990
rect 46060 8094 46062 8146
rect 46114 8094 46116 8146
rect 44604 7410 44660 7420
rect 44828 6916 44884 6926
rect 44716 6804 44772 6814
rect 44156 6078 44158 6130
rect 44210 6078 44212 6130
rect 44156 5012 44212 6078
rect 44604 6578 44660 6590
rect 44604 6526 44606 6578
rect 44658 6526 44660 6578
rect 44604 6132 44660 6526
rect 44604 6066 44660 6076
rect 44716 5794 44772 6748
rect 44716 5742 44718 5794
rect 44770 5742 44772 5794
rect 44716 5730 44772 5742
rect 44828 5234 44884 6860
rect 45948 6916 46004 6926
rect 45948 6578 46004 6860
rect 46060 6804 46116 8094
rect 46060 6738 46116 6748
rect 46284 8258 46340 9884
rect 46620 9826 46676 9838
rect 46620 9774 46622 9826
rect 46674 9774 46676 9826
rect 46620 8428 46676 9774
rect 46732 9156 46788 9166
rect 46732 9062 46788 9100
rect 47068 9042 47124 9054
rect 47068 8990 47070 9042
rect 47122 8990 47124 9042
rect 47068 8482 47124 8990
rect 47068 8430 47070 8482
rect 47122 8430 47124 8482
rect 46620 8372 46788 8428
rect 47068 8418 47124 8430
rect 46284 8206 46286 8258
rect 46338 8206 46340 8258
rect 46284 6690 46340 8206
rect 46732 8260 46788 8372
rect 46732 8166 46788 8204
rect 47404 8260 47460 10670
rect 47292 7364 47348 7374
rect 47404 7364 47460 8204
rect 47292 7362 47460 7364
rect 47292 7310 47294 7362
rect 47346 7310 47460 7362
rect 47292 7308 47460 7310
rect 47292 7298 47348 7308
rect 46732 6804 46788 6814
rect 46732 6710 46788 6748
rect 46284 6638 46286 6690
rect 46338 6638 46340 6690
rect 46284 6626 46340 6638
rect 47068 6692 47124 6702
rect 47964 6692 48020 6702
rect 47068 6690 48020 6692
rect 47068 6638 47070 6690
rect 47122 6638 47966 6690
rect 48018 6638 48020 6690
rect 47068 6636 48020 6638
rect 47068 6626 47124 6636
rect 47964 6626 48020 6636
rect 45948 6526 45950 6578
rect 46002 6526 46004 6578
rect 45948 6514 46004 6526
rect 47740 6466 47796 6478
rect 47740 6414 47742 6466
rect 47794 6414 47796 6466
rect 46844 6020 46900 6030
rect 46844 5926 46900 5964
rect 47740 6020 47796 6414
rect 47740 5954 47796 5964
rect 44828 5182 44830 5234
rect 44882 5182 44884 5234
rect 44828 5170 44884 5182
rect 47516 5906 47572 5918
rect 47516 5854 47518 5906
rect 47570 5854 47572 5906
rect 44268 5124 44324 5134
rect 44268 5030 44324 5068
rect 45500 5124 45556 5134
rect 45500 5030 45556 5068
rect 46620 5122 46676 5134
rect 46620 5070 46622 5122
rect 46674 5070 46676 5122
rect 44156 4946 44212 4956
rect 46620 4676 46676 5070
rect 47516 5122 47572 5854
rect 47516 5070 47518 5122
rect 47570 5070 47572 5122
rect 46620 4610 46676 4620
rect 46956 5012 47012 5022
rect 38780 4510 38782 4562
rect 38834 4510 38836 4562
rect 38780 4498 38836 4510
rect 44604 4564 44660 4574
rect 44604 4470 44660 4508
rect 46956 4562 47012 4956
rect 47516 5012 47572 5070
rect 47516 4946 47572 4956
rect 46956 4510 46958 4562
rect 47010 4510 47012 4562
rect 46956 4498 47012 4510
rect 47292 4898 47348 4910
rect 47292 4846 47294 4898
rect 47346 4846 47348 4898
rect 47292 4564 47348 4846
rect 47292 4498 47348 4508
rect 44940 4452 44996 4462
rect 44940 4450 45108 4452
rect 44940 4398 44942 4450
rect 44994 4398 45108 4450
rect 44940 4396 45108 4398
rect 44940 4386 44996 4396
rect 38444 3490 38500 3500
rect 44268 3556 44324 3566
rect 44268 3462 44324 3500
rect 44940 3556 44996 3566
rect 44940 3462 44996 3500
rect 8652 3332 8708 3342
rect 14140 3332 14196 3342
rect 19628 3332 19684 3342
rect 25340 3332 25396 3342
rect 8428 3330 8708 3332
rect 8428 3278 8654 3330
rect 8706 3278 8708 3330
rect 8428 3276 8708 3278
rect 8428 800 8484 3276
rect 8652 3266 8708 3276
rect 13916 3330 14196 3332
rect 13916 3278 14142 3330
rect 14194 3278 14196 3330
rect 13916 3276 14196 3278
rect 13916 800 13972 3276
rect 14140 3266 14196 3276
rect 19404 3330 19684 3332
rect 19404 3278 19630 3330
rect 19682 3278 19684 3330
rect 19404 3276 19684 3278
rect 19404 800 19460 3276
rect 19628 3266 19684 3276
rect 24892 3330 25396 3332
rect 24892 3278 25342 3330
rect 25394 3278 25396 3330
rect 24892 3276 25396 3278
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 24892 800 24948 3276
rect 25340 3266 25396 3276
rect 45052 1652 45108 4396
rect 46060 3442 46116 3454
rect 46060 3390 46062 3442
rect 46114 3390 46116 3442
rect 46060 3108 46116 3390
rect 46060 3042 46116 3052
rect 45052 1586 45108 1596
rect 2912 0 3024 800
rect 8400 0 8512 800
rect 13888 0 14000 800
rect 19376 0 19488 800
rect 24864 0 24976 800
rect 30352 0 30464 800
rect 35840 0 35952 800
rect 41328 0 41440 800
rect 46816 0 46928 800
<< via2 >>
rect 47852 48188 47908 48244
rect 45948 46732 46004 46788
rect 1820 46508 1876 46564
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 39900 41132 39956 41188
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 1932 40348 1988 40404
rect 1820 34188 1876 34244
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35644 36764 35700 36820
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 32732 35586 32788 35588
rect 32732 35534 32734 35586
rect 32734 35534 32786 35586
rect 32786 35534 32788 35586
rect 32732 35532 32788 35534
rect 33964 35532 34020 35588
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 29708 34914 29764 34916
rect 29708 34862 29710 34914
rect 29710 34862 29762 34914
rect 29762 34862 29764 34914
rect 29708 34860 29764 34862
rect 31276 34860 31332 34916
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 30828 34242 30884 34244
rect 30828 34190 30830 34242
rect 30830 34190 30882 34242
rect 30882 34190 30884 34242
rect 30828 34188 30884 34190
rect 4060 33964 4116 34020
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 32508 34300 32564 34356
rect 32508 33964 32564 34020
rect 32620 34972 32676 35028
rect 31276 33346 31332 33348
rect 31276 33294 31278 33346
rect 31278 33294 31330 33346
rect 31330 33294 31332 33346
rect 31276 33292 31332 33294
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 33740 34972 33796 35028
rect 32844 34354 32900 34356
rect 32844 34302 32846 34354
rect 32846 34302 32898 34354
rect 32898 34302 32900 34354
rect 32844 34300 32900 34302
rect 33516 34300 33572 34356
rect 33180 34188 33236 34244
rect 34076 35474 34132 35476
rect 34076 35422 34078 35474
rect 34078 35422 34130 35474
rect 34130 35422 34132 35474
rect 34076 35420 34132 35422
rect 34860 35532 34916 35588
rect 36876 36652 36932 36708
rect 35644 35532 35700 35588
rect 35196 35420 35252 35476
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35868 35308 35924 35364
rect 34300 34914 34356 34916
rect 34300 34862 34302 34914
rect 34302 34862 34354 34914
rect 34354 34862 34356 34914
rect 34300 34860 34356 34862
rect 35980 34972 36036 35028
rect 36540 34860 36596 34916
rect 34076 34130 34132 34132
rect 34076 34078 34078 34130
rect 34078 34078 34130 34130
rect 34130 34078 34132 34130
rect 34076 34076 34132 34078
rect 34748 34242 34804 34244
rect 34748 34190 34750 34242
rect 34750 34190 34802 34242
rect 34802 34190 34804 34242
rect 34748 34188 34804 34190
rect 35644 34188 35700 34244
rect 34636 34076 34692 34132
rect 36652 34748 36708 34804
rect 36764 34972 36820 35028
rect 36540 34076 36596 34132
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 34636 33292 34692 33348
rect 35644 33628 35700 33684
rect 34860 32562 34916 32564
rect 34860 32510 34862 32562
rect 34862 32510 34914 32562
rect 34914 32510 34916 32562
rect 34860 32508 34916 32510
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 1820 28082 1876 28084
rect 1820 28030 1822 28082
rect 1822 28030 1874 28082
rect 1874 28030 1876 28082
rect 1820 28028 1876 28030
rect 35532 32562 35588 32564
rect 35532 32510 35534 32562
rect 35534 32510 35586 32562
rect 35586 32510 35588 32562
rect 35532 32508 35588 32510
rect 38332 36706 38388 36708
rect 38332 36654 38334 36706
rect 38334 36654 38386 36706
rect 38386 36654 38388 36706
rect 38332 36652 38388 36654
rect 37884 36204 37940 36260
rect 37996 35308 38052 35364
rect 42028 37436 42084 37492
rect 42476 37436 42532 37492
rect 38668 36370 38724 36372
rect 38668 36318 38670 36370
rect 38670 36318 38722 36370
rect 38722 36318 38724 36370
rect 38668 36316 38724 36318
rect 40348 36316 40404 36372
rect 39900 36258 39956 36260
rect 39900 36206 39902 36258
rect 39902 36206 39954 36258
rect 39954 36206 39956 36258
rect 39900 36204 39956 36206
rect 37548 34802 37604 34804
rect 37548 34750 37550 34802
rect 37550 34750 37602 34802
rect 37602 34750 37604 34802
rect 37548 34748 37604 34750
rect 38780 34690 38836 34692
rect 38780 34638 38782 34690
rect 38782 34638 38834 34690
rect 38834 34638 38836 34690
rect 38780 34636 38836 34638
rect 38556 34130 38612 34132
rect 38556 34078 38558 34130
rect 38558 34078 38610 34130
rect 38610 34078 38612 34130
rect 38556 34076 38612 34078
rect 37884 34018 37940 34020
rect 37884 33966 37886 34018
rect 37886 33966 37938 34018
rect 37938 33966 37940 34018
rect 37884 33964 37940 33966
rect 36764 33628 36820 33684
rect 36652 33404 36708 33460
rect 35868 32508 35924 32564
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 37660 33516 37716 33572
rect 39228 34636 39284 34692
rect 39452 34636 39508 34692
rect 39228 34412 39284 34468
rect 38780 33628 38836 33684
rect 39116 34076 39172 34132
rect 37884 33404 37940 33460
rect 38332 32450 38388 32452
rect 38332 32398 38334 32450
rect 38334 32398 38386 32450
rect 38386 32398 38388 32450
rect 38332 32396 38388 32398
rect 39676 34018 39732 34020
rect 39676 33966 39678 34018
rect 39678 33966 39730 34018
rect 39730 33966 39732 34018
rect 39676 33964 39732 33966
rect 39228 32396 39284 32452
rect 42140 36876 42196 36932
rect 42364 36428 42420 36484
rect 41020 36370 41076 36372
rect 41020 36318 41022 36370
rect 41022 36318 41074 36370
rect 41074 36318 41076 36370
rect 41020 36316 41076 36318
rect 43372 37490 43428 37492
rect 43372 37438 43374 37490
rect 43374 37438 43426 37490
rect 43426 37438 43428 37490
rect 43372 37436 43428 37438
rect 42812 36876 42868 36932
rect 42476 36316 42532 36372
rect 42924 36428 42980 36484
rect 43484 36482 43540 36484
rect 43484 36430 43486 36482
rect 43486 36430 43538 36482
rect 43538 36430 43540 36482
rect 43484 36428 43540 36430
rect 43708 35868 43764 35924
rect 40796 34636 40852 34692
rect 41692 34636 41748 34692
rect 44156 35868 44212 35924
rect 44268 36876 44324 36932
rect 46060 45276 46116 45332
rect 44716 44322 44772 44324
rect 44716 44270 44718 44322
rect 44718 44270 44770 44322
rect 44770 44270 44772 44322
rect 44716 44268 44772 44270
rect 45500 44322 45556 44324
rect 45500 44270 45502 44322
rect 45502 44270 45554 44322
rect 45554 44270 45556 44322
rect 45500 44268 45556 44270
rect 44716 42700 44772 42756
rect 44380 36764 44436 36820
rect 44716 41186 44772 41188
rect 44716 41134 44718 41186
rect 44718 41134 44770 41186
rect 44770 41134 44772 41186
rect 44716 41132 44772 41134
rect 44716 38556 44772 38612
rect 44716 37436 44772 37492
rect 44940 36876 44996 36932
rect 44604 36652 44660 36708
rect 43708 34412 43764 34468
rect 43820 34690 43876 34692
rect 43820 34638 43822 34690
rect 43822 34638 43874 34690
rect 43874 34638 43876 34690
rect 43820 34636 43876 34638
rect 41916 34188 41972 34244
rect 42364 34242 42420 34244
rect 42364 34190 42366 34242
rect 42366 34190 42418 34242
rect 42418 34190 42420 34242
rect 42364 34188 42420 34190
rect 43820 34076 43876 34132
rect 40460 33964 40516 34020
rect 40460 33458 40516 33460
rect 40460 33406 40462 33458
rect 40462 33406 40514 33458
rect 40514 33406 40516 33458
rect 40460 33404 40516 33406
rect 44044 33628 44100 33684
rect 44044 33180 44100 33236
rect 39900 31554 39956 31556
rect 39900 31502 39902 31554
rect 39902 31502 39954 31554
rect 39954 31502 39956 31554
rect 39900 31500 39956 31502
rect 44716 35084 44772 35140
rect 44716 34188 44772 34244
rect 45052 34130 45108 34132
rect 45052 34078 45054 34130
rect 45054 34078 45106 34130
rect 45106 34078 45108 34130
rect 45052 34076 45108 34078
rect 44380 33516 44436 33572
rect 45500 42754 45556 42756
rect 45500 42702 45502 42754
rect 45502 42702 45554 42754
rect 45554 42702 45556 42754
rect 45500 42700 45556 42702
rect 45500 41186 45556 41188
rect 45500 41134 45502 41186
rect 45502 41134 45554 41186
rect 45554 41134 45556 41186
rect 45500 41132 45556 41134
rect 45500 38556 45556 38612
rect 46060 37996 46116 38052
rect 45724 36876 45780 36932
rect 45724 36428 45780 36484
rect 45276 35196 45332 35252
rect 46172 35532 46228 35588
rect 45948 35138 46004 35140
rect 45948 35086 45950 35138
rect 45950 35086 46002 35138
rect 46002 35086 46004 35138
rect 45948 35084 46004 35086
rect 46620 43820 46676 43876
rect 46620 42364 46676 42420
rect 46620 40908 46676 40964
rect 46620 39506 46676 39508
rect 46620 39454 46622 39506
rect 46622 39454 46674 39506
rect 46674 39454 46676 39506
rect 46620 39452 46676 39454
rect 46620 36540 46676 36596
rect 47180 36876 47236 36932
rect 46396 34300 46452 34356
rect 46508 36370 46564 36372
rect 46508 36318 46510 36370
rect 46510 36318 46562 36370
rect 46562 36318 46564 36370
rect 46508 36316 46564 36318
rect 47628 36370 47684 36372
rect 47628 36318 47630 36370
rect 47630 36318 47682 36370
rect 47682 36318 47684 36370
rect 47628 36316 47684 36318
rect 46732 35756 46788 35812
rect 47068 35644 47124 35700
rect 47516 35756 47572 35812
rect 47180 35586 47236 35588
rect 47180 35534 47182 35586
rect 47182 35534 47234 35586
rect 47234 35534 47236 35586
rect 47180 35532 47236 35534
rect 45836 34242 45892 34244
rect 45836 34190 45838 34242
rect 45838 34190 45890 34242
rect 45890 34190 45892 34242
rect 45836 34188 45892 34190
rect 45164 33404 45220 33460
rect 45388 34076 45444 34132
rect 44716 33346 44772 33348
rect 44716 33294 44718 33346
rect 44718 33294 44770 33346
rect 44770 33294 44772 33346
rect 44716 33292 44772 33294
rect 45948 33570 46004 33572
rect 45948 33518 45950 33570
rect 45950 33518 46002 33570
rect 46002 33518 46004 33570
rect 45948 33516 46004 33518
rect 46284 33346 46340 33348
rect 46284 33294 46286 33346
rect 46286 33294 46338 33346
rect 46338 33294 46340 33346
rect 46284 33292 46340 33294
rect 46956 33964 47012 34020
rect 46956 33292 47012 33348
rect 46844 33234 46900 33236
rect 46844 33182 46846 33234
rect 46846 33182 46898 33234
rect 46898 33182 46900 33234
rect 46844 33180 46900 33182
rect 42252 32450 42308 32452
rect 42252 32398 42254 32450
rect 42254 32398 42306 32450
rect 42306 32398 42308 32450
rect 42252 32396 42308 32398
rect 42812 32396 42868 32452
rect 40796 31500 40852 31556
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 34860 28476 34916 28532
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 3388 26908 3444 26964
rect 6412 26908 6468 26964
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 5740 22988 5796 23044
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 8988 23042 9044 23044
rect 8988 22990 8990 23042
rect 8990 22990 9042 23042
rect 9042 22990 9044 23042
rect 8988 22988 9044 22990
rect 8540 22428 8596 22484
rect 10444 22428 10500 22484
rect 1820 21868 1876 21924
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 1820 15708 1876 15764
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 33628 26962 33684 26964
rect 33628 26910 33630 26962
rect 33630 26910 33682 26962
rect 33682 26910 33684 26962
rect 33628 26908 33684 26910
rect 36876 27858 36932 27860
rect 36876 27806 36878 27858
rect 36878 27806 36930 27858
rect 36930 27806 36932 27858
rect 36876 27804 36932 27806
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 34860 26908 34916 26964
rect 37660 26908 37716 26964
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 39788 28364 39844 28420
rect 38444 26684 38500 26740
rect 38780 27020 38836 27076
rect 39452 26684 39508 26740
rect 40124 27804 40180 27860
rect 42476 31554 42532 31556
rect 42476 31502 42478 31554
rect 42478 31502 42530 31554
rect 42530 31502 42532 31554
rect 42476 31500 42532 31502
rect 42588 28588 42644 28644
rect 43260 32172 43316 32228
rect 43372 32396 43428 32452
rect 43372 31948 43428 32004
rect 43036 31554 43092 31556
rect 43036 31502 43038 31554
rect 43038 31502 43090 31554
rect 43090 31502 43092 31554
rect 43036 31500 43092 31502
rect 43932 31948 43988 32004
rect 43596 30044 43652 30100
rect 43260 29372 43316 29428
rect 43820 29426 43876 29428
rect 43820 29374 43822 29426
rect 43822 29374 43874 29426
rect 43874 29374 43876 29426
rect 43820 29372 43876 29374
rect 44380 30156 44436 30212
rect 45836 30210 45892 30212
rect 45836 30158 45838 30210
rect 45838 30158 45890 30210
rect 45890 30158 45892 30210
rect 45836 30156 45892 30158
rect 48076 35756 48132 35812
rect 47964 35698 48020 35700
rect 47964 35646 47966 35698
rect 47966 35646 48018 35698
rect 48018 35646 48020 35698
rect 47964 35644 48020 35646
rect 47740 34076 47796 34132
rect 47964 34018 48020 34020
rect 47964 33966 47966 34018
rect 47966 33966 48018 34018
rect 48018 33966 48020 34018
rect 47964 33964 48020 33966
rect 46620 30716 46676 30772
rect 44716 29484 44772 29540
rect 44044 29260 44100 29316
rect 43260 28476 43316 28532
rect 43484 28364 43540 28420
rect 40124 27132 40180 27188
rect 40236 27244 40292 27300
rect 40460 26796 40516 26852
rect 41692 27244 41748 27300
rect 41580 27132 41636 27188
rect 41132 27074 41188 27076
rect 41132 27022 41134 27074
rect 41134 27022 41186 27074
rect 41186 27022 41188 27074
rect 41132 27020 41188 27022
rect 41468 26796 41524 26852
rect 42028 27244 42084 27300
rect 46396 30098 46452 30100
rect 46396 30046 46398 30098
rect 46398 30046 46450 30098
rect 46450 30046 46452 30098
rect 46396 30044 46452 30046
rect 47516 30098 47572 30100
rect 47516 30046 47518 30098
rect 47518 30046 47570 30098
rect 47570 30046 47572 30098
rect 47516 30044 47572 30046
rect 46732 29484 46788 29540
rect 45612 28642 45668 28644
rect 45612 28590 45614 28642
rect 45614 28590 45666 28642
rect 45666 28590 45668 28642
rect 45612 28588 45668 28590
rect 44716 28028 44772 28084
rect 45612 28252 45668 28308
rect 44604 27804 44660 27860
rect 42812 27186 42868 27188
rect 42812 27134 42814 27186
rect 42814 27134 42866 27186
rect 42866 27134 42868 27186
rect 42812 27132 42868 27134
rect 42140 27020 42196 27076
rect 42252 26908 42308 26964
rect 43820 26908 43876 26964
rect 44492 26908 44548 26964
rect 45500 26908 45556 26964
rect 45052 26796 45108 26852
rect 46284 28082 46340 28084
rect 46284 28030 46286 28082
rect 46286 28030 46338 28082
rect 46338 28030 46340 28082
rect 46284 28028 46340 28030
rect 46172 27244 46228 27300
rect 46172 26402 46228 26404
rect 46172 26350 46174 26402
rect 46174 26350 46226 26402
rect 46226 26350 46228 26402
rect 46172 26348 46228 26350
rect 44492 24780 44548 24836
rect 46620 24892 46676 24948
rect 45948 24780 46004 24836
rect 43932 23772 43988 23828
rect 42252 23212 42308 23268
rect 43596 23212 43652 23268
rect 33628 22988 33684 23044
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 20188 15036 20244 15092
rect 3388 13804 3444 13860
rect 6860 13858 6916 13860
rect 6860 13806 6862 13858
rect 6862 13806 6914 13858
rect 6914 13806 6916 13858
rect 6860 13804 6916 13806
rect 10444 13804 10500 13860
rect 11788 13858 11844 13860
rect 11788 13806 11790 13858
rect 11790 13806 11842 13858
rect 11842 13806 11844 13858
rect 11788 13804 11844 13806
rect 6188 13746 6244 13748
rect 6188 13694 6190 13746
rect 6190 13694 6242 13746
rect 6242 13694 6244 13746
rect 6188 13692 6244 13694
rect 9660 13692 9716 13748
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 8988 12236 9044 12292
rect 11004 13746 11060 13748
rect 11004 13694 11006 13746
rect 11006 13694 11058 13746
rect 11058 13694 11060 13746
rect 11004 13692 11060 13694
rect 13468 13692 13524 13748
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 1820 9602 1876 9604
rect 1820 9550 1822 9602
rect 1822 9550 1874 9602
rect 1874 9550 1876 9602
rect 1820 9548 1876 9550
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 14364 13746 14420 13748
rect 14364 13694 14366 13746
rect 14366 13694 14418 13746
rect 14418 13694 14420 13746
rect 14364 13692 14420 13694
rect 16716 13692 16772 13748
rect 13916 13634 13972 13636
rect 13916 13582 13918 13634
rect 13918 13582 13970 13634
rect 13970 13582 13972 13634
rect 13916 13580 13972 13582
rect 17052 13692 17108 13748
rect 17836 14476 17892 14532
rect 19964 14364 20020 14420
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 19404 13746 19460 13748
rect 19404 13694 19406 13746
rect 19406 13694 19458 13746
rect 19458 13694 19460 13746
rect 19404 13692 19460 13694
rect 17836 13580 17892 13636
rect 18844 13634 18900 13636
rect 18844 13582 18846 13634
rect 18846 13582 18898 13634
rect 18898 13582 18900 13634
rect 18844 13580 18900 13582
rect 14140 12290 14196 12292
rect 14140 12238 14142 12290
rect 14142 12238 14194 12290
rect 14194 12238 14196 12290
rect 14140 12236 14196 12238
rect 16268 12066 16324 12068
rect 16268 12014 16270 12066
rect 16270 12014 16322 12066
rect 16322 12014 16324 12066
rect 16268 12012 16324 12014
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 3388 5180 3444 5236
rect 1932 3442 1988 3444
rect 1932 3390 1934 3442
rect 1934 3390 1986 3442
rect 1986 3390 1988 3442
rect 1932 3388 1988 3390
rect 2940 4172 2996 4228
rect 6524 5234 6580 5236
rect 6524 5182 6526 5234
rect 6526 5182 6578 5234
rect 6578 5182 6580 5234
rect 6524 5180 6580 5182
rect 5852 5122 5908 5124
rect 5852 5070 5854 5122
rect 5854 5070 5906 5122
rect 5906 5070 5908 5122
rect 5852 5068 5908 5070
rect 16604 8370 16660 8372
rect 16604 8318 16606 8370
rect 16606 8318 16658 8370
rect 16658 8318 16660 8370
rect 16604 8316 16660 8318
rect 20972 15036 21028 15092
rect 20524 14530 20580 14532
rect 20524 14478 20526 14530
rect 20526 14478 20578 14530
rect 20578 14478 20580 14530
rect 20524 14476 20580 14478
rect 21756 15036 21812 15092
rect 22092 15202 22148 15204
rect 22092 15150 22094 15202
rect 22094 15150 22146 15202
rect 22146 15150 22148 15202
rect 22092 15148 22148 15150
rect 20636 14418 20692 14420
rect 20636 14366 20638 14418
rect 20638 14366 20690 14418
rect 20690 14366 20692 14418
rect 20636 14364 20692 14366
rect 20300 13692 20356 13748
rect 20188 13580 20244 13636
rect 21644 13580 21700 13636
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 21532 12012 21588 12068
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 18844 8316 18900 8372
rect 13804 8258 13860 8260
rect 13804 8206 13806 8258
rect 13806 8206 13858 8258
rect 13858 8206 13860 8258
rect 13804 8204 13860 8206
rect 17052 8258 17108 8260
rect 17052 8206 17054 8258
rect 17054 8206 17106 8258
rect 17106 8206 17108 8258
rect 17052 8204 17108 8206
rect 9212 5068 9268 5124
rect 8652 4956 8708 5012
rect 21532 8092 21588 8148
rect 22764 13634 22820 13636
rect 22764 13582 22766 13634
rect 22766 13582 22818 13634
rect 22818 13582 22820 13634
rect 22764 13580 22820 13582
rect 24444 12178 24500 12180
rect 24444 12126 24446 12178
rect 24446 12126 24498 12178
rect 24498 12126 24500 12178
rect 24444 12124 24500 12126
rect 24892 12178 24948 12180
rect 24892 12126 24894 12178
rect 24894 12126 24946 12178
rect 24946 12126 24948 12178
rect 24892 12124 24948 12126
rect 21644 8204 21700 8260
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 22316 8258 22372 8260
rect 22316 8206 22318 8258
rect 22318 8206 22370 8258
rect 22370 8206 22372 8258
rect 22316 8204 22372 8206
rect 21756 8146 21812 8148
rect 21756 8094 21758 8146
rect 21758 8094 21810 8146
rect 21810 8094 21812 8146
rect 21756 8092 21812 8094
rect 23100 8146 23156 8148
rect 23100 8094 23102 8146
rect 23102 8094 23154 8146
rect 23154 8094 23156 8146
rect 23100 8092 23156 8094
rect 26012 8092 26068 8148
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 14476 4956 14532 5012
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 30268 19852 30324 19908
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 43372 22876 43428 22932
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 33740 19852 33796 19908
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 38780 17612 38836 17668
rect 37884 16882 37940 16884
rect 37884 16830 37886 16882
rect 37886 16830 37938 16882
rect 37938 16830 37940 16882
rect 37884 16828 37940 16830
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 38444 16882 38500 16884
rect 38444 16830 38446 16882
rect 38446 16830 38498 16882
rect 38498 16830 38500 16882
rect 38444 16828 38500 16830
rect 44044 21980 44100 22036
rect 43596 21868 43652 21924
rect 43932 21868 43988 21924
rect 42476 19964 42532 20020
rect 39788 16828 39844 16884
rect 40236 17612 40292 17668
rect 37884 15148 37940 15204
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 39340 12290 39396 12292
rect 39340 12238 39342 12290
rect 39342 12238 39394 12290
rect 39394 12238 39396 12290
rect 39340 12236 39396 12238
rect 33740 12124 33796 12180
rect 34300 12178 34356 12180
rect 34300 12126 34302 12178
rect 34302 12126 34354 12178
rect 34354 12126 34356 12178
rect 34300 12124 34356 12126
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 26348 8034 26404 8036
rect 26348 7982 26350 8034
rect 26350 7982 26402 8034
rect 26402 7982 26404 8034
rect 26348 7980 26404 7982
rect 34860 7980 34916 8036
rect 37324 7474 37380 7476
rect 37324 7422 37326 7474
rect 37326 7422 37378 7474
rect 37378 7422 37380 7474
rect 37324 7420 37380 7422
rect 39116 9266 39172 9268
rect 39116 9214 39118 9266
rect 39118 9214 39170 9266
rect 39170 9214 39172 9266
rect 39116 9212 39172 9214
rect 37660 7420 37716 7476
rect 38332 7420 38388 7476
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 34860 6524 34916 6580
rect 33964 5180 34020 5236
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35532 5180 35588 5236
rect 36652 6690 36708 6692
rect 36652 6638 36654 6690
rect 36654 6638 36706 6690
rect 36706 6638 36708 6690
rect 36652 6636 36708 6638
rect 37324 6636 37380 6692
rect 36428 6578 36484 6580
rect 36428 6526 36430 6578
rect 36430 6526 36482 6578
rect 36482 6526 36484 6578
rect 36428 6524 36484 6526
rect 35868 4956 35924 5012
rect 36764 4956 36820 5012
rect 37548 5906 37604 5908
rect 37548 5854 37550 5906
rect 37550 5854 37602 5906
rect 37602 5854 37604 5906
rect 37548 5852 37604 5854
rect 38220 5852 38276 5908
rect 37436 4956 37492 5012
rect 36204 4450 36260 4452
rect 36204 4398 36206 4450
rect 36206 4398 36258 4450
rect 36258 4398 36260 4450
rect 36204 4396 36260 4398
rect 37548 4396 37604 4452
rect 26236 4172 26292 4228
rect 39676 9884 39732 9940
rect 41804 17666 41860 17668
rect 41804 17614 41806 17666
rect 41806 17614 41858 17666
rect 41858 17614 41860 17666
rect 41804 17612 41860 17614
rect 43260 20018 43316 20020
rect 43260 19966 43262 20018
rect 43262 19966 43314 20018
rect 43314 19966 43316 20018
rect 43260 19964 43316 19966
rect 43148 18450 43204 18452
rect 43148 18398 43150 18450
rect 43150 18398 43202 18450
rect 43202 18398 43204 18450
rect 43148 18396 43204 18398
rect 44492 23826 44548 23828
rect 44492 23774 44494 23826
rect 44494 23774 44546 23826
rect 44546 23774 44548 23826
rect 44492 23772 44548 23774
rect 46284 24556 46340 24612
rect 47404 24610 47460 24612
rect 47404 24558 47406 24610
rect 47406 24558 47458 24610
rect 47458 24558 47460 24610
rect 47404 24556 47460 24558
rect 46284 23772 46340 23828
rect 44604 23212 44660 23268
rect 45948 23548 46004 23604
rect 44716 22370 44772 22372
rect 44716 22318 44718 22370
rect 44718 22318 44770 22370
rect 44770 22318 44772 22370
rect 44716 22316 44772 22318
rect 45388 22092 45444 22148
rect 46508 23548 46564 23604
rect 44492 20802 44548 20804
rect 44492 20750 44494 20802
rect 44494 20750 44546 20802
rect 44546 20750 44548 20802
rect 44492 20748 44548 20750
rect 44380 20636 44436 20692
rect 43820 20018 43876 20020
rect 43820 19966 43822 20018
rect 43822 19966 43874 20018
rect 43874 19966 43876 20018
rect 43820 19964 43876 19966
rect 45836 20802 45892 20804
rect 45836 20750 45838 20802
rect 45838 20750 45890 20802
rect 45890 20750 45892 20802
rect 45836 20748 45892 20750
rect 46732 22988 46788 23044
rect 47516 23042 47572 23044
rect 47516 22990 47518 23042
rect 47518 22990 47570 23042
rect 47570 22990 47572 23042
rect 47516 22988 47572 22990
rect 46732 22370 46788 22372
rect 46732 22318 46734 22370
rect 46734 22318 46786 22370
rect 46786 22318 46788 22370
rect 46732 22316 46788 22318
rect 45948 20636 46004 20692
rect 47740 22146 47796 22148
rect 47740 22094 47742 22146
rect 47742 22094 47794 22146
rect 47794 22094 47796 22146
rect 47740 22092 47796 22094
rect 45276 20524 45332 20580
rect 46396 20690 46452 20692
rect 46396 20638 46398 20690
rect 46398 20638 46450 20690
rect 46450 20638 46452 20690
rect 46396 20636 46452 20638
rect 43372 18396 43428 18452
rect 43708 18450 43764 18452
rect 43708 18398 43710 18450
rect 43710 18398 43762 18450
rect 43762 18398 43764 18450
rect 43708 18396 43764 18398
rect 44716 17836 44772 17892
rect 45612 17890 45668 17892
rect 45612 17838 45614 17890
rect 45614 17838 45666 17890
rect 45666 17838 45668 17890
rect 45612 17836 45668 17838
rect 46620 19122 46676 19124
rect 46620 19070 46622 19122
rect 46622 19070 46674 19122
rect 46674 19070 46676 19122
rect 46620 19068 46676 19070
rect 42924 17778 42980 17780
rect 42924 17726 42926 17778
rect 42926 17726 42978 17778
rect 42978 17726 42980 17778
rect 42924 17724 42980 17726
rect 45052 17724 45108 17780
rect 42476 17666 42532 17668
rect 42476 17614 42478 17666
rect 42478 17614 42530 17666
rect 42530 17614 42532 17666
rect 42476 17612 42532 17614
rect 44604 17666 44660 17668
rect 44604 17614 44606 17666
rect 44606 17614 44658 17666
rect 44658 17614 44660 17666
rect 44604 17612 44660 17614
rect 44156 17500 44212 17556
rect 41244 16828 41300 16884
rect 41916 15484 41972 15540
rect 42476 15538 42532 15540
rect 42476 15486 42478 15538
rect 42478 15486 42530 15538
rect 42530 15486 42532 15538
rect 42476 15484 42532 15486
rect 44492 16828 44548 16884
rect 42924 15484 42980 15540
rect 44044 15372 44100 15428
rect 44716 15932 44772 15988
rect 44716 15372 44772 15428
rect 42812 15314 42868 15316
rect 42812 15262 42814 15314
rect 42814 15262 42866 15314
rect 42866 15262 42868 15314
rect 42812 15260 42868 15262
rect 44380 15314 44436 15316
rect 44380 15262 44382 15314
rect 44382 15262 44434 15314
rect 44434 15262 44436 15314
rect 44380 15260 44436 15262
rect 46172 17724 46228 17780
rect 45612 15986 45668 15988
rect 45612 15934 45614 15986
rect 45614 15934 45666 15986
rect 45666 15934 45668 15986
rect 45612 15932 45668 15934
rect 46508 17554 46564 17556
rect 46508 17502 46510 17554
rect 46510 17502 46562 17554
rect 46562 17502 46564 17554
rect 46508 17500 46564 17502
rect 46284 16994 46340 16996
rect 46284 16942 46286 16994
rect 46286 16942 46338 16994
rect 46338 16942 46340 16994
rect 46284 16940 46340 16942
rect 46732 17052 46788 17108
rect 47852 17052 47908 17108
rect 47628 16994 47684 16996
rect 47628 16942 47630 16994
rect 47630 16942 47682 16994
rect 47682 16942 47684 16994
rect 47628 16940 47684 16942
rect 47068 16882 47124 16884
rect 47068 16830 47070 16882
rect 47070 16830 47122 16882
rect 47122 16830 47124 16882
rect 47068 16828 47124 16830
rect 44716 14642 44772 14644
rect 44716 14590 44718 14642
rect 44718 14590 44770 14642
rect 44770 14590 44772 14642
rect 44716 14588 44772 14590
rect 45948 14588 46004 14644
rect 47292 14700 47348 14756
rect 43820 13858 43876 13860
rect 43820 13806 43822 13858
rect 43822 13806 43874 13858
rect 43874 13806 43876 13858
rect 43820 13804 43876 13806
rect 45612 13804 45668 13860
rect 45276 13244 45332 13300
rect 43820 12348 43876 12404
rect 41244 12236 41300 12292
rect 42364 12236 42420 12292
rect 43260 12290 43316 12292
rect 43260 12238 43262 12290
rect 43262 12238 43314 12290
rect 43314 12238 43316 12290
rect 43260 12236 43316 12238
rect 40236 9884 40292 9940
rect 39676 9266 39732 9268
rect 39676 9214 39678 9266
rect 39678 9214 39730 9266
rect 39730 9214 39732 9266
rect 39676 9212 39732 9214
rect 39788 7980 39844 8036
rect 38892 7308 38948 7364
rect 38668 6636 38724 6692
rect 39564 6690 39620 6692
rect 39564 6638 39566 6690
rect 39566 6638 39618 6690
rect 39618 6638 39620 6690
rect 39564 6636 39620 6638
rect 40124 7362 40180 7364
rect 40124 7310 40126 7362
rect 40126 7310 40178 7362
rect 40178 7310 40180 7362
rect 40124 7308 40180 7310
rect 41132 8034 41188 8036
rect 41132 7982 41134 8034
rect 41134 7982 41186 8034
rect 41186 7982 41188 8034
rect 41132 7980 41188 7982
rect 40572 7474 40628 7476
rect 40572 7422 40574 7474
rect 40574 7422 40626 7474
rect 40626 7422 40628 7474
rect 40572 7420 40628 7422
rect 44716 11282 44772 11284
rect 44716 11230 44718 11282
rect 44718 11230 44770 11282
rect 44770 11230 44772 11282
rect 44716 11228 44772 11230
rect 45612 11282 45668 11284
rect 45612 11230 45614 11282
rect 45614 11230 45666 11282
rect 45666 11230 45668 11282
rect 45612 11228 45668 11230
rect 43820 10780 43876 10836
rect 46620 11788 46676 11844
rect 46508 10834 46564 10836
rect 46508 10782 46510 10834
rect 46510 10782 46562 10834
rect 46562 10782 46564 10834
rect 46508 10780 46564 10782
rect 46284 10668 46340 10724
rect 46060 10332 46116 10388
rect 43596 9938 43652 9940
rect 43596 9886 43598 9938
rect 43598 9886 43650 9938
rect 43650 9886 43652 9938
rect 43596 9884 43652 9886
rect 44716 9938 44772 9940
rect 44716 9886 44718 9938
rect 44718 9886 44770 9938
rect 44770 9886 44772 9938
rect 44716 9884 44772 9886
rect 47068 10722 47124 10724
rect 47068 10670 47070 10722
rect 47070 10670 47122 10722
rect 47122 10670 47124 10722
rect 47068 10668 47124 10670
rect 46284 9884 46340 9940
rect 43596 9212 43652 9268
rect 44156 9212 44212 9268
rect 45164 9100 45220 9156
rect 42924 8034 42980 8036
rect 42924 7982 42926 8034
rect 42926 7982 42978 8034
rect 42978 7982 42980 8034
rect 42924 7980 42980 7982
rect 43596 7980 43652 8036
rect 42364 7420 42420 7476
rect 40460 7308 40516 7364
rect 43484 7308 43540 7364
rect 40012 6636 40068 6692
rect 43820 7474 43876 7476
rect 43820 7422 43822 7474
rect 43822 7422 43874 7474
rect 43874 7422 43876 7474
rect 43820 7420 43876 7422
rect 44156 7420 44212 7476
rect 43596 6860 43652 6916
rect 38892 6524 38948 6580
rect 39676 6578 39732 6580
rect 39676 6526 39678 6578
rect 39678 6526 39730 6578
rect 39730 6526 39732 6578
rect 39676 6524 39732 6526
rect 40348 6524 40404 6580
rect 38892 5852 38948 5908
rect 38332 5234 38388 5236
rect 38332 5182 38334 5234
rect 38334 5182 38386 5234
rect 38386 5182 38388 5234
rect 38332 5180 38388 5182
rect 38444 4956 38500 5012
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 38780 5180 38836 5236
rect 40348 5068 40404 5124
rect 44380 7474 44436 7476
rect 44380 7422 44382 7474
rect 44382 7422 44434 7474
rect 44434 7422 44436 7474
rect 44380 7420 44436 7422
rect 45276 8930 45332 8932
rect 45276 8878 45278 8930
rect 45278 8878 45330 8930
rect 45330 8878 45332 8930
rect 45276 8876 45332 8878
rect 44604 7420 44660 7476
rect 44828 6860 44884 6916
rect 44716 6748 44772 6804
rect 44604 6076 44660 6132
rect 45948 6860 46004 6916
rect 46060 6748 46116 6804
rect 46732 9154 46788 9156
rect 46732 9102 46734 9154
rect 46734 9102 46786 9154
rect 46786 9102 46788 9154
rect 46732 9100 46788 9102
rect 46732 8258 46788 8260
rect 46732 8206 46734 8258
rect 46734 8206 46786 8258
rect 46786 8206 46788 8258
rect 46732 8204 46788 8206
rect 47404 8204 47460 8260
rect 46732 6802 46788 6804
rect 46732 6750 46734 6802
rect 46734 6750 46786 6802
rect 46786 6750 46788 6802
rect 46732 6748 46788 6750
rect 46844 6018 46900 6020
rect 46844 5966 46846 6018
rect 46846 5966 46898 6018
rect 46898 5966 46900 6018
rect 46844 5964 46900 5966
rect 47740 5964 47796 6020
rect 44268 5122 44324 5124
rect 44268 5070 44270 5122
rect 44270 5070 44322 5122
rect 44322 5070 44324 5122
rect 44268 5068 44324 5070
rect 45500 5122 45556 5124
rect 45500 5070 45502 5122
rect 45502 5070 45554 5122
rect 45554 5070 45556 5122
rect 45500 5068 45556 5070
rect 44156 4956 44212 5012
rect 46620 4620 46676 4676
rect 46956 4956 47012 5012
rect 44604 4562 44660 4564
rect 44604 4510 44606 4562
rect 44606 4510 44658 4562
rect 44658 4510 44660 4562
rect 44604 4508 44660 4510
rect 47516 4956 47572 5012
rect 47292 4508 47348 4564
rect 38444 3500 38500 3556
rect 44268 3554 44324 3556
rect 44268 3502 44270 3554
rect 44270 3502 44322 3554
rect 44322 3502 44324 3554
rect 44268 3500 44324 3502
rect 44940 3554 44996 3556
rect 44940 3502 44942 3554
rect 44942 3502 44994 3554
rect 44994 3502 44996 3554
rect 44940 3500 44996 3502
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 46060 3052 46116 3108
rect 45052 1596 45108 1652
<< metal3 >>
rect 49200 48244 50000 48272
rect 47842 48188 47852 48244
rect 47908 48188 50000 48244
rect 49200 48160 50000 48188
rect 49200 46788 50000 46816
rect 45938 46732 45948 46788
rect 46004 46732 50000 46788
rect 49200 46704 50000 46732
rect 0 46564 800 46592
rect 0 46508 1820 46564
rect 1876 46508 1886 46564
rect 0 46480 800 46508
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 49200 45332 50000 45360
rect 46050 45276 46060 45332
rect 46116 45276 50000 45332
rect 49200 45248 50000 45276
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 44706 44268 44716 44324
rect 44772 44268 45500 44324
rect 45556 44268 45566 44324
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 49200 43876 50000 43904
rect 46610 43820 46620 43876
rect 46676 43820 50000 43876
rect 49200 43792 50000 43820
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 44706 42700 44716 42756
rect 44772 42700 45500 42756
rect 45556 42700 45566 42756
rect 49200 42420 50000 42448
rect 46610 42364 46620 42420
rect 46676 42364 50000 42420
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 49200 42336 50000 42364
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 39890 41132 39900 41188
rect 39956 41132 44716 41188
rect 44772 41132 45500 41188
rect 45556 41132 45566 41188
rect 49200 40964 50000 40992
rect 46610 40908 46620 40964
rect 46676 40908 50000 40964
rect 49200 40880 50000 40908
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 0 40404 800 40432
rect 0 40348 1932 40404
rect 1988 40348 1998 40404
rect 0 40320 800 40348
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 49200 39508 50000 39536
rect 46610 39452 46620 39508
rect 46676 39452 50000 39508
rect 49200 39424 50000 39452
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 44706 38556 44716 38612
rect 44772 38556 45500 38612
rect 45556 38556 45566 38612
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 49200 38052 50000 38080
rect 46050 37996 46060 38052
rect 46116 37996 50000 38052
rect 49200 37968 50000 37996
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 42018 37436 42028 37492
rect 42084 37436 42476 37492
rect 42532 37436 43372 37492
rect 43428 37436 44716 37492
rect 44772 37436 44782 37492
rect 42130 36876 42140 36932
rect 42196 36876 42812 36932
rect 42868 36876 44268 36932
rect 44324 36876 44940 36932
rect 44996 36876 45006 36932
rect 45714 36876 45724 36932
rect 45780 36876 47180 36932
rect 47236 36876 47246 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 35634 36764 35644 36820
rect 35700 36764 44380 36820
rect 44436 36764 44446 36820
rect 36866 36652 36876 36708
rect 36932 36652 38332 36708
rect 38388 36652 44604 36708
rect 44660 36652 44670 36708
rect 49200 36596 50000 36624
rect 46610 36540 46620 36596
rect 46676 36540 50000 36596
rect 49200 36512 50000 36540
rect 40348 36428 42364 36484
rect 42420 36428 42430 36484
rect 42914 36428 42924 36484
rect 42980 36428 43484 36484
rect 43540 36428 45724 36484
rect 45780 36428 45790 36484
rect 40348 36372 40404 36428
rect 38658 36316 38668 36372
rect 38724 36316 40348 36372
rect 40404 36316 40414 36372
rect 41010 36316 41020 36372
rect 41076 36316 42476 36372
rect 42532 36316 42542 36372
rect 46498 36316 46508 36372
rect 46564 36316 47628 36372
rect 47684 36316 47694 36372
rect 37874 36204 37884 36260
rect 37940 36204 39900 36260
rect 39956 36204 39966 36260
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 32722 35532 32732 35588
rect 32788 35532 33964 35588
rect 34020 35532 34030 35588
rect 34850 35532 34860 35588
rect 34916 35532 35644 35588
rect 35700 35532 35710 35588
rect 34860 35476 34916 35532
rect 34066 35420 34076 35476
rect 34132 35420 34916 35476
rect 35186 35420 35196 35476
rect 35252 35420 38276 35476
rect 35858 35308 35868 35364
rect 35924 35308 37996 35364
rect 38052 35308 38062 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 38220 35252 38276 35420
rect 43652 35252 43708 35924
rect 43764 35868 44156 35924
rect 44212 35868 44222 35924
rect 46722 35756 46732 35812
rect 46788 35756 47516 35812
rect 47572 35756 48076 35812
rect 48132 35756 48142 35812
rect 47058 35644 47068 35700
rect 47124 35644 47964 35700
rect 48020 35644 48030 35700
rect 46162 35532 46172 35588
rect 46228 35532 47180 35588
rect 47236 35532 47246 35588
rect 38220 35196 43708 35252
rect 45266 35196 45276 35252
rect 45332 35196 46228 35252
rect 46172 35140 46228 35196
rect 49200 35140 50000 35168
rect 44706 35084 44716 35140
rect 44772 35084 45948 35140
rect 46004 35084 46014 35140
rect 46172 35084 50000 35140
rect 49200 35056 50000 35084
rect 32610 34972 32620 35028
rect 32676 34972 33740 35028
rect 33796 34972 33806 35028
rect 35970 34972 35980 35028
rect 36036 34972 36764 35028
rect 36820 34972 36830 35028
rect 29698 34860 29708 34916
rect 29764 34860 31276 34916
rect 31332 34860 31342 34916
rect 34290 34860 34300 34916
rect 34356 34860 36540 34916
rect 36596 34860 36606 34916
rect 36642 34748 36652 34804
rect 36708 34748 37548 34804
rect 37604 34748 37614 34804
rect 38770 34636 38780 34692
rect 38836 34636 39228 34692
rect 39284 34636 39452 34692
rect 39508 34636 40796 34692
rect 40852 34636 41692 34692
rect 41748 34636 43820 34692
rect 43876 34636 43886 34692
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 39218 34412 39228 34468
rect 39284 34412 43708 34468
rect 43764 34412 43774 34468
rect 32498 34300 32508 34356
rect 32564 34300 32844 34356
rect 32900 34300 33516 34356
rect 33572 34300 46396 34356
rect 46452 34300 46462 34356
rect 0 34244 800 34272
rect 0 34188 1820 34244
rect 1876 34188 1886 34244
rect 30818 34188 30828 34244
rect 30884 34188 33180 34244
rect 33236 34188 33246 34244
rect 34738 34188 34748 34244
rect 34804 34188 35644 34244
rect 35700 34188 35710 34244
rect 41906 34188 41916 34244
rect 41972 34188 42364 34244
rect 42420 34188 42430 34244
rect 44706 34188 44716 34244
rect 44772 34188 45836 34244
rect 45892 34188 45902 34244
rect 0 34160 800 34188
rect 34066 34076 34076 34132
rect 34132 34076 34636 34132
rect 34692 34076 34702 34132
rect 36530 34076 36540 34132
rect 36596 34076 38556 34132
rect 38612 34076 39116 34132
rect 39172 34076 39182 34132
rect 43810 34076 43820 34132
rect 43876 34076 45052 34132
rect 45108 34076 45118 34132
rect 45378 34076 45388 34132
rect 45444 34076 47740 34132
rect 47796 34076 47806 34132
rect 4050 33964 4060 34020
rect 4116 33964 32508 34020
rect 32564 33964 32574 34020
rect 37874 33964 37884 34020
rect 37940 33964 39676 34020
rect 39732 33964 40460 34020
rect 40516 33964 40526 34020
rect 46946 33964 46956 34020
rect 47012 33964 47964 34020
rect 48020 33964 48030 34020
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 49200 33684 50000 33712
rect 35634 33628 35644 33684
rect 35700 33628 36764 33684
rect 36820 33628 38780 33684
rect 38836 33628 38846 33684
rect 44034 33628 44044 33684
rect 44100 33628 50000 33684
rect 37660 33572 37716 33628
rect 49200 33600 50000 33628
rect 37650 33516 37660 33572
rect 37716 33516 37726 33572
rect 44370 33516 44380 33572
rect 44436 33516 45948 33572
rect 46004 33516 46014 33572
rect 36642 33404 36652 33460
rect 36708 33404 37884 33460
rect 37940 33404 37950 33460
rect 40450 33404 40460 33460
rect 40516 33404 45164 33460
rect 45220 33404 45230 33460
rect 31266 33292 31276 33348
rect 31332 33292 34636 33348
rect 34692 33292 34702 33348
rect 44706 33292 44716 33348
rect 44772 33292 46284 33348
rect 46340 33292 46956 33348
rect 47012 33292 47022 33348
rect 44034 33180 44044 33236
rect 44100 33180 46844 33236
rect 46900 33180 46910 33236
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 34850 32508 34860 32564
rect 34916 32508 35532 32564
rect 35588 32508 35598 32564
rect 35858 32508 35868 32564
rect 35924 32508 35934 32564
rect 35868 32452 35924 32508
rect 35868 32396 38332 32452
rect 38388 32396 39228 32452
rect 39284 32396 39294 32452
rect 42242 32396 42252 32452
rect 42308 32396 42812 32452
rect 42868 32396 43372 32452
rect 43428 32396 43438 32452
rect 49200 32228 50000 32256
rect 43250 32172 43260 32228
rect 43316 32172 50000 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 49200 32144 50000 32172
rect 43362 31948 43372 32004
rect 43428 31948 43932 32004
rect 43988 31948 43998 32004
rect 39890 31500 39900 31556
rect 39956 31500 40796 31556
rect 40852 31500 42476 31556
rect 42532 31500 43036 31556
rect 43092 31500 43102 31556
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 49200 30772 50000 30800
rect 46610 30716 46620 30772
rect 46676 30716 50000 30772
rect 49200 30688 50000 30716
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 44370 30156 44380 30212
rect 44436 30156 45836 30212
rect 45892 30156 45902 30212
rect 43586 30044 43596 30100
rect 43652 30044 46396 30100
rect 46452 30044 47516 30100
rect 47572 30044 47582 30100
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 44706 29484 44716 29540
rect 44772 29484 46732 29540
rect 46788 29484 46798 29540
rect 43250 29372 43260 29428
rect 43316 29372 43820 29428
rect 43876 29372 43886 29428
rect 49200 29316 50000 29344
rect 44034 29260 44044 29316
rect 44100 29260 50000 29316
rect 49200 29232 50000 29260
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 42578 28588 42588 28644
rect 42644 28588 45612 28644
rect 45668 28588 45678 28644
rect 34850 28476 34860 28532
rect 34916 28476 43260 28532
rect 43316 28476 43326 28532
rect 39778 28364 39788 28420
rect 39844 28364 43484 28420
rect 43540 28364 43708 28420
rect 43652 28308 43708 28364
rect 43652 28252 45612 28308
rect 45668 28252 45678 28308
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 0 28084 800 28112
rect 0 28028 1820 28084
rect 1876 28028 1886 28084
rect 44706 28028 44716 28084
rect 44772 28028 46284 28084
rect 46340 28028 46350 28084
rect 0 28000 800 28028
rect 49200 27860 50000 27888
rect 36866 27804 36876 27860
rect 36932 27804 40124 27860
rect 40180 27804 40190 27860
rect 44594 27804 44604 27860
rect 44660 27804 50000 27860
rect 49200 27776 50000 27804
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 40226 27244 40236 27300
rect 40292 27244 41692 27300
rect 41748 27244 42028 27300
rect 42084 27244 46172 27300
rect 46228 27244 46238 27300
rect 40114 27132 40124 27188
rect 40180 27132 41580 27188
rect 41636 27132 42812 27188
rect 42868 27132 42878 27188
rect 38770 27020 38780 27076
rect 38836 27020 41132 27076
rect 41188 27020 41198 27076
rect 42130 27020 42140 27076
rect 42196 27020 43708 27076
rect 43652 26964 43708 27020
rect 3378 26908 3388 26964
rect 3444 26908 6412 26964
rect 6468 26908 6478 26964
rect 33618 26908 33628 26964
rect 33684 26908 34860 26964
rect 34916 26908 34926 26964
rect 37650 26908 37660 26964
rect 37716 26908 42252 26964
rect 42308 26908 42318 26964
rect 43652 26908 43820 26964
rect 43876 26908 44492 26964
rect 44548 26908 45500 26964
rect 45556 26908 45566 26964
rect 40450 26796 40460 26852
rect 40516 26796 41468 26852
rect 41524 26796 45052 26852
rect 45108 26796 45118 26852
rect 38434 26684 38444 26740
rect 38500 26684 39452 26740
rect 39508 26684 39518 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 49200 26404 50000 26432
rect 46162 26348 46172 26404
rect 46228 26348 50000 26404
rect 49200 26320 50000 26348
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 49200 24948 50000 24976
rect 46610 24892 46620 24948
rect 46676 24892 50000 24948
rect 49200 24864 50000 24892
rect 44482 24780 44492 24836
rect 44548 24780 45948 24836
rect 46004 24780 46014 24836
rect 46274 24556 46284 24612
rect 46340 24556 47404 24612
rect 47460 24556 47470 24612
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 43922 23772 43932 23828
rect 43988 23772 44492 23828
rect 44548 23772 46284 23828
rect 46340 23772 46350 23828
rect 45938 23548 45948 23604
rect 46004 23548 46508 23604
rect 46564 23548 46574 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 49200 23492 50000 23520
rect 47740 23436 50000 23492
rect 42242 23212 42252 23268
rect 42308 23212 43596 23268
rect 43652 23212 44604 23268
rect 44660 23212 44670 23268
rect 5730 22988 5740 23044
rect 5796 22988 8988 23044
rect 9044 22988 33628 23044
rect 33684 22988 33694 23044
rect 46722 22988 46732 23044
rect 46788 22988 47516 23044
rect 47572 22988 47582 23044
rect 47740 22932 47796 23436
rect 49200 23408 50000 23436
rect 43362 22876 43372 22932
rect 43428 22876 47796 22932
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 8530 22428 8540 22484
rect 8596 22428 10444 22484
rect 10500 22428 10510 22484
rect 44706 22316 44716 22372
rect 44772 22316 46732 22372
rect 46788 22316 46798 22372
rect 45378 22092 45388 22148
rect 45444 22092 47740 22148
rect 47796 22092 47806 22148
rect 49200 22036 50000 22064
rect 44034 21980 44044 22036
rect 44100 21980 50000 22036
rect 0 21924 800 21952
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 49200 21952 50000 21980
rect 0 21868 1820 21924
rect 1876 21868 1886 21924
rect 43586 21868 43596 21924
rect 43652 21868 43932 21924
rect 43988 21868 43998 21924
rect 0 21840 800 21868
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 44482 20748 44492 20804
rect 44548 20748 45836 20804
rect 45892 20748 45902 20804
rect 44370 20636 44380 20692
rect 44436 20636 45948 20692
rect 46004 20636 46396 20692
rect 46452 20636 46462 20692
rect 49200 20580 50000 20608
rect 45266 20524 45276 20580
rect 45332 20524 50000 20580
rect 49200 20496 50000 20524
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 42466 19964 42476 20020
rect 42532 19964 43260 20020
rect 43316 19964 43820 20020
rect 43876 19964 43886 20020
rect 30258 19852 30268 19908
rect 30324 19852 33740 19908
rect 33796 19852 33806 19908
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 49200 19124 50000 19152
rect 46610 19068 46620 19124
rect 46676 19068 50000 19124
rect 49200 19040 50000 19068
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 43138 18396 43148 18452
rect 43204 18396 43372 18452
rect 43428 18396 43708 18452
rect 43764 18396 43774 18452
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 44706 17836 44716 17892
rect 44772 17836 45612 17892
rect 45668 17836 45678 17892
rect 42914 17724 42924 17780
rect 42980 17724 45052 17780
rect 45108 17724 46172 17780
rect 46228 17724 46238 17780
rect 49200 17668 50000 17696
rect 38770 17612 38780 17668
rect 38836 17612 40236 17668
rect 40292 17612 41804 17668
rect 41860 17612 42476 17668
rect 42532 17612 42542 17668
rect 44594 17612 44604 17668
rect 44660 17612 50000 17668
rect 49200 17584 50000 17612
rect 44146 17500 44156 17556
rect 44212 17500 46508 17556
rect 46564 17500 46574 17556
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 46722 17052 46732 17108
rect 46788 17052 47852 17108
rect 47908 17052 47918 17108
rect 46274 16940 46284 16996
rect 46340 16940 47628 16996
rect 47684 16940 47694 16996
rect 37874 16828 37884 16884
rect 37940 16828 38444 16884
rect 38500 16828 39788 16884
rect 39844 16828 39854 16884
rect 41234 16828 41244 16884
rect 41300 16828 44492 16884
rect 44548 16828 47068 16884
rect 47124 16828 47134 16884
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 49200 16212 50000 16240
rect 49084 16156 50000 16212
rect 44706 15932 44716 15988
rect 44772 15932 45612 15988
rect 45668 15932 45678 15988
rect 49084 15876 49140 16156
rect 49200 16128 50000 16156
rect 49084 15820 49364 15876
rect 0 15764 800 15792
rect 0 15708 1820 15764
rect 1876 15708 1886 15764
rect 0 15680 800 15708
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 49308 15540 49364 15820
rect 41906 15484 41916 15540
rect 41972 15484 42476 15540
rect 42532 15484 42542 15540
rect 42914 15484 42924 15540
rect 42980 15484 49364 15540
rect 44034 15372 44044 15428
rect 44100 15372 44716 15428
rect 44772 15372 44782 15428
rect 42802 15260 42812 15316
rect 42868 15260 44380 15316
rect 44436 15260 44446 15316
rect 22082 15148 22092 15204
rect 22148 15148 37884 15204
rect 37940 15148 37950 15204
rect 20178 15036 20188 15092
rect 20244 15036 20972 15092
rect 21028 15036 21756 15092
rect 21812 15036 21822 15092
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 49200 14756 50000 14784
rect 47282 14700 47292 14756
rect 47348 14700 50000 14756
rect 49200 14672 50000 14700
rect 44706 14588 44716 14644
rect 44772 14588 45948 14644
rect 46004 14588 46014 14644
rect 17826 14476 17836 14532
rect 17892 14476 20524 14532
rect 20580 14476 20590 14532
rect 19954 14364 19964 14420
rect 20020 14364 20636 14420
rect 20692 14364 20702 14420
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 3378 13804 3388 13860
rect 3444 13804 6860 13860
rect 6916 13804 6926 13860
rect 10434 13804 10444 13860
rect 10500 13804 11788 13860
rect 11844 13804 11854 13860
rect 43810 13804 43820 13860
rect 43876 13804 45612 13860
rect 45668 13804 45678 13860
rect 6178 13692 6188 13748
rect 6244 13692 9660 13748
rect 9716 13692 11004 13748
rect 11060 13692 13468 13748
rect 13524 13692 14364 13748
rect 14420 13692 16716 13748
rect 16772 13692 17052 13748
rect 17108 13692 19404 13748
rect 19460 13692 20300 13748
rect 20356 13692 21700 13748
rect 21644 13636 21700 13692
rect 13906 13580 13916 13636
rect 13972 13580 17836 13636
rect 17892 13580 17902 13636
rect 18834 13580 18844 13636
rect 18900 13580 20188 13636
rect 20244 13580 20254 13636
rect 21634 13580 21644 13636
rect 21700 13580 22764 13636
rect 22820 13580 22830 13636
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 49200 13300 50000 13328
rect 45266 13244 45276 13300
rect 45332 13244 50000 13300
rect 49200 13216 50000 13244
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 43260 12348 43820 12404
rect 43876 12348 43886 12404
rect 43260 12292 43316 12348
rect 8978 12236 8988 12292
rect 9044 12236 14140 12292
rect 14196 12236 14206 12292
rect 39330 12236 39340 12292
rect 39396 12236 41244 12292
rect 41300 12236 42364 12292
rect 42420 12236 43260 12292
rect 43316 12236 43326 12292
rect 24434 12124 24444 12180
rect 24500 12124 24892 12180
rect 24948 12124 33740 12180
rect 33796 12124 34300 12180
rect 34356 12124 34366 12180
rect 16258 12012 16268 12068
rect 16324 12012 21532 12068
rect 21588 12012 21598 12068
rect 49200 11844 50000 11872
rect 46610 11788 46620 11844
rect 46676 11788 50000 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 49200 11760 50000 11788
rect 44706 11228 44716 11284
rect 44772 11228 45612 11284
rect 45668 11228 45678 11284
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 43810 10780 43820 10836
rect 43876 10780 46508 10836
rect 46564 10780 46574 10836
rect 46274 10668 46284 10724
rect 46340 10668 47068 10724
rect 47124 10668 47134 10724
rect 49200 10388 50000 10416
rect 46050 10332 46060 10388
rect 46116 10332 50000 10388
rect 49200 10304 50000 10332
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 39666 9884 39676 9940
rect 39732 9884 40236 9940
rect 40292 9884 43596 9940
rect 43652 9884 43662 9940
rect 44706 9884 44716 9940
rect 44772 9884 46284 9940
rect 46340 9884 46350 9940
rect 0 9604 800 9632
rect 0 9548 1820 9604
rect 1876 9548 1886 9604
rect 0 9520 800 9548
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 39106 9212 39116 9268
rect 39172 9212 39676 9268
rect 39732 9212 39742 9268
rect 43586 9212 43596 9268
rect 43652 9212 44156 9268
rect 44212 9212 44222 9268
rect 45154 9100 45164 9156
rect 45220 9100 46732 9156
rect 46788 9100 46798 9156
rect 49200 8932 50000 8960
rect 45266 8876 45276 8932
rect 45332 8876 50000 8932
rect 49200 8848 50000 8876
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 16594 8316 16604 8372
rect 16660 8316 18844 8372
rect 18900 8316 18910 8372
rect 13794 8204 13804 8260
rect 13860 8204 17052 8260
rect 17108 8204 21644 8260
rect 21700 8204 22316 8260
rect 22372 8204 22382 8260
rect 46722 8204 46732 8260
rect 46788 8204 47404 8260
rect 47460 8204 47470 8260
rect 21522 8092 21532 8148
rect 21588 8092 21756 8148
rect 21812 8092 23100 8148
rect 23156 8092 26012 8148
rect 26068 8092 26078 8148
rect 26338 7980 26348 8036
rect 26404 7980 34860 8036
rect 34916 7980 34926 8036
rect 39778 7980 39788 8036
rect 39844 7980 41132 8036
rect 41188 7980 42924 8036
rect 42980 7980 43596 8036
rect 43652 7980 43662 8036
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 49200 7476 50000 7504
rect 37314 7420 37324 7476
rect 37380 7420 37660 7476
rect 37716 7420 38332 7476
rect 38388 7420 40572 7476
rect 40628 7420 42364 7476
rect 42420 7420 43820 7476
rect 43876 7420 44156 7476
rect 44212 7420 44380 7476
rect 44436 7420 44446 7476
rect 44594 7420 44604 7476
rect 44660 7420 50000 7476
rect 49200 7392 50000 7420
rect 38882 7308 38892 7364
rect 38948 7308 40124 7364
rect 40180 7308 40460 7364
rect 40516 7308 43484 7364
rect 43540 7308 43550 7364
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 43586 6860 43596 6916
rect 43652 6860 44828 6916
rect 44884 6860 45948 6916
rect 46004 6860 46014 6916
rect 44706 6748 44716 6804
rect 44772 6748 46060 6804
rect 46116 6748 46732 6804
rect 46788 6748 46798 6804
rect 36642 6636 36652 6692
rect 36708 6636 37324 6692
rect 37380 6636 38668 6692
rect 38724 6636 39564 6692
rect 39620 6636 40012 6692
rect 40068 6636 40078 6692
rect 34850 6524 34860 6580
rect 34916 6524 36428 6580
rect 36484 6524 36494 6580
rect 38882 6524 38892 6580
rect 38948 6524 39676 6580
rect 39732 6524 40348 6580
rect 40404 6524 40414 6580
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 44594 6076 44604 6132
rect 44660 6076 48020 6132
rect 47964 6020 48020 6076
rect 49200 6020 50000 6048
rect 46834 5964 46844 6020
rect 46900 5964 47740 6020
rect 47796 5964 47806 6020
rect 47964 5964 50000 6020
rect 49200 5936 50000 5964
rect 37538 5852 37548 5908
rect 37604 5852 38220 5908
rect 38276 5852 38892 5908
rect 38948 5852 38958 5908
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 3378 5180 3388 5236
rect 3444 5180 6524 5236
rect 6580 5180 6590 5236
rect 33954 5180 33964 5236
rect 34020 5180 35532 5236
rect 35588 5180 38332 5236
rect 38388 5180 38780 5236
rect 38836 5180 38846 5236
rect 5842 5068 5852 5124
rect 5908 5068 9212 5124
rect 9268 5068 9278 5124
rect 40338 5068 40348 5124
rect 40404 5068 44268 5124
rect 44324 5068 45500 5124
rect 45556 5068 45566 5124
rect 8642 4956 8652 5012
rect 8708 4956 14476 5012
rect 14532 4956 14542 5012
rect 35858 4956 35868 5012
rect 35924 4956 36764 5012
rect 36820 4956 37436 5012
rect 37492 4956 38444 5012
rect 38500 4956 38510 5012
rect 44146 4956 44156 5012
rect 44212 4956 46956 5012
rect 47012 4956 47516 5012
rect 47572 4956 47582 5012
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 46610 4620 46620 4676
rect 46676 4620 48020 4676
rect 47964 4564 48020 4620
rect 49200 4564 50000 4592
rect 44594 4508 44604 4564
rect 44660 4508 47292 4564
rect 47348 4508 47358 4564
rect 47964 4508 50000 4564
rect 49200 4480 50000 4508
rect 36194 4396 36204 4452
rect 36260 4396 37548 4452
rect 37604 4396 37614 4452
rect 2930 4172 2940 4228
rect 2996 4172 26236 4228
rect 26292 4172 26302 4228
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 38434 3500 38444 3556
rect 38500 3500 44268 3556
rect 44324 3500 44940 3556
rect 44996 3500 45006 3556
rect 0 3444 800 3472
rect 0 3388 1932 3444
rect 1988 3388 1998 3444
rect 0 3360 800 3388
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 49200 3108 50000 3136
rect 46050 3052 46060 3108
rect 46116 3052 50000 3108
rect 49200 3024 50000 3052
rect 49200 1652 50000 1680
rect 45042 1596 45052 1652
rect 45108 1596 50000 1652
rect 49200 1568 50000 1596
<< via3 >>
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 46284 4768 46316
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 45500 20128 46316
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 46284 35488 46316
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__078__A2 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 25760 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__081__A2
timestamp 1669390400
transform 1 0 20944 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__082__I
timestamp 1669390400
transform 1 0 37856 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__083__I
timestamp 1669390400
transform -1 0 39760 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__084__I0
timestamp 1669390400
transform 1 0 34832 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__084__I1
timestamp 1669390400
transform 1 0 37408 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__086__I0
timestamp 1669390400
transform 1 0 38416 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__086__I1
timestamp 1669390400
transform 1 0 38864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__088__I0
timestamp 1669390400
transform -1 0 40432 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__090__I1
timestamp 1669390400
transform 1 0 41104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__092__I
timestamp 1669390400
transform 1 0 43568 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__093__I0
timestamp 1669390400
transform -1 0 44912 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__101__I
timestamp 1669390400
transform 1 0 41776 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__110__I
timestamp 1669390400
transform 1 0 43232 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__119__I
timestamp 1669390400
transform 1 0 39760 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__120__I
timestamp 1669390400
transform 1 0 40768 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__129__I
timestamp 1669390400
transform 1 0 42448 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__130__S
timestamp 1669390400
transform 1 0 47488 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__132__S
timestamp 1669390400
transform 1 0 47600 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__134__S
timestamp 1669390400
transform 1 0 47600 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__136__I1
timestamp 1669390400
transform 1 0 48048 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__136__S
timestamp 1669390400
transform 1 0 47600 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__138__I
timestamp 1669390400
transform 1 0 41440 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__139__I0
timestamp 1669390400
transform 1 0 43456 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__141__I1
timestamp 1669390400
transform 1 0 43344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__143__I0
timestamp 1669390400
transform 1 0 42336 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__143__I1
timestamp 1669390400
transform 1 0 39424 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__145__I0
timestamp 1669390400
transform 1 0 39872 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__145__I1
timestamp 1669390400
transform -1 0 36960 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__147__I
timestamp 1669390400
transform 1 0 39872 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__148__I0
timestamp 1669390400
transform 1 0 38304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__148__I1
timestamp 1669390400
transform 1 0 39648 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__150__I0
timestamp 1669390400
transform -1 0 36960 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__150__I1
timestamp 1669390400
transform 1 0 39200 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__152__I0
timestamp 1669390400
transform 1 0 35168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__152__I1
timestamp 1669390400
transform 1 0 35616 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__154__I0
timestamp 1669390400
transform 1 0 34832 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__154__I1
timestamp 1669390400
transform -1 0 32928 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__156__CLK
timestamp 1669390400
transform 1 0 9632 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__157__CLK
timestamp 1669390400
transform 1 0 16688 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__158__CLK
timestamp 1669390400
transform 1 0 21728 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__158__D
timestamp 1669390400
transform 1 0 21728 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__159__CLK
timestamp 1669390400
transform 1 0 8960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__160__CLK
timestamp 1669390400
transform 1 0 14336 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__160__D
timestamp 1669390400
transform 1 0 10416 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__161__CLK
timestamp 1669390400
transform -1 0 20384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__162__CLK
timestamp 1669390400
transform -1 0 9296 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__163__CLK
timestamp 1669390400
transform 1 0 17024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__164__CLK
timestamp 1669390400
transform 1 0 22736 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__164__D
timestamp 1669390400
transform 1 0 18816 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__165__CLK
timestamp 1669390400
transform 1 0 38304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__166__CLK
timestamp 1669390400
transform 1 0 38752 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__167__CLK
timestamp 1669390400
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__168__CLK
timestamp 1669390400
transform 1 0 37632 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__169__CLK
timestamp 1669390400
transform 1 0 44128 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__170__CLK
timestamp 1669390400
transform 1 0 43792 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__171__CLK
timestamp 1669390400
transform 1 0 42336 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__172__CLK
timestamp 1669390400
transform 1 0 43232 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__173__CLK
timestamp 1669390400
transform 1 0 41216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__174__CLK
timestamp 1669390400
transform 1 0 40544 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__175__CLK
timestamp 1669390400
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__176__CLK
timestamp 1669390400
transform 1 0 43120 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__177__CLK
timestamp 1669390400
transform 1 0 43344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__178__CLK
timestamp 1669390400
transform 1 0 42224 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__179__CLK
timestamp 1669390400
transform 1 0 43904 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__180__CLK
timestamp 1669390400
transform 1 0 41216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__181__CLK
timestamp 1669390400
transform 1 0 42784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__182__CLK
timestamp 1669390400
transform 1 0 40096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__183__CLK
timestamp 1669390400
transform 1 0 43232 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__184__CLK
timestamp 1669390400
transform 1 0 43232 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__185__CLK
timestamp 1669390400
transform 1 0 43344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__186__CLK
timestamp 1669390400
transform 1 0 43792 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__187__CLK
timestamp 1669390400
transform -1 0 43904 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__188__CLK
timestamp 1669390400
transform 1 0 42224 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__189__CLK
timestamp 1669390400
transform 1 0 40768 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__190__CLK
timestamp 1669390400
transform 1 0 39200 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__191__CLK
timestamp 1669390400
transform -1 0 36288 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__192__CLK
timestamp 1669390400
transform 1 0 38752 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__193__CLK
timestamp 1669390400
transform 1 0 36736 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__194__CLK
timestamp 1669390400
transform 1 0 34832 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__195__CLK
timestamp 1669390400
transform 1 0 34608 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__196__CLK
timestamp 1669390400
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__205__I
timestamp 1669390400
transform 1 0 46928 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__I
timestamp 1669390400
transform 1 0 4032 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clock_I
timestamp 1669390400
transform -1 0 26432 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_0__f_clock_I
timestamp 1669390400
transform 1 0 33712 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_1__f_clock_I
timestamp 1669390400
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_2__f_clock_I
timestamp 1669390400
transform 1 0 33712 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_3__f_clock_I
timestamp 1669390400
transform 1 0 29904 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1669390400
transform -1 0 1904 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1669390400
transform -1 0 1904 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1669390400
transform -1 0 1904 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output5_I
timestamp 1669390400
transform -1 0 44352 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output16_I
timestamp 1669390400
transform 1 0 44240 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output20_I
timestamp 1669390400
transform 1 0 47152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output22_I
timestamp 1669390400
transform 1 0 44688 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output23_I
timestamp 1669390400
transform 1 0 44688 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output24_I
timestamp 1669390400
transform 1 0 44688 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output25_I
timestamp 1669390400
transform 1 0 44688 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output26_I
timestamp 1669390400
transform 1 0 44128 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output28_I
timestamp 1669390400
transform -1 0 44576 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output29_I
timestamp 1669390400
transform 1 0 46592 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output30_I
timestamp 1669390400
transform 1 0 42896 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1568 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 3472 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37
timestamp 1669390400
transform 1 0 5488 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 7280 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 8176 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63
timestamp 1669390400
transform 1 0 8400 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68
timestamp 1669390400
transform 1 0 8960 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_72 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 9408 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1669390400
transform 1 0 12992 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_107 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 13328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_111
timestamp 1669390400
transform 1 0 13776 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_117
timestamp 1669390400
transform 1 0 14448 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_133
timestamp 1669390400
transform 1 0 16240 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_137
timestamp 1669390400
transform 1 0 16688 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_139
timestamp 1669390400
transform 1 0 16912 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_142
timestamp 1669390400
transform 1 0 17248 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_158
timestamp 1669390400
transform 1 0 19040 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_166
timestamp 1669390400
transform 1 0 19936 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_174
timestamp 1669390400
transform 1 0 20832 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_177
timestamp 1669390400
transform 1 0 21168 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_209
timestamp 1669390400
transform 1 0 24752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_212
timestamp 1669390400
transform 1 0 25088 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_217
timestamp 1669390400
transform 1 0 25648 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_233
timestamp 1669390400
transform 1 0 27440 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_241
timestamp 1669390400
transform 1 0 28336 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_247
timestamp 1669390400
transform 1 0 29008 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_279
timestamp 1669390400
transform 1 0 32592 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_282
timestamp 1669390400
transform 1 0 32928 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_314
timestamp 1669390400
transform 1 0 36512 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_317
timestamp 1669390400
transform 1 0 36848 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_349
timestamp 1669390400
transform 1 0 40432 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_352
timestamp 1669390400
transform 1 0 40768 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_368
timestamp 1669390400
transform 1 0 42560 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_376
timestamp 1669390400
transform 1 0 43456 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_380
timestamp 1669390400
transform 1 0 43904 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_384
timestamp 1669390400
transform 1 0 44352 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_387
timestamp 1669390400
transform 1 0 44688 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_402
timestamp 1669390400
transform 1 0 46368 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_418
timestamp 1669390400
transform 1 0 48160 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_2
timestamp 1669390400
transform 1 0 1568 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_5 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1904 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_69
timestamp 1669390400
transform 1 0 9072 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_73
timestamp 1669390400
transform 1 0 9520 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_137
timestamp 1669390400
transform 1 0 16688 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_141
timestamp 1669390400
transform 1 0 17136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_144
timestamp 1669390400
transform 1 0 17472 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_208
timestamp 1669390400
transform 1 0 24640 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_212
timestamp 1669390400
transform 1 0 25088 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_215
timestamp 1669390400
transform 1 0 25424 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_279
timestamp 1669390400
transform 1 0 32592 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_283
timestamp 1669390400
transform 1 0 33040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_286
timestamp 1669390400
transform 1 0 33376 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_302
timestamp 1669390400
transform 1 0 35168 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_332
timestamp 1669390400
transform 1 0 38528 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_336
timestamp 1669390400
transform 1 0 38976 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_352
timestamp 1669390400
transform 1 0 40768 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_354
timestamp 1669390400
transform 1 0 40992 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_357
timestamp 1669390400
transform 1 0 41328 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_373
timestamp 1669390400
transform 1 0 43120 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_381
timestamp 1669390400
transform 1 0 44016 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_391
timestamp 1669390400
transform 1 0 45136 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_409
timestamp 1669390400
transform 1 0 47152 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_417
timestamp 1669390400
transform 1 0 48048 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_419
timestamp 1669390400
transform 1 0 48272 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_2
timestamp 1669390400
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1669390400
transform 1 0 5152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_37
timestamp 1669390400
transform 1 0 5488 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_67
timestamp 1669390400
transform 1 0 8848 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_71
timestamp 1669390400
transform 1 0 9296 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_103
timestamp 1669390400
transform 1 0 12880 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1669390400
transform 1 0 13104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_108
timestamp 1669390400
transform 1 0 13440 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_172
timestamp 1669390400
transform 1 0 20608 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_176
timestamp 1669390400
transform 1 0 21056 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_179
timestamp 1669390400
transform 1 0 21392 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_243
timestamp 1669390400
transform 1 0 28560 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_247
timestamp 1669390400
transform 1 0 29008 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_250
timestamp 1669390400
transform 1 0 29344 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_282
timestamp 1669390400
transform 1 0 32928 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_286
timestamp 1669390400
transform 1 0 33376 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_288
timestamp 1669390400
transform 1 0 33600 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_318
timestamp 1669390400
transform 1 0 36960 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_321
timestamp 1669390400
transform 1 0 37296 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_328
timestamp 1669390400
transform 1 0 38080 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_332
timestamp 1669390400
transform 1 0 38528 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_364
timestamp 1669390400
transform 1 0 42112 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_380
timestamp 1669390400
transform 1 0 43904 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_382
timestamp 1669390400
transform 1 0 44128 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_385
timestamp 1669390400
transform 1 0 44464 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_389
timestamp 1669390400
transform 1 0 44912 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_392
timestamp 1669390400
transform 1 0 45248 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_407
timestamp 1669390400
transform 1 0 46928 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_415
timestamp 1669390400
transform 1 0 47824 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_419
timestamp 1669390400
transform 1 0 48272 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_2
timestamp 1669390400
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_66
timestamp 1669390400
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1669390400
transform 1 0 9184 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_73
timestamp 1669390400
transform 1 0 9520 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_137
timestamp 1669390400
transform 1 0 16688 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_141
timestamp 1669390400
transform 1 0 17136 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_144
timestamp 1669390400
transform 1 0 17472 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_208
timestamp 1669390400
transform 1 0 24640 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_212
timestamp 1669390400
transform 1 0 25088 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_215
timestamp 1669390400
transform 1 0 25424 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_279
timestamp 1669390400
transform 1 0 32592 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_283
timestamp 1669390400
transform 1 0 33040 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_286
timestamp 1669390400
transform 1 0 33376 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_294
timestamp 1669390400
transform 1 0 34272 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_298
timestamp 1669390400
transform 1 0 34720 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_306
timestamp 1669390400
transform 1 0 35616 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_329
timestamp 1669390400
transform 1 0 38192 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_333
timestamp 1669390400
transform 1 0 38640 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_337
timestamp 1669390400
transform 1 0 39088 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_353
timestamp 1669390400
transform 1 0 40880 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_357
timestamp 1669390400
transform 1 0 41328 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_373
timestamp 1669390400
transform 1 0 43120 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_381
timestamp 1669390400
transform 1 0 44016 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_384
timestamp 1669390400
transform 1 0 44352 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_415
timestamp 1669390400
transform 1 0 47824 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_419
timestamp 1669390400
transform 1 0 48272 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_2
timestamp 1669390400
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1669390400
transform 1 0 5152 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_37
timestamp 1669390400
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_101
timestamp 1669390400
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1669390400
transform 1 0 13104 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_108
timestamp 1669390400
transform 1 0 13440 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_172
timestamp 1669390400
transform 1 0 20608 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_176
timestamp 1669390400
transform 1 0 21056 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_179
timestamp 1669390400
transform 1 0 21392 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_243
timestamp 1669390400
transform 1 0 28560 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_247
timestamp 1669390400
transform 1 0 29008 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_250
timestamp 1669390400
transform 1 0 29344 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_282
timestamp 1669390400
transform 1 0 32928 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_298
timestamp 1669390400
transform 1 0 34720 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_301
timestamp 1669390400
transform 1 0 35056 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_318
timestamp 1669390400
transform 1 0 36960 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_321
timestamp 1669390400
transform 1 0 37296 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_324
timestamp 1669390400
transform 1 0 37632 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_328
timestamp 1669390400
transform 1 0 38080 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_345
timestamp 1669390400
transform 1 0 39984 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_349
timestamp 1669390400
transform 1 0 40432 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_365
timestamp 1669390400
transform 1 0 42224 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_373
timestamp 1669390400
transform 1 0 43120 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_389
timestamp 1669390400
transform 1 0 44912 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_392
timestamp 1669390400
transform 1 0 45248 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_411
timestamp 1669390400
transform 1 0 47376 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_419
timestamp 1669390400
transform 1 0 48272 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_2
timestamp 1669390400
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_66
timestamp 1669390400
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1669390400
transform 1 0 9184 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_73
timestamp 1669390400
transform 1 0 9520 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_137
timestamp 1669390400
transform 1 0 16688 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_141
timestamp 1669390400
transform 1 0 17136 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_144
timestamp 1669390400
transform 1 0 17472 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_176
timestamp 1669390400
transform 1 0 21056 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_180
timestamp 1669390400
transform 1 0 21504 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_184
timestamp 1669390400
transform 1 0 21952 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_200
timestamp 1669390400
transform 1 0 23744 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_208
timestamp 1669390400
transform 1 0 24640 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_212
timestamp 1669390400
transform 1 0 25088 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_215
timestamp 1669390400
transform 1 0 25424 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_218
timestamp 1669390400
transform 1 0 25760 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_282
timestamp 1669390400
transform 1 0 32928 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_286
timestamp 1669390400
transform 1 0 33376 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_318
timestamp 1669390400
transform 1 0 36960 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_348
timestamp 1669390400
transform 1 0 40320 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_352
timestamp 1669390400
transform 1 0 40768 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_354
timestamp 1669390400
transform 1 0 40992 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_357
timestamp 1669390400
transform 1 0 41328 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_373
timestamp 1669390400
transform 1 0 43120 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_377
timestamp 1669390400
transform 1 0 43568 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_381
timestamp 1669390400
transform 1 0 44016 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_412
timestamp 1669390400
transform 1 0 47488 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1669390400
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1669390400
transform 1 0 5152 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_37
timestamp 1669390400
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_101
timestamp 1669390400
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_105
timestamp 1669390400
transform 1 0 13104 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_108
timestamp 1669390400
transform 1 0 13440 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_138
timestamp 1669390400
transform 1 0 16800 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_142
timestamp 1669390400
transform 1 0 17248 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_174
timestamp 1669390400
transform 1 0 20832 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_176
timestamp 1669390400
transform 1 0 21056 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_179
timestamp 1669390400
transform 1 0 21392 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_181
timestamp 1669390400
transform 1 0 21616 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_184
timestamp 1669390400
transform 1 0 21952 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_215
timestamp 1669390400
transform 1 0 25424 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_225
timestamp 1669390400
transform 1 0 26544 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_241
timestamp 1669390400
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_245
timestamp 1669390400
transform 1 0 28784 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_247
timestamp 1669390400
transform 1 0 29008 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_250
timestamp 1669390400
transform 1 0 29344 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_314
timestamp 1669390400
transform 1 0 36512 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_318
timestamp 1669390400
transform 1 0 36960 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_321
timestamp 1669390400
transform 1 0 37296 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_325
timestamp 1669390400
transform 1 0 37744 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_332
timestamp 1669390400
transform 1 0 38528 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_336
timestamp 1669390400
transform 1 0 38976 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_353
timestamp 1669390400
transform 1 0 40880 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_357
timestamp 1669390400
transform 1 0 41328 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_365
timestamp 1669390400
transform 1 0 42224 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_369
timestamp 1669390400
transform 1 0 42672 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_373
timestamp 1669390400
transform 1 0 43120 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_389
timestamp 1669390400
transform 1 0 44912 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_392
timestamp 1669390400
transform 1 0 45248 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_411
timestamp 1669390400
transform 1 0 47376 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_419
timestamp 1669390400
transform 1 0 48272 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_2
timestamp 1669390400
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_66
timestamp 1669390400
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_70
timestamp 1669390400
transform 1 0 9184 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_73
timestamp 1669390400
transform 1 0 9520 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_137
timestamp 1669390400
transform 1 0 16688 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_141
timestamp 1669390400
transform 1 0 17136 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_144
timestamp 1669390400
transform 1 0 17472 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_208
timestamp 1669390400
transform 1 0 24640 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_212
timestamp 1669390400
transform 1 0 25088 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_215
timestamp 1669390400
transform 1 0 25424 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_279
timestamp 1669390400
transform 1 0 32592 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_283
timestamp 1669390400
transform 1 0 33040 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_286
timestamp 1669390400
transform 1 0 33376 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_318
timestamp 1669390400
transform 1 0 36960 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_326
timestamp 1669390400
transform 1 0 37856 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_330
timestamp 1669390400
transform 1 0 38304 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_339
timestamp 1669390400
transform 1 0 39312 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_343
timestamp 1669390400
transform 1 0 39760 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_351
timestamp 1669390400
transform 1 0 40656 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_357
timestamp 1669390400
transform 1 0 41328 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_373
timestamp 1669390400
transform 1 0 43120 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_381
timestamp 1669390400
transform 1 0 44016 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_385
timestamp 1669390400
transform 1 0 44464 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_387
timestamp 1669390400
transform 1 0 44688 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_402
timestamp 1669390400
transform 1 0 46368 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_410
timestamp 1669390400
transform 1 0 47264 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_418
timestamp 1669390400
transform 1 0 48160 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_2
timestamp 1669390400
transform 1 0 1568 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_7
timestamp 1669390400
transform 1 0 2128 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_23
timestamp 1669390400
transform 1 0 3920 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_31
timestamp 1669390400
transform 1 0 4816 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_37
timestamp 1669390400
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_101
timestamp 1669390400
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1669390400
transform 1 0 13104 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_108
timestamp 1669390400
transform 1 0 13440 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_172
timestamp 1669390400
transform 1 0 20608 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_176
timestamp 1669390400
transform 1 0 21056 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_179
timestamp 1669390400
transform 1 0 21392 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_243
timestamp 1669390400
transform 1 0 28560 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_247
timestamp 1669390400
transform 1 0 29008 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_250
timestamp 1669390400
transform 1 0 29344 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_314
timestamp 1669390400
transform 1 0 36512 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_318
timestamp 1669390400
transform 1 0 36960 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_321
timestamp 1669390400
transform 1 0 37296 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_323
timestamp 1669390400
transform 1 0 37520 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_326
timestamp 1669390400
transform 1 0 37856 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_357
timestamp 1669390400
transform 1 0 41328 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_373
timestamp 1669390400
transform 1 0 43120 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_379
timestamp 1669390400
transform 1 0 43792 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_389
timestamp 1669390400
transform 1 0 44912 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_392
timestamp 1669390400
transform 1 0 45248 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_407
timestamp 1669390400
transform 1 0 46928 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_415
timestamp 1669390400
transform 1 0 47824 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_419
timestamp 1669390400
transform 1 0 48272 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_2
timestamp 1669390400
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_66
timestamp 1669390400
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_70
timestamp 1669390400
transform 1 0 9184 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_73
timestamp 1669390400
transform 1 0 9520 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_137
timestamp 1669390400
transform 1 0 16688 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_141
timestamp 1669390400
transform 1 0 17136 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_144
timestamp 1669390400
transform 1 0 17472 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_208
timestamp 1669390400
transform 1 0 24640 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_212
timestamp 1669390400
transform 1 0 25088 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_215
timestamp 1669390400
transform 1 0 25424 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_279
timestamp 1669390400
transform 1 0 32592 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_283
timestamp 1669390400
transform 1 0 33040 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_286
timestamp 1669390400
transform 1 0 33376 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_318
timestamp 1669390400
transform 1 0 36960 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_334
timestamp 1669390400
transform 1 0 38752 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_342
timestamp 1669390400
transform 1 0 39648 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_350
timestamp 1669390400
transform 1 0 40544 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_354
timestamp 1669390400
transform 1 0 40992 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_357
timestamp 1669390400
transform 1 0 41328 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_365
timestamp 1669390400
transform 1 0 42224 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_368
timestamp 1669390400
transform 1 0 42560 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_399
timestamp 1669390400
transform 1 0 46032 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_416
timestamp 1669390400
transform 1 0 47936 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_2
timestamp 1669390400
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1669390400
transform 1 0 5152 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_37
timestamp 1669390400
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_101
timestamp 1669390400
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1669390400
transform 1 0 13104 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_108
timestamp 1669390400
transform 1 0 13440 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_172
timestamp 1669390400
transform 1 0 20608 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_176
timestamp 1669390400
transform 1 0 21056 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_179
timestamp 1669390400
transform 1 0 21392 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_243
timestamp 1669390400
transform 1 0 28560 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_247
timestamp 1669390400
transform 1 0 29008 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_250
timestamp 1669390400
transform 1 0 29344 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_314
timestamp 1669390400
transform 1 0 36512 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_318
timestamp 1669390400
transform 1 0 36960 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_321
timestamp 1669390400
transform 1 0 37296 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_353
timestamp 1669390400
transform 1 0 40880 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_369
timestamp 1669390400
transform 1 0 42672 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_373
timestamp 1669390400
transform 1 0 43120 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_381
timestamp 1669390400
transform 1 0 44016 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_389
timestamp 1669390400
transform 1 0 44912 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_392
timestamp 1669390400
transform 1 0 45248 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_408
timestamp 1669390400
transform 1 0 47040 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_416
timestamp 1669390400
transform 1 0 47936 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_2
timestamp 1669390400
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_66
timestamp 1669390400
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_70
timestamp 1669390400
transform 1 0 9184 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_73
timestamp 1669390400
transform 1 0 9520 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_105
timestamp 1669390400
transform 1 0 13104 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_135
timestamp 1669390400
transform 1 0 16464 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_139
timestamp 1669390400
transform 1 0 16912 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_141
timestamp 1669390400
transform 1 0 17136 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_144
timestamp 1669390400
transform 1 0 17472 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_152
timestamp 1669390400
transform 1 0 18368 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_156
timestamp 1669390400
transform 1 0 18816 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_208
timestamp 1669390400
transform 1 0 24640 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_212
timestamp 1669390400
transform 1 0 25088 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_215
timestamp 1669390400
transform 1 0 25424 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_279
timestamp 1669390400
transform 1 0 32592 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_283
timestamp 1669390400
transform 1 0 33040 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_286
timestamp 1669390400
transform 1 0 33376 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_288
timestamp 1669390400
transform 1 0 33600 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_291
timestamp 1669390400
transform 1 0 33936 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_343
timestamp 1669390400
transform 1 0 39760 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_351
timestamp 1669390400
transform 1 0 40656 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_357
timestamp 1669390400
transform 1 0 41328 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_373
timestamp 1669390400
transform 1 0 43120 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_376
timestamp 1669390400
transform 1 0 43456 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_407
timestamp 1669390400
transform 1 0 46928 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_415
timestamp 1669390400
transform 1 0 47824 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_419
timestamp 1669390400
transform 1 0 48272 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_2
timestamp 1669390400
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1669390400
transform 1 0 5152 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_37
timestamp 1669390400
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_101
timestamp 1669390400
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_105
timestamp 1669390400
transform 1 0 13104 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_108
timestamp 1669390400
transform 1 0 13440 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_172
timestamp 1669390400
transform 1 0 20608 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_176
timestamp 1669390400
transform 1 0 21056 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_179
timestamp 1669390400
transform 1 0 21392 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_243
timestamp 1669390400
transform 1 0 28560 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_247
timestamp 1669390400
transform 1 0 29008 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_250
timestamp 1669390400
transform 1 0 29344 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_314
timestamp 1669390400
transform 1 0 36512 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_318
timestamp 1669390400
transform 1 0 36960 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_321
timestamp 1669390400
transform 1 0 37296 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_385
timestamp 1669390400
transform 1 0 44464 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_389
timestamp 1669390400
transform 1 0 44912 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_392
timestamp 1669390400
transform 1 0 45248 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_407
timestamp 1669390400
transform 1 0 46928 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_415
timestamp 1669390400
transform 1 0 47824 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_419
timestamp 1669390400
transform 1 0 48272 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_2
timestamp 1669390400
transform 1 0 1568 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_34
timestamp 1669390400
transform 1 0 5152 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_38
timestamp 1669390400
transform 1 0 5600 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_40
timestamp 1669390400
transform 1 0 5824 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_70
timestamp 1669390400
transform 1 0 9184 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_73
timestamp 1669390400
transform 1 0 9520 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_76
timestamp 1669390400
transform 1 0 9856 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_80
timestamp 1669390400
transform 1 0 10304 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_83
timestamp 1669390400
transform 1 0 10640 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_114
timestamp 1669390400
transform 1 0 14112 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_118
timestamp 1669390400
transform 1 0 14560 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_134
timestamp 1669390400
transform 1 0 16352 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_144
timestamp 1669390400
transform 1 0 17472 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_152
timestamp 1669390400
transform 1 0 18368 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_158
timestamp 1669390400
transform 1 0 19040 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_189
timestamp 1669390400
transform 1 0 22512 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_193
timestamp 1669390400
transform 1 0 22960 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_209
timestamp 1669390400
transform 1 0 24752 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_215
timestamp 1669390400
transform 1 0 25424 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_279
timestamp 1669390400
transform 1 0 32592 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_283
timestamp 1669390400
transform 1 0 33040 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_286
timestamp 1669390400
transform 1 0 33376 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_350
timestamp 1669390400
transform 1 0 40544 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_354
timestamp 1669390400
transform 1 0 40992 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_357
timestamp 1669390400
transform 1 0 41328 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_373
timestamp 1669390400
transform 1 0 43120 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_381
timestamp 1669390400
transform 1 0 44016 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_385
timestamp 1669390400
transform 1 0 44464 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_387
timestamp 1669390400
transform 1 0 44688 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_402
timestamp 1669390400
transform 1 0 46368 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_418
timestamp 1669390400
transform 1 0 48160 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_2
timestamp 1669390400
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_34
timestamp 1669390400
transform 1 0 5152 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_37
timestamp 1669390400
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_101
timestamp 1669390400
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_105
timestamp 1669390400
transform 1 0 13104 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_108
timestamp 1669390400
transform 1 0 13440 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_124
timestamp 1669390400
transform 1 0 15232 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_132
timestamp 1669390400
transform 1 0 16128 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_136
timestamp 1669390400
transform 1 0 16576 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_138
timestamp 1669390400
transform 1 0 16800 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_168
timestamp 1669390400
transform 1 0 20160 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_175
timestamp 1669390400
transform 1 0 20944 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_179
timestamp 1669390400
transform 1 0 21392 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_183
timestamp 1669390400
transform 1 0 21840 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_188
timestamp 1669390400
transform 1 0 22400 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_220
timestamp 1669390400
transform 1 0 25984 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_236
timestamp 1669390400
transform 1 0 27776 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_244
timestamp 1669390400
transform 1 0 28672 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_250
timestamp 1669390400
transform 1 0 29344 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_314
timestamp 1669390400
transform 1 0 36512 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_318
timestamp 1669390400
transform 1 0 36960 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_321
timestamp 1669390400
transform 1 0 37296 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_353
timestamp 1669390400
transform 1 0 40880 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_355
timestamp 1669390400
transform 1 0 41104 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_358
timestamp 1669390400
transform 1 0 41440 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_389
timestamp 1669390400
transform 1 0 44912 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_392
timestamp 1669390400
transform 1 0 45248 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_408
timestamp 1669390400
transform 1 0 47040 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_416
timestamp 1669390400
transform 1 0 47936 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_2
timestamp 1669390400
transform 1 0 1568 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_5
timestamp 1669390400
transform 1 0 1904 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_69
timestamp 1669390400
transform 1 0 9072 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_73
timestamp 1669390400
transform 1 0 9520 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_137
timestamp 1669390400
transform 1 0 16688 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_141
timestamp 1669390400
transform 1 0 17136 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_144
timestamp 1669390400
transform 1 0 17472 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_160
timestamp 1669390400
transform 1 0 19264 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_170
timestamp 1669390400
transform 1 0 20384 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_174
timestamp 1669390400
transform 1 0 20832 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_177
timestamp 1669390400
transform 1 0 21168 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_186
timestamp 1669390400
transform 1 0 22176 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_202
timestamp 1669390400
transform 1 0 23968 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_210
timestamp 1669390400
transform 1 0 24864 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_212
timestamp 1669390400
transform 1 0 25088 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_215
timestamp 1669390400
transform 1 0 25424 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_279
timestamp 1669390400
transform 1 0 32592 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_283
timestamp 1669390400
transform 1 0 33040 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_286
timestamp 1669390400
transform 1 0 33376 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_350
timestamp 1669390400
transform 1 0 40544 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_354
timestamp 1669390400
transform 1 0 40992 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_357
timestamp 1669390400
transform 1 0 41328 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_365
timestamp 1669390400
transform 1 0 42224 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_372
timestamp 1669390400
transform 1 0 43008 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_380
timestamp 1669390400
transform 1 0 43904 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_397
timestamp 1669390400
transform 1 0 45808 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_413
timestamp 1669390400
transform 1 0 47600 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_417
timestamp 1669390400
transform 1 0 48048 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_419
timestamp 1669390400
transform 1 0 48272 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_2
timestamp 1669390400
transform 1 0 1568 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_19
timestamp 1669390400
transform 1 0 3472 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_37
timestamp 1669390400
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_101
timestamp 1669390400
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_105
timestamp 1669390400
transform 1 0 13104 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_108
timestamp 1669390400
transform 1 0 13440 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_172
timestamp 1669390400
transform 1 0 20608 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_176
timestamp 1669390400
transform 1 0 21056 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_179
timestamp 1669390400
transform 1 0 21392 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_243
timestamp 1669390400
transform 1 0 28560 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_247
timestamp 1669390400
transform 1 0 29008 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_250
timestamp 1669390400
transform 1 0 29344 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_314
timestamp 1669390400
transform 1 0 36512 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_318
timestamp 1669390400
transform 1 0 36960 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_321
timestamp 1669390400
transform 1 0 37296 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_337
timestamp 1669390400
transform 1 0 39088 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_345
timestamp 1669390400
transform 1 0 39984 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_349
timestamp 1669390400
transform 1 0 40432 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_352
timestamp 1669390400
transform 1 0 40768 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_383
timestamp 1669390400
transform 1 0 44240 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_387
timestamp 1669390400
transform 1 0 44688 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_389
timestamp 1669390400
transform 1 0 44912 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_392
timestamp 1669390400
transform 1 0 45248 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_408
timestamp 1669390400
transform 1 0 47040 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_416
timestamp 1669390400
transform 1 0 47936 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_2
timestamp 1669390400
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_66
timestamp 1669390400
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_70
timestamp 1669390400
transform 1 0 9184 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_73
timestamp 1669390400
transform 1 0 9520 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_137
timestamp 1669390400
transform 1 0 16688 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_141
timestamp 1669390400
transform 1 0 17136 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_144
timestamp 1669390400
transform 1 0 17472 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_208
timestamp 1669390400
transform 1 0 24640 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_212
timestamp 1669390400
transform 1 0 25088 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_215
timestamp 1669390400
transform 1 0 25424 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_279
timestamp 1669390400
transform 1 0 32592 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_283
timestamp 1669390400
transform 1 0 33040 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_17_286
timestamp 1669390400
transform 1 0 33376 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_318
timestamp 1669390400
transform 1 0 36960 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_328
timestamp 1669390400
transform 1 0 38080 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_336
timestamp 1669390400
transform 1 0 38976 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_352
timestamp 1669390400
transform 1 0 40768 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_354
timestamp 1669390400
transform 1 0 40992 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_357
timestamp 1669390400
transform 1 0 41328 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_379
timestamp 1669390400
transform 1 0 43792 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_410
timestamp 1669390400
transform 1 0 47264 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_418
timestamp 1669390400
transform 1 0 48160 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_18_2
timestamp 1669390400
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_34
timestamp 1669390400
transform 1 0 5152 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_37
timestamp 1669390400
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_101
timestamp 1669390400
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_105
timestamp 1669390400
transform 1 0 13104 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_108
timestamp 1669390400
transform 1 0 13440 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_172
timestamp 1669390400
transform 1 0 20608 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_176
timestamp 1669390400
transform 1 0 21056 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_179
timestamp 1669390400
transform 1 0 21392 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_243
timestamp 1669390400
transform 1 0 28560 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_247
timestamp 1669390400
transform 1 0 29008 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_250
timestamp 1669390400
transform 1 0 29344 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_314
timestamp 1669390400
transform 1 0 36512 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_318
timestamp 1669390400
transform 1 0 36960 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_18_321
timestamp 1669390400
transform 1 0 37296 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_353
timestamp 1669390400
transform 1 0 40880 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_363
timestamp 1669390400
transform 1 0 42000 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_373
timestamp 1669390400
transform 1 0 43120 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_389
timestamp 1669390400
transform 1 0 44912 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_392
timestamp 1669390400
transform 1 0 45248 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_408
timestamp 1669390400
transform 1 0 47040 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_416
timestamp 1669390400
transform 1 0 47936 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_2
timestamp 1669390400
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_66
timestamp 1669390400
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_70
timestamp 1669390400
transform 1 0 9184 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_73
timestamp 1669390400
transform 1 0 9520 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_137
timestamp 1669390400
transform 1 0 16688 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_141
timestamp 1669390400
transform 1 0 17136 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_144
timestamp 1669390400
transform 1 0 17472 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_208
timestamp 1669390400
transform 1 0 24640 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_212
timestamp 1669390400
transform 1 0 25088 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_215
timestamp 1669390400
transform 1 0 25424 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_279
timestamp 1669390400
transform 1 0 32592 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_283
timestamp 1669390400
transform 1 0 33040 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_286
timestamp 1669390400
transform 1 0 33376 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_350
timestamp 1669390400
transform 1 0 40544 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_354
timestamp 1669390400
transform 1 0 40992 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_357
timestamp 1669390400
transform 1 0 41328 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_375
timestamp 1669390400
transform 1 0 43344 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_406
timestamp 1669390400
transform 1 0 46816 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_414
timestamp 1669390400
transform 1 0 47712 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_418
timestamp 1669390400
transform 1 0 48160 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_2
timestamp 1669390400
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_34
timestamp 1669390400
transform 1 0 5152 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_37
timestamp 1669390400
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_101
timestamp 1669390400
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_105
timestamp 1669390400
transform 1 0 13104 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_108
timestamp 1669390400
transform 1 0 13440 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_172
timestamp 1669390400
transform 1 0 20608 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_176
timestamp 1669390400
transform 1 0 21056 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_179
timestamp 1669390400
transform 1 0 21392 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_243
timestamp 1669390400
transform 1 0 28560 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_247
timestamp 1669390400
transform 1 0 29008 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_250
timestamp 1669390400
transform 1 0 29344 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_314
timestamp 1669390400
transform 1 0 36512 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_318
timestamp 1669390400
transform 1 0 36960 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_321
timestamp 1669390400
transform 1 0 37296 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_353
timestamp 1669390400
transform 1 0 40880 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_369
timestamp 1669390400
transform 1 0 42672 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_377
timestamp 1669390400
transform 1 0 43568 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_381
timestamp 1669390400
transform 1 0 44016 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_389
timestamp 1669390400
transform 1 0 44912 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_392
timestamp 1669390400
transform 1 0 45248 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_407
timestamp 1669390400
transform 1 0 46928 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_415
timestamp 1669390400
transform 1 0 47824 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_419
timestamp 1669390400
transform 1 0 48272 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_2
timestamp 1669390400
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_66
timestamp 1669390400
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_70
timestamp 1669390400
transform 1 0 9184 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_73
timestamp 1669390400
transform 1 0 9520 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_137
timestamp 1669390400
transform 1 0 16688 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_141
timestamp 1669390400
transform 1 0 17136 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_144
timestamp 1669390400
transform 1 0 17472 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_208
timestamp 1669390400
transform 1 0 24640 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_212
timestamp 1669390400
transform 1 0 25088 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_215
timestamp 1669390400
transform 1 0 25424 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_219
timestamp 1669390400
transform 1 0 25872 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_221
timestamp 1669390400
transform 1 0 26096 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_224
timestamp 1669390400
transform 1 0 26432 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_276
timestamp 1669390400
transform 1 0 32256 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_286
timestamp 1669390400
transform 1 0 33376 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_350
timestamp 1669390400
transform 1 0 40544 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_354
timestamp 1669390400
transform 1 0 40992 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_357
timestamp 1669390400
transform 1 0 41328 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_373
timestamp 1669390400
transform 1 0 43120 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_376
timestamp 1669390400
transform 1 0 43456 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_386
timestamp 1669390400
transform 1 0 44576 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_402
timestamp 1669390400
transform 1 0 46368 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_418
timestamp 1669390400
transform 1 0 48160 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_2
timestamp 1669390400
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_34
timestamp 1669390400
transform 1 0 5152 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_37
timestamp 1669390400
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_101
timestamp 1669390400
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_105
timestamp 1669390400
transform 1 0 13104 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_108
timestamp 1669390400
transform 1 0 13440 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_172
timestamp 1669390400
transform 1 0 20608 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_176
timestamp 1669390400
transform 1 0 21056 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_179
timestamp 1669390400
transform 1 0 21392 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_243
timestamp 1669390400
transform 1 0 28560 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_247
timestamp 1669390400
transform 1 0 29008 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_250
timestamp 1669390400
transform 1 0 29344 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_314
timestamp 1669390400
transform 1 0 36512 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_318
timestamp 1669390400
transform 1 0 36960 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_321
timestamp 1669390400
transform 1 0 37296 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_353
timestamp 1669390400
transform 1 0 40880 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_369
timestamp 1669390400
transform 1 0 42672 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_377
timestamp 1669390400
transform 1 0 43568 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_381
timestamp 1669390400
transform 1 0 44016 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_389
timestamp 1669390400
transform 1 0 44912 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_392
timestamp 1669390400
transform 1 0 45248 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_394
timestamp 1669390400
transform 1 0 45472 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_410
timestamp 1669390400
transform 1 0 47264 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_418
timestamp 1669390400
transform 1 0 48160 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_2
timestamp 1669390400
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_66
timestamp 1669390400
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_70
timestamp 1669390400
transform 1 0 9184 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_73
timestamp 1669390400
transform 1 0 9520 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_137
timestamp 1669390400
transform 1 0 16688 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_141
timestamp 1669390400
transform 1 0 17136 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_144
timestamp 1669390400
transform 1 0 17472 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_208
timestamp 1669390400
transform 1 0 24640 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_212
timestamp 1669390400
transform 1 0 25088 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_215
timestamp 1669390400
transform 1 0 25424 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_279
timestamp 1669390400
transform 1 0 32592 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_283
timestamp 1669390400
transform 1 0 33040 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_286
timestamp 1669390400
transform 1 0 33376 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_350
timestamp 1669390400
transform 1 0 40544 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_354
timestamp 1669390400
transform 1 0 40992 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_357
timestamp 1669390400
transform 1 0 41328 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_373
timestamp 1669390400
transform 1 0 43120 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_377
timestamp 1669390400
transform 1 0 43568 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_408
timestamp 1669390400
transform 1 0 47040 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_416
timestamp 1669390400
transform 1 0 47936 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_2
timestamp 1669390400
transform 1 0 1568 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_7
timestamp 1669390400
transform 1 0 2128 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_23
timestamp 1669390400
transform 1 0 3920 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_31
timestamp 1669390400
transform 1 0 4816 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_37
timestamp 1669390400
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_101
timestamp 1669390400
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_105
timestamp 1669390400
transform 1 0 13104 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_108
timestamp 1669390400
transform 1 0 13440 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_172
timestamp 1669390400
transform 1 0 20608 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_176
timestamp 1669390400
transform 1 0 21056 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_179
timestamp 1669390400
transform 1 0 21392 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_243
timestamp 1669390400
transform 1 0 28560 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_247
timestamp 1669390400
transform 1 0 29008 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_250
timestamp 1669390400
transform 1 0 29344 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_314
timestamp 1669390400
transform 1 0 36512 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_318
timestamp 1669390400
transform 1 0 36960 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_321
timestamp 1669390400
transform 1 0 37296 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_337
timestamp 1669390400
transform 1 0 39088 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_341
timestamp 1669390400
transform 1 0 39536 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_345
timestamp 1669390400
transform 1 0 39984 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_361
timestamp 1669390400
transform 1 0 41776 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_369
timestamp 1669390400
transform 1 0 42672 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_373
timestamp 1669390400
transform 1 0 43120 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_389
timestamp 1669390400
transform 1 0 44912 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_392
timestamp 1669390400
transform 1 0 45248 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_411
timestamp 1669390400
transform 1 0 47376 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_419
timestamp 1669390400
transform 1 0 48272 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_25_2
timestamp 1669390400
transform 1 0 1568 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_34
timestamp 1669390400
transform 1 0 5152 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_36
timestamp 1669390400
transform 1 0 5376 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_66
timestamp 1669390400
transform 1 0 8736 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_70
timestamp 1669390400
transform 1 0 9184 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_73
timestamp 1669390400
transform 1 0 9520 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_137
timestamp 1669390400
transform 1 0 16688 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_141
timestamp 1669390400
transform 1 0 17136 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_144
timestamp 1669390400
transform 1 0 17472 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_208
timestamp 1669390400
transform 1 0 24640 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_212
timestamp 1669390400
transform 1 0 25088 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_215
timestamp 1669390400
transform 1 0 25424 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_279
timestamp 1669390400
transform 1 0 32592 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_283
timestamp 1669390400
transform 1 0 33040 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_286
timestamp 1669390400
transform 1 0 33376 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_288
timestamp 1669390400
transform 1 0 33600 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_291
timestamp 1669390400
transform 1 0 33936 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_343
timestamp 1669390400
transform 1 0 39760 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_351
timestamp 1669390400
transform 1 0 40656 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_357
timestamp 1669390400
transform 1 0 41328 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_367
timestamp 1669390400
transform 1 0 42448 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_383
timestamp 1669390400
transform 1 0 44240 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_414
timestamp 1669390400
transform 1 0 47712 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_418
timestamp 1669390400
transform 1 0 48160 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_2
timestamp 1669390400
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_34
timestamp 1669390400
transform 1 0 5152 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_37
timestamp 1669390400
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_101
timestamp 1669390400
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_105
timestamp 1669390400
transform 1 0 13104 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_108
timestamp 1669390400
transform 1 0 13440 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_172
timestamp 1669390400
transform 1 0 20608 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_176
timestamp 1669390400
transform 1 0 21056 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_179
timestamp 1669390400
transform 1 0 21392 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_243
timestamp 1669390400
transform 1 0 28560 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_247
timestamp 1669390400
transform 1 0 29008 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_250
timestamp 1669390400
transform 1 0 29344 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_314
timestamp 1669390400
transform 1 0 36512 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_318
timestamp 1669390400
transform 1 0 36960 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_321
timestamp 1669390400
transform 1 0 37296 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_353
timestamp 1669390400
transform 1 0 40880 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_369
timestamp 1669390400
transform 1 0 42672 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_373
timestamp 1669390400
transform 1 0 43120 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_389
timestamp 1669390400
transform 1 0 44912 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_392
timestamp 1669390400
transform 1 0 45248 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_411
timestamp 1669390400
transform 1 0 47376 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_419
timestamp 1669390400
transform 1 0 48272 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_2
timestamp 1669390400
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_66
timestamp 1669390400
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_70
timestamp 1669390400
transform 1 0 9184 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_73
timestamp 1669390400
transform 1 0 9520 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_137
timestamp 1669390400
transform 1 0 16688 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_141
timestamp 1669390400
transform 1 0 17136 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_144
timestamp 1669390400
transform 1 0 17472 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_208
timestamp 1669390400
transform 1 0 24640 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_212
timestamp 1669390400
transform 1 0 25088 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_215
timestamp 1669390400
transform 1 0 25424 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_279
timestamp 1669390400
transform 1 0 32592 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_283
timestamp 1669390400
transform 1 0 33040 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_286
timestamp 1669390400
transform 1 0 33376 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_350
timestamp 1669390400
transform 1 0 40544 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_354
timestamp 1669390400
transform 1 0 40992 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_357
timestamp 1669390400
transform 1 0 41328 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_373
timestamp 1669390400
transform 1 0 43120 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_377
timestamp 1669390400
transform 1 0 43568 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_379
timestamp 1669390400
transform 1 0 43792 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_382
timestamp 1669390400
transform 1 0 44128 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_413
timestamp 1669390400
transform 1 0 47600 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_417
timestamp 1669390400
transform 1 0 48048 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_419
timestamp 1669390400
transform 1 0 48272 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_2
timestamp 1669390400
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_34
timestamp 1669390400
transform 1 0 5152 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_37
timestamp 1669390400
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_101
timestamp 1669390400
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_105
timestamp 1669390400
transform 1 0 13104 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_108
timestamp 1669390400
transform 1 0 13440 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_172
timestamp 1669390400
transform 1 0 20608 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_176
timestamp 1669390400
transform 1 0 21056 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_179
timestamp 1669390400
transform 1 0 21392 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_243
timestamp 1669390400
transform 1 0 28560 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_247
timestamp 1669390400
transform 1 0 29008 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_250
timestamp 1669390400
transform 1 0 29344 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_314
timestamp 1669390400
transform 1 0 36512 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_318
timestamp 1669390400
transform 1 0 36960 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_321
timestamp 1669390400
transform 1 0 37296 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_353
timestamp 1669390400
transform 1 0 40880 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_355
timestamp 1669390400
transform 1 0 41104 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_358
timestamp 1669390400
transform 1 0 41440 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_366
timestamp 1669390400
transform 1 0 42336 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_373
timestamp 1669390400
transform 1 0 43120 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_381
timestamp 1669390400
transform 1 0 44016 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_389
timestamp 1669390400
transform 1 0 44912 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_392
timestamp 1669390400
transform 1 0 45248 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_407
timestamp 1669390400
transform 1 0 46928 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_415
timestamp 1669390400
transform 1 0 47824 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_419
timestamp 1669390400
transform 1 0 48272 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_2
timestamp 1669390400
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_66
timestamp 1669390400
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_70
timestamp 1669390400
transform 1 0 9184 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_73
timestamp 1669390400
transform 1 0 9520 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_137
timestamp 1669390400
transform 1 0 16688 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_141
timestamp 1669390400
transform 1 0 17136 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_144
timestamp 1669390400
transform 1 0 17472 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_208
timestamp 1669390400
transform 1 0 24640 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_212
timestamp 1669390400
transform 1 0 25088 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_215
timestamp 1669390400
transform 1 0 25424 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_279
timestamp 1669390400
transform 1 0 32592 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_283
timestamp 1669390400
transform 1 0 33040 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_29_286
timestamp 1669390400
transform 1 0 33376 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_318
timestamp 1669390400
transform 1 0 36960 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_326
timestamp 1669390400
transform 1 0 37856 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_336
timestamp 1669390400
transform 1 0 38976 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_353
timestamp 1669390400
transform 1 0 40880 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_357
timestamp 1669390400
transform 1 0 41328 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_387
timestamp 1669390400
transform 1 0 44688 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_403
timestamp 1669390400
transform 1 0 46480 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_419
timestamp 1669390400
transform 1 0 48272 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_2
timestamp 1669390400
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_34
timestamp 1669390400
transform 1 0 5152 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_37
timestamp 1669390400
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_101
timestamp 1669390400
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_105
timestamp 1669390400
transform 1 0 13104 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_108
timestamp 1669390400
transform 1 0 13440 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_172
timestamp 1669390400
transform 1 0 20608 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_176
timestamp 1669390400
transform 1 0 21056 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_179
timestamp 1669390400
transform 1 0 21392 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_243
timestamp 1669390400
transform 1 0 28560 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_247
timestamp 1669390400
transform 1 0 29008 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_250
timestamp 1669390400
transform 1 0 29344 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_254
timestamp 1669390400
transform 1 0 29792 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_257
timestamp 1669390400
transform 1 0 30128 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_309
timestamp 1669390400
transform 1 0 35952 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_317
timestamp 1669390400
transform 1 0 36848 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_321
timestamp 1669390400
transform 1 0 37296 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_351
timestamp 1669390400
transform 1 0 40656 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_368
timestamp 1669390400
transform 1 0 42560 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_372
timestamp 1669390400
transform 1 0 43008 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_376
timestamp 1669390400
transform 1 0 43456 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_384
timestamp 1669390400
transform 1 0 44352 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_388
timestamp 1669390400
transform 1 0 44800 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_392
timestamp 1669390400
transform 1 0 45248 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_408
timestamp 1669390400
transform 1 0 47040 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_416
timestamp 1669390400
transform 1 0 47936 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_2
timestamp 1669390400
transform 1 0 1568 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_5
timestamp 1669390400
transform 1 0 1904 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_69
timestamp 1669390400
transform 1 0 9072 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_73
timestamp 1669390400
transform 1 0 9520 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_137
timestamp 1669390400
transform 1 0 16688 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_141
timestamp 1669390400
transform 1 0 17136 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_144
timestamp 1669390400
transform 1 0 17472 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_208
timestamp 1669390400
transform 1 0 24640 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_212
timestamp 1669390400
transform 1 0 25088 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_215
timestamp 1669390400
transform 1 0 25424 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_279
timestamp 1669390400
transform 1 0 32592 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_283
timestamp 1669390400
transform 1 0 33040 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_286
timestamp 1669390400
transform 1 0 33376 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_302
timestamp 1669390400
transform 1 0 35168 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_310
timestamp 1669390400
transform 1 0 36064 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_314
timestamp 1669390400
transform 1 0 36512 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_344
timestamp 1669390400
transform 1 0 39872 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_348
timestamp 1669390400
transform 1 0 40320 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_354
timestamp 1669390400
transform 1 0 40992 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_357
timestamp 1669390400
transform 1 0 41328 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_366
timestamp 1669390400
transform 1 0 42336 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_368
timestamp 1669390400
transform 1 0 42560 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_398
timestamp 1669390400
transform 1 0 45920 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_406
timestamp 1669390400
transform 1 0 46816 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_414
timestamp 1669390400
transform 1 0 47712 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_418
timestamp 1669390400
transform 1 0 48160 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_2
timestamp 1669390400
transform 1 0 1568 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_19
timestamp 1669390400
transform 1 0 3472 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_37
timestamp 1669390400
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_101
timestamp 1669390400
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_105
timestamp 1669390400
transform 1 0 13104 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_108
timestamp 1669390400
transform 1 0 13440 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_172
timestamp 1669390400
transform 1 0 20608 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_176
timestamp 1669390400
transform 1 0 21056 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_179
timestamp 1669390400
transform 1 0 21392 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_243
timestamp 1669390400
transform 1 0 28560 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_247
timestamp 1669390400
transform 1 0 29008 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_250
timestamp 1669390400
transform 1 0 29344 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_314
timestamp 1669390400
transform 1 0 36512 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_318
timestamp 1669390400
transform 1 0 36960 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_321
timestamp 1669390400
transform 1 0 37296 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_325
timestamp 1669390400
transform 1 0 37744 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_333
timestamp 1669390400
transform 1 0 38640 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_365
timestamp 1669390400
transform 1 0 42224 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_373
timestamp 1669390400
transform 1 0 43120 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_389
timestamp 1669390400
transform 1 0 44912 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_392
timestamp 1669390400
transform 1 0 45248 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_408
timestamp 1669390400
transform 1 0 47040 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_416
timestamp 1669390400
transform 1 0 47936 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_2
timestamp 1669390400
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_66
timestamp 1669390400
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_70
timestamp 1669390400
transform 1 0 9184 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_73
timestamp 1669390400
transform 1 0 9520 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_137
timestamp 1669390400
transform 1 0 16688 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_141
timestamp 1669390400
transform 1 0 17136 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_144
timestamp 1669390400
transform 1 0 17472 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_208
timestamp 1669390400
transform 1 0 24640 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_212
timestamp 1669390400
transform 1 0 25088 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_215
timestamp 1669390400
transform 1 0 25424 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_279
timestamp 1669390400
transform 1 0 32592 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_283
timestamp 1669390400
transform 1 0 33040 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_286
timestamp 1669390400
transform 1 0 33376 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_350
timestamp 1669390400
transform 1 0 40544 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_354
timestamp 1669390400
transform 1 0 40992 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_357
timestamp 1669390400
transform 1 0 41328 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_373
timestamp 1669390400
transform 1 0 43120 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_376
timestamp 1669390400
transform 1 0 43456 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_407
timestamp 1669390400
transform 1 0 46928 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_415
timestamp 1669390400
transform 1 0 47824 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_419
timestamp 1669390400
transform 1 0 48272 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_2
timestamp 1669390400
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_34
timestamp 1669390400
transform 1 0 5152 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_37
timestamp 1669390400
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_101
timestamp 1669390400
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_105
timestamp 1669390400
transform 1 0 13104 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_108
timestamp 1669390400
transform 1 0 13440 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_172
timestamp 1669390400
transform 1 0 20608 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_176
timestamp 1669390400
transform 1 0 21056 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_179
timestamp 1669390400
transform 1 0 21392 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_243
timestamp 1669390400
transform 1 0 28560 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_247
timestamp 1669390400
transform 1 0 29008 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_250
timestamp 1669390400
transform 1 0 29344 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_314
timestamp 1669390400
transform 1 0 36512 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_318
timestamp 1669390400
transform 1 0 36960 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_321
timestamp 1669390400
transform 1 0 37296 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_353
timestamp 1669390400
transform 1 0 40880 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_369
timestamp 1669390400
transform 1 0 42672 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_373
timestamp 1669390400
transform 1 0 43120 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_389
timestamp 1669390400
transform 1 0 44912 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_392
timestamp 1669390400
transform 1 0 45248 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_394
timestamp 1669390400
transform 1 0 45472 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_410
timestamp 1669390400
transform 1 0 47264 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_414
timestamp 1669390400
transform 1 0 47712 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_418
timestamp 1669390400
transform 1 0 48160 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_2
timestamp 1669390400
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_66
timestamp 1669390400
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_70
timestamp 1669390400
transform 1 0 9184 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_73
timestamp 1669390400
transform 1 0 9520 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_137
timestamp 1669390400
transform 1 0 16688 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_141
timestamp 1669390400
transform 1 0 17136 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_144
timestamp 1669390400
transform 1 0 17472 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_208
timestamp 1669390400
transform 1 0 24640 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_212
timestamp 1669390400
transform 1 0 25088 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_215
timestamp 1669390400
transform 1 0 25424 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_279
timestamp 1669390400
transform 1 0 32592 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_283
timestamp 1669390400
transform 1 0 33040 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_286
timestamp 1669390400
transform 1 0 33376 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_350
timestamp 1669390400
transform 1 0 40544 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_354
timestamp 1669390400
transform 1 0 40992 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_357
timestamp 1669390400
transform 1 0 41328 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_373
timestamp 1669390400
transform 1 0 43120 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_377
timestamp 1669390400
transform 1 0 43568 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_408
timestamp 1669390400
transform 1 0 47040 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_416
timestamp 1669390400
transform 1 0 47936 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_2
timestamp 1669390400
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_34
timestamp 1669390400
transform 1 0 5152 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_37
timestamp 1669390400
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_101
timestamp 1669390400
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_105
timestamp 1669390400
transform 1 0 13104 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_108
timestamp 1669390400
transform 1 0 13440 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_172
timestamp 1669390400
transform 1 0 20608 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_176
timestamp 1669390400
transform 1 0 21056 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_179
timestamp 1669390400
transform 1 0 21392 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_243
timestamp 1669390400
transform 1 0 28560 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_247
timestamp 1669390400
transform 1 0 29008 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_250
timestamp 1669390400
transform 1 0 29344 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_282
timestamp 1669390400
transform 1 0 32928 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_298
timestamp 1669390400
transform 1 0 34720 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_306
timestamp 1669390400
transform 1 0 35616 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_314
timestamp 1669390400
transform 1 0 36512 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_318
timestamp 1669390400
transform 1 0 36960 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_321
timestamp 1669390400
transform 1 0 37296 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_328
timestamp 1669390400
transform 1 0 38080 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_346
timestamp 1669390400
transform 1 0 40096 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_362
timestamp 1669390400
transform 1 0 41888 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_366
timestamp 1669390400
transform 1 0 42336 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_369
timestamp 1669390400
transform 1 0 42672 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_379
timestamp 1669390400
transform 1 0 43792 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_389
timestamp 1669390400
transform 1 0 44912 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_392
timestamp 1669390400
transform 1 0 45248 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_407
timestamp 1669390400
transform 1 0 46928 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_415
timestamp 1669390400
transform 1 0 47824 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_419
timestamp 1669390400
transform 1 0 48272 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_2
timestamp 1669390400
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_66
timestamp 1669390400
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_70
timestamp 1669390400
transform 1 0 9184 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_73
timestamp 1669390400
transform 1 0 9520 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_137
timestamp 1669390400
transform 1 0 16688 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_141
timestamp 1669390400
transform 1 0 17136 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_144
timestamp 1669390400
transform 1 0 17472 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_208
timestamp 1669390400
transform 1 0 24640 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_212
timestamp 1669390400
transform 1 0 25088 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_215
timestamp 1669390400
transform 1 0 25424 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_247
timestamp 1669390400
transform 1 0 29008 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_263
timestamp 1669390400
transform 1 0 30800 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_271
timestamp 1669390400
transform 1 0 31696 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_281
timestamp 1669390400
transform 1 0 32816 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_283
timestamp 1669390400
transform 1 0 33040 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_286
timestamp 1669390400
transform 1 0 33376 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_294
timestamp 1669390400
transform 1 0 34272 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_298
timestamp 1669390400
transform 1 0 34720 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_301
timestamp 1669390400
transform 1 0 35056 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_332
timestamp 1669390400
transform 1 0 38528 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_344
timestamp 1669390400
transform 1 0 39872 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_354
timestamp 1669390400
transform 1 0 40992 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_357
timestamp 1669390400
transform 1 0 41328 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_360
timestamp 1669390400
transform 1 0 41664 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_364
timestamp 1669390400
transform 1 0 42112 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_367
timestamp 1669390400
transform 1 0 42448 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_383
timestamp 1669390400
transform 1 0 44240 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_414
timestamp 1669390400
transform 1 0 47712 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_418
timestamp 1669390400
transform 1 0 48160 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_2
timestamp 1669390400
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_34
timestamp 1669390400
transform 1 0 5152 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_37
timestamp 1669390400
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_101
timestamp 1669390400
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_105
timestamp 1669390400
transform 1 0 13104 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_108
timestamp 1669390400
transform 1 0 13440 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_172
timestamp 1669390400
transform 1 0 20608 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_176
timestamp 1669390400
transform 1 0 21056 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_179
timestamp 1669390400
transform 1 0 21392 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_243
timestamp 1669390400
transform 1 0 28560 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_247
timestamp 1669390400
transform 1 0 29008 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_250
timestamp 1669390400
transform 1 0 29344 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_295
timestamp 1669390400
transform 1 0 34384 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_299
timestamp 1669390400
transform 1 0 34832 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_318
timestamp 1669390400
transform 1 0 36960 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_321
timestamp 1669390400
transform 1 0 37296 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_351
timestamp 1669390400
transform 1 0 40656 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_367
timestamp 1669390400
transform 1 0 42448 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_389
timestamp 1669390400
transform 1 0 44912 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_392
timestamp 1669390400
transform 1 0 45248 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_411
timestamp 1669390400
transform 1 0 47376 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_415
timestamp 1669390400
transform 1 0 47824 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_419
timestamp 1669390400
transform 1 0 48272 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_2
timestamp 1669390400
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_66
timestamp 1669390400
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_70
timestamp 1669390400
transform 1 0 9184 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_73
timestamp 1669390400
transform 1 0 9520 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_137
timestamp 1669390400
transform 1 0 16688 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_141
timestamp 1669390400
transform 1 0 17136 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_144
timestamp 1669390400
transform 1 0 17472 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_208
timestamp 1669390400
transform 1 0 24640 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_212
timestamp 1669390400
transform 1 0 25088 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_39_215
timestamp 1669390400
transform 1 0 25424 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_247
timestamp 1669390400
transform 1 0 29008 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_255
timestamp 1669390400
transform 1 0 29904 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_265
timestamp 1669390400
transform 1 0 31024 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_273
timestamp 1669390400
transform 1 0 31920 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_277
timestamp 1669390400
transform 1 0 32368 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_279
timestamp 1669390400
transform 1 0 32592 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_282
timestamp 1669390400
transform 1 0 32928 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_286
timestamp 1669390400
transform 1 0 33376 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_319
timestamp 1669390400
transform 1 0 37072 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_336
timestamp 1669390400
transform 1 0 38976 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_340
timestamp 1669390400
transform 1 0 39424 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_344
timestamp 1669390400
transform 1 0 39872 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_354
timestamp 1669390400
transform 1 0 40992 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_357
timestamp 1669390400
transform 1 0 41328 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_387
timestamp 1669390400
transform 1 0 44688 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_418
timestamp 1669390400
transform 1 0 48160 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_2
timestamp 1669390400
transform 1 0 1568 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_7
timestamp 1669390400
transform 1 0 2128 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_23
timestamp 1669390400
transform 1 0 3920 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_31
timestamp 1669390400
transform 1 0 4816 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_37
timestamp 1669390400
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_101
timestamp 1669390400
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_105
timestamp 1669390400
transform 1 0 13104 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_108
timestamp 1669390400
transform 1 0 13440 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_172
timestamp 1669390400
transform 1 0 20608 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_176
timestamp 1669390400
transform 1 0 21056 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_179
timestamp 1669390400
transform 1 0 21392 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_243
timestamp 1669390400
transform 1 0 28560 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_247
timestamp 1669390400
transform 1 0 29008 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_250
timestamp 1669390400
transform 1 0 29344 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_280
timestamp 1669390400
transform 1 0 32704 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_297
timestamp 1669390400
transform 1 0 34608 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_301
timestamp 1669390400
transform 1 0 35056 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_311
timestamp 1669390400
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_315
timestamp 1669390400
transform 1 0 36624 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_318
timestamp 1669390400
transform 1 0 36960 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_321
timestamp 1669390400
transform 1 0 37296 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_328
timestamp 1669390400
transform 1 0 38080 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_332
timestamp 1669390400
transform 1 0 38528 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_336
timestamp 1669390400
transform 1 0 38976 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_367
timestamp 1669390400
transform 1 0 42448 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_375
timestamp 1669390400
transform 1 0 43344 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_381
timestamp 1669390400
transform 1 0 44016 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_389
timestamp 1669390400
transform 1 0 44912 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_392
timestamp 1669390400
transform 1 0 45248 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_411
timestamp 1669390400
transform 1 0 47376 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_415
timestamp 1669390400
transform 1 0 47824 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_419
timestamp 1669390400
transform 1 0 48272 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_2
timestamp 1669390400
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_66
timestamp 1669390400
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_70
timestamp 1669390400
transform 1 0 9184 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_73
timestamp 1669390400
transform 1 0 9520 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_137
timestamp 1669390400
transform 1 0 16688 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_141
timestamp 1669390400
transform 1 0 17136 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_144
timestamp 1669390400
transform 1 0 17472 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_208
timestamp 1669390400
transform 1 0 24640 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_212
timestamp 1669390400
transform 1 0 25088 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_215
timestamp 1669390400
transform 1 0 25424 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_279
timestamp 1669390400
transform 1 0 32592 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_282
timestamp 1669390400
transform 1 0 32928 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_286
timestamp 1669390400
transform 1 0 33376 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_302
timestamp 1669390400
transform 1 0 35168 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_306
timestamp 1669390400
transform 1 0 35616 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_336
timestamp 1669390400
transform 1 0 38976 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_340
timestamp 1669390400
transform 1 0 39424 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_344
timestamp 1669390400
transform 1 0 39872 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_351
timestamp 1669390400
transform 1 0 40656 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_357
timestamp 1669390400
transform 1 0 41328 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_364
timestamp 1669390400
transform 1 0 42112 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_368
timestamp 1669390400
transform 1 0 42560 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_376
timestamp 1669390400
transform 1 0 43456 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_380
timestamp 1669390400
transform 1 0 43904 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_411
timestamp 1669390400
transform 1 0 47376 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_419
timestamp 1669390400
transform 1 0 48272 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_2
timestamp 1669390400
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_34
timestamp 1669390400
transform 1 0 5152 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_37
timestamp 1669390400
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_101
timestamp 1669390400
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_105
timestamp 1669390400
transform 1 0 13104 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_108
timestamp 1669390400
transform 1 0 13440 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_172
timestamp 1669390400
transform 1 0 20608 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_176
timestamp 1669390400
transform 1 0 21056 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_179
timestamp 1669390400
transform 1 0 21392 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_243
timestamp 1669390400
transform 1 0 28560 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_247
timestamp 1669390400
transform 1 0 29008 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_250
timestamp 1669390400
transform 1 0 29344 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_282
timestamp 1669390400
transform 1 0 32928 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_298
timestamp 1669390400
transform 1 0 34720 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_304
timestamp 1669390400
transform 1 0 35392 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_308
timestamp 1669390400
transform 1 0 35840 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_312
timestamp 1669390400
transform 1 0 36288 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_318
timestamp 1669390400
transform 1 0 36960 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_321
timestamp 1669390400
transform 1 0 37296 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_340
timestamp 1669390400
transform 1 0 39424 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_357
timestamp 1669390400
transform 1 0 41328 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_374
timestamp 1669390400
transform 1 0 43232 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_378
timestamp 1669390400
transform 1 0 43680 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_382
timestamp 1669390400
transform 1 0 44128 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_389
timestamp 1669390400
transform 1 0 44912 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_392
timestamp 1669390400
transform 1 0 45248 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_411
timestamp 1669390400
transform 1 0 47376 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_415
timestamp 1669390400
transform 1 0 47824 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_419
timestamp 1669390400
transform 1 0 48272 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_2
timestamp 1669390400
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_66
timestamp 1669390400
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_70
timestamp 1669390400
transform 1 0 9184 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_73
timestamp 1669390400
transform 1 0 9520 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_137
timestamp 1669390400
transform 1 0 16688 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_141
timestamp 1669390400
transform 1 0 17136 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_144
timestamp 1669390400
transform 1 0 17472 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_208
timestamp 1669390400
transform 1 0 24640 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_212
timestamp 1669390400
transform 1 0 25088 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_215
timestamp 1669390400
transform 1 0 25424 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_279
timestamp 1669390400
transform 1 0 32592 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_283
timestamp 1669390400
transform 1 0 33040 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_43_286
timestamp 1669390400
transform 1 0 33376 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_318
timestamp 1669390400
transform 1 0 36960 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_334
timestamp 1669390400
transform 1 0 38752 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_338
timestamp 1669390400
transform 1 0 39200 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_342
timestamp 1669390400
transform 1 0 39648 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_346
timestamp 1669390400
transform 1 0 40096 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_354
timestamp 1669390400
transform 1 0 40992 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_357
timestamp 1669390400
transform 1 0 41328 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_373
timestamp 1669390400
transform 1 0 43120 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_377
timestamp 1669390400
transform 1 0 43568 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_385
timestamp 1669390400
transform 1 0 44464 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_387
timestamp 1669390400
transform 1 0 44688 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_402
timestamp 1669390400
transform 1 0 46368 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_418
timestamp 1669390400
transform 1 0 48160 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_44_2
timestamp 1669390400
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_34
timestamp 1669390400
transform 1 0 5152 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_37
timestamp 1669390400
transform 1 0 5488 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_101
timestamp 1669390400
transform 1 0 12656 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_105
timestamp 1669390400
transform 1 0 13104 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_108
timestamp 1669390400
transform 1 0 13440 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_172
timestamp 1669390400
transform 1 0 20608 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_176
timestamp 1669390400
transform 1 0 21056 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_179
timestamp 1669390400
transform 1 0 21392 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_243
timestamp 1669390400
transform 1 0 28560 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_247
timestamp 1669390400
transform 1 0 29008 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_250
timestamp 1669390400
transform 1 0 29344 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_314
timestamp 1669390400
transform 1 0 36512 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_318
timestamp 1669390400
transform 1 0 36960 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_321
timestamp 1669390400
transform 1 0 37296 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_385
timestamp 1669390400
transform 1 0 44464 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_389
timestamp 1669390400
transform 1 0 44912 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_392
timestamp 1669390400
transform 1 0 45248 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_407
timestamp 1669390400
transform 1 0 46928 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_411
timestamp 1669390400
transform 1 0 47376 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_419
timestamp 1669390400
transform 1 0 48272 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_2
timestamp 1669390400
transform 1 0 1568 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_66
timestamp 1669390400
transform 1 0 8736 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_70
timestamp 1669390400
transform 1 0 9184 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_73
timestamp 1669390400
transform 1 0 9520 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_137
timestamp 1669390400
transform 1 0 16688 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_141
timestamp 1669390400
transform 1 0 17136 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_144
timestamp 1669390400
transform 1 0 17472 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_208
timestamp 1669390400
transform 1 0 24640 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_212
timestamp 1669390400
transform 1 0 25088 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_215
timestamp 1669390400
transform 1 0 25424 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_279
timestamp 1669390400
transform 1 0 32592 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_283
timestamp 1669390400
transform 1 0 33040 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_286
timestamp 1669390400
transform 1 0 33376 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_350
timestamp 1669390400
transform 1 0 40544 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_354
timestamp 1669390400
transform 1 0 40992 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_357
timestamp 1669390400
transform 1 0 41328 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_373
timestamp 1669390400
transform 1 0 43120 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_381
timestamp 1669390400
transform 1 0 44016 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_385
timestamp 1669390400
transform 1 0 44464 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_387
timestamp 1669390400
transform 1 0 44688 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_402
timestamp 1669390400
transform 1 0 46368 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_418
timestamp 1669390400
transform 1 0 48160 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_46_2
timestamp 1669390400
transform 1 0 1568 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_34
timestamp 1669390400
transform 1 0 5152 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_37
timestamp 1669390400
transform 1 0 5488 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_101
timestamp 1669390400
transform 1 0 12656 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_105
timestamp 1669390400
transform 1 0 13104 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_108
timestamp 1669390400
transform 1 0 13440 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_172
timestamp 1669390400
transform 1 0 20608 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_176
timestamp 1669390400
transform 1 0 21056 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_179
timestamp 1669390400
transform 1 0 21392 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_243
timestamp 1669390400
transform 1 0 28560 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_247
timestamp 1669390400
transform 1 0 29008 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_250
timestamp 1669390400
transform 1 0 29344 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_314
timestamp 1669390400
transform 1 0 36512 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_318
timestamp 1669390400
transform 1 0 36960 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_321
timestamp 1669390400
transform 1 0 37296 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_385
timestamp 1669390400
transform 1 0 44464 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_389
timestamp 1669390400
transform 1 0 44912 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_392
timestamp 1669390400
transform 1 0 45248 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_407
timestamp 1669390400
transform 1 0 46928 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_415
timestamp 1669390400
transform 1 0 47824 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_419
timestamp 1669390400
transform 1 0 48272 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_2
timestamp 1669390400
transform 1 0 1568 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_10
timestamp 1669390400
transform 1 0 2464 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_14
timestamp 1669390400
transform 1 0 2912 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_22
timestamp 1669390400
transform 1 0 3808 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_26
timestamp 1669390400
transform 1 0 4256 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_58
timestamp 1669390400
transform 1 0 7840 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_66
timestamp 1669390400
transform 1 0 8736 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_70
timestamp 1669390400
transform 1 0 9184 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_73
timestamp 1669390400
transform 1 0 9520 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_137
timestamp 1669390400
transform 1 0 16688 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_141
timestamp 1669390400
transform 1 0 17136 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_144
timestamp 1669390400
transform 1 0 17472 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_208
timestamp 1669390400
transform 1 0 24640 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_212
timestamp 1669390400
transform 1 0 25088 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_215
timestamp 1669390400
transform 1 0 25424 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_279
timestamp 1669390400
transform 1 0 32592 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_283
timestamp 1669390400
transform 1 0 33040 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_286
timestamp 1669390400
transform 1 0 33376 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_350
timestamp 1669390400
transform 1 0 40544 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_354
timestamp 1669390400
transform 1 0 40992 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_357
timestamp 1669390400
transform 1 0 41328 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_389
timestamp 1669390400
transform 1 0 44912 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_405
timestamp 1669390400
transform 1 0 46704 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_413
timestamp 1669390400
transform 1 0 47600 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_417
timestamp 1669390400
transform 1 0 48048 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_419
timestamp 1669390400
transform 1 0 48272 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_2
timestamp 1669390400
transform 1 0 1568 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_17
timestamp 1669390400
transform 1 0 3248 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_33
timestamp 1669390400
transform 1 0 5040 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_37
timestamp 1669390400
transform 1 0 5488 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_101
timestamp 1669390400
transform 1 0 12656 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_105
timestamp 1669390400
transform 1 0 13104 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_108
timestamp 1669390400
transform 1 0 13440 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_172
timestamp 1669390400
transform 1 0 20608 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_176
timestamp 1669390400
transform 1 0 21056 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_179
timestamp 1669390400
transform 1 0 21392 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_243
timestamp 1669390400
transform 1 0 28560 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_247
timestamp 1669390400
transform 1 0 29008 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_250
timestamp 1669390400
transform 1 0 29344 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_314
timestamp 1669390400
transform 1 0 36512 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_318
timestamp 1669390400
transform 1 0 36960 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_321
timestamp 1669390400
transform 1 0 37296 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_385
timestamp 1669390400
transform 1 0 44464 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_389
timestamp 1669390400
transform 1 0 44912 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_392
timestamp 1669390400
transform 1 0 45248 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_407
timestamp 1669390400
transform 1 0 46928 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_415
timestamp 1669390400
transform 1 0 47824 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_419
timestamp 1669390400
transform 1 0 48272 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_2
timestamp 1669390400
transform 1 0 1568 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_66
timestamp 1669390400
transform 1 0 8736 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_70
timestamp 1669390400
transform 1 0 9184 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_73
timestamp 1669390400
transform 1 0 9520 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_137
timestamp 1669390400
transform 1 0 16688 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_141
timestamp 1669390400
transform 1 0 17136 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_144
timestamp 1669390400
transform 1 0 17472 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_208
timestamp 1669390400
transform 1 0 24640 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_212
timestamp 1669390400
transform 1 0 25088 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_215
timestamp 1669390400
transform 1 0 25424 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_279
timestamp 1669390400
transform 1 0 32592 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_283
timestamp 1669390400
transform 1 0 33040 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_286
timestamp 1669390400
transform 1 0 33376 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_350
timestamp 1669390400
transform 1 0 40544 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_354
timestamp 1669390400
transform 1 0 40992 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_49_357
timestamp 1669390400
transform 1 0 41328 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_389
timestamp 1669390400
transform 1 0 44912 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_405
timestamp 1669390400
transform 1 0 46704 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_413
timestamp 1669390400
transform 1 0 47600 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_417
timestamp 1669390400
transform 1 0 48048 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_419
timestamp 1669390400
transform 1 0 48272 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_2
timestamp 1669390400
transform 1 0 1568 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_34
timestamp 1669390400
transform 1 0 5152 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_37
timestamp 1669390400
transform 1 0 5488 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_101
timestamp 1669390400
transform 1 0 12656 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_105
timestamp 1669390400
transform 1 0 13104 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_108
timestamp 1669390400
transform 1 0 13440 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_172
timestamp 1669390400
transform 1 0 20608 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_176
timestamp 1669390400
transform 1 0 21056 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_179
timestamp 1669390400
transform 1 0 21392 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_243
timestamp 1669390400
transform 1 0 28560 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_247
timestamp 1669390400
transform 1 0 29008 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_250
timestamp 1669390400
transform 1 0 29344 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_314
timestamp 1669390400
transform 1 0 36512 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_318
timestamp 1669390400
transform 1 0 36960 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_321
timestamp 1669390400
transform 1 0 37296 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_385
timestamp 1669390400
transform 1 0 44464 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_389
timestamp 1669390400
transform 1 0 44912 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_392
timestamp 1669390400
transform 1 0 45248 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_407
timestamp 1669390400
transform 1 0 46928 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_415
timestamp 1669390400
transform 1 0 47824 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_419
timestamp 1669390400
transform 1 0 48272 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_2
timestamp 1669390400
transform 1 0 1568 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_66
timestamp 1669390400
transform 1 0 8736 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_70
timestamp 1669390400
transform 1 0 9184 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_73
timestamp 1669390400
transform 1 0 9520 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_137
timestamp 1669390400
transform 1 0 16688 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_141
timestamp 1669390400
transform 1 0 17136 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_144
timestamp 1669390400
transform 1 0 17472 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_208
timestamp 1669390400
transform 1 0 24640 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_212
timestamp 1669390400
transform 1 0 25088 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_215
timestamp 1669390400
transform 1 0 25424 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_279
timestamp 1669390400
transform 1 0 32592 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_283
timestamp 1669390400
transform 1 0 33040 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_286
timestamp 1669390400
transform 1 0 33376 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_350
timestamp 1669390400
transform 1 0 40544 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_354
timestamp 1669390400
transform 1 0 40992 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_51_357
timestamp 1669390400
transform 1 0 41328 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_389
timestamp 1669390400
transform 1 0 44912 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_405
timestamp 1669390400
transform 1 0 46704 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_413
timestamp 1669390400
transform 1 0 47600 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_417
timestamp 1669390400
transform 1 0 48048 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_419
timestamp 1669390400
transform 1 0 48272 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_52_2
timestamp 1669390400
transform 1 0 1568 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_34
timestamp 1669390400
transform 1 0 5152 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_37
timestamp 1669390400
transform 1 0 5488 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_101
timestamp 1669390400
transform 1 0 12656 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_105
timestamp 1669390400
transform 1 0 13104 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_108
timestamp 1669390400
transform 1 0 13440 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_172
timestamp 1669390400
transform 1 0 20608 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_176
timestamp 1669390400
transform 1 0 21056 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_179
timestamp 1669390400
transform 1 0 21392 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_243
timestamp 1669390400
transform 1 0 28560 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_247
timestamp 1669390400
transform 1 0 29008 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_250
timestamp 1669390400
transform 1 0 29344 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_314
timestamp 1669390400
transform 1 0 36512 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_318
timestamp 1669390400
transform 1 0 36960 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_321
timestamp 1669390400
transform 1 0 37296 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_385
timestamp 1669390400
transform 1 0 44464 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_389
timestamp 1669390400
transform 1 0 44912 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_392
timestamp 1669390400
transform 1 0 45248 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_407
timestamp 1669390400
transform 1 0 46928 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_415
timestamp 1669390400
transform 1 0 47824 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_419
timestamp 1669390400
transform 1 0 48272 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_2
timestamp 1669390400
transform 1 0 1568 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_66
timestamp 1669390400
transform 1 0 8736 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_70
timestamp 1669390400
transform 1 0 9184 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_73
timestamp 1669390400
transform 1 0 9520 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_137
timestamp 1669390400
transform 1 0 16688 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_141
timestamp 1669390400
transform 1 0 17136 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_144
timestamp 1669390400
transform 1 0 17472 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_208
timestamp 1669390400
transform 1 0 24640 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_212
timestamp 1669390400
transform 1 0 25088 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_215
timestamp 1669390400
transform 1 0 25424 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_279
timestamp 1669390400
transform 1 0 32592 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_283
timestamp 1669390400
transform 1 0 33040 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_286
timestamp 1669390400
transform 1 0 33376 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_350
timestamp 1669390400
transform 1 0 40544 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_354
timestamp 1669390400
transform 1 0 40992 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_357
timestamp 1669390400
transform 1 0 41328 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_373
timestamp 1669390400
transform 1 0 43120 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_381
timestamp 1669390400
transform 1 0 44016 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_383
timestamp 1669390400
transform 1 0 44240 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_386
timestamp 1669390400
transform 1 0 44576 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_402
timestamp 1669390400
transform 1 0 46368 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_406
timestamp 1669390400
transform 1 0 46816 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_414
timestamp 1669390400
transform 1 0 47712 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_418
timestamp 1669390400
transform 1 0 48160 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_2
timestamp 1669390400
transform 1 0 1568 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_7
timestamp 1669390400
transform 1 0 2128 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_23
timestamp 1669390400
transform 1 0 3920 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_31
timestamp 1669390400
transform 1 0 4816 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_37
timestamp 1669390400
transform 1 0 5488 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_69
timestamp 1669390400
transform 1 0 9072 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_72
timestamp 1669390400
transform 1 0 9408 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_104
timestamp 1669390400
transform 1 0 12992 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_107
timestamp 1669390400
transform 1 0 13328 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_139
timestamp 1669390400
transform 1 0 16912 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_142
timestamp 1669390400
transform 1 0 17248 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_174
timestamp 1669390400
transform 1 0 20832 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_177
timestamp 1669390400
transform 1 0 21168 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_209
timestamp 1669390400
transform 1 0 24752 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_212
timestamp 1669390400
transform 1 0 25088 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_244
timestamp 1669390400
transform 1 0 28672 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_247
timestamp 1669390400
transform 1 0 29008 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_279
timestamp 1669390400
transform 1 0 32592 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_282
timestamp 1669390400
transform 1 0 32928 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_314
timestamp 1669390400
transform 1 0 36512 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_317
timestamp 1669390400
transform 1 0 36848 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_349
timestamp 1669390400
transform 1 0 40432 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_352
timestamp 1669390400
transform 1 0 40768 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_368
timestamp 1669390400
transform 1 0 42560 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_376
timestamp 1669390400
transform 1 0 43456 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_380
timestamp 1669390400
transform 1 0 43904 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_384
timestamp 1669390400
transform 1 0 44352 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_387
timestamp 1669390400
transform 1 0 44688 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_402
timestamp 1669390400
transform 1 0 46368 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_418
timestamp 1669390400
transform 1 0 48160 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1669390400
transform -1 0 48608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1669390400
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1669390400
transform -1 0 48608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1669390400
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1669390400
transform -1 0 48608 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1669390400
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1669390400
transform -1 0 48608 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1669390400
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1669390400
transform -1 0 48608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1669390400
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1669390400
transform -1 0 48608 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1669390400
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1669390400
transform -1 0 48608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1669390400
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1669390400
transform -1 0 48608 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1669390400
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1669390400
transform -1 0 48608 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1669390400
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1669390400
transform -1 0 48608 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1669390400
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1669390400
transform -1 0 48608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1669390400
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1669390400
transform -1 0 48608 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1669390400
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1669390400
transform -1 0 48608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1669390400
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1669390400
transform -1 0 48608 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1669390400
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1669390400
transform -1 0 48608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1669390400
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1669390400
transform -1 0 48608 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1669390400
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1669390400
transform -1 0 48608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_34
timestamp 1669390400
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_35
timestamp 1669390400
transform -1 0 48608 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_36
timestamp 1669390400
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_37
timestamp 1669390400
transform -1 0 48608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_38
timestamp 1669390400
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_39
timestamp 1669390400
transform -1 0 48608 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_40
timestamp 1669390400
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_41
timestamp 1669390400
transform -1 0 48608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_42
timestamp 1669390400
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_43
timestamp 1669390400
transform -1 0 48608 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_44
timestamp 1669390400
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_45
timestamp 1669390400
transform -1 0 48608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_46
timestamp 1669390400
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_47
timestamp 1669390400
transform -1 0 48608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_48
timestamp 1669390400
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_49
timestamp 1669390400
transform -1 0 48608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_50
timestamp 1669390400
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_51
timestamp 1669390400
transform -1 0 48608 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_52
timestamp 1669390400
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_53
timestamp 1669390400
transform -1 0 48608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_54
timestamp 1669390400
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_55
timestamp 1669390400
transform -1 0 48608 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_56
timestamp 1669390400
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_57
timestamp 1669390400
transform -1 0 48608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_58
timestamp 1669390400
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_59
timestamp 1669390400
transform -1 0 48608 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_60
timestamp 1669390400
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_61
timestamp 1669390400
transform -1 0 48608 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_62
timestamp 1669390400
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_63
timestamp 1669390400
transform -1 0 48608 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_64
timestamp 1669390400
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_65
timestamp 1669390400
transform -1 0 48608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_66
timestamp 1669390400
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_67
timestamp 1669390400
transform -1 0 48608 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_68
timestamp 1669390400
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_69
timestamp 1669390400
transform -1 0 48608 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_70
timestamp 1669390400
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_71
timestamp 1669390400
transform -1 0 48608 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_72
timestamp 1669390400
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_73
timestamp 1669390400
transform -1 0 48608 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_74
timestamp 1669390400
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_75
timestamp 1669390400
transform -1 0 48608 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_76
timestamp 1669390400
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_77
timestamp 1669390400
transform -1 0 48608 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_78
timestamp 1669390400
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_79
timestamp 1669390400
transform -1 0 48608 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_80
timestamp 1669390400
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_81
timestamp 1669390400
transform -1 0 48608 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_82
timestamp 1669390400
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_83
timestamp 1669390400
transform -1 0 48608 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_84
timestamp 1669390400
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_85
timestamp 1669390400
transform -1 0 48608 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_86
timestamp 1669390400
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_87
timestamp 1669390400
transform -1 0 48608 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_88
timestamp 1669390400
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_89
timestamp 1669390400
transform -1 0 48608 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_90
timestamp 1669390400
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_91
timestamp 1669390400
transform -1 0 48608 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_92
timestamp 1669390400
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_93
timestamp 1669390400
transform -1 0 48608 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_94
timestamp 1669390400
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_95
timestamp 1669390400
transform -1 0 48608 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_96
timestamp 1669390400
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_97
timestamp 1669390400
transform -1 0 48608 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_98
timestamp 1669390400
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_99
timestamp 1669390400
transform -1 0 48608 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_100
timestamp 1669390400
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_101
timestamp 1669390400
transform -1 0 48608 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_102
timestamp 1669390400
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_103
timestamp 1669390400
transform -1 0 48608 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_104
timestamp 1669390400
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_105
timestamp 1669390400
transform -1 0 48608 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_106
timestamp 1669390400
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_107
timestamp 1669390400
transform -1 0 48608 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_108
timestamp 1669390400
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_109
timestamp 1669390400
transform -1 0 48608 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_110 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_111
timestamp 1669390400
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_112
timestamp 1669390400
transform 1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_113
timestamp 1669390400
transform 1 0 17024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_114
timestamp 1669390400
transform 1 0 20944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_115
timestamp 1669390400
transform 1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_116
timestamp 1669390400
transform 1 0 28784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_117
timestamp 1669390400
transform 1 0 32704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_118
timestamp 1669390400
transform 1 0 36624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_119
timestamp 1669390400
transform 1 0 40544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_120
timestamp 1669390400
transform 1 0 44464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_121
timestamp 1669390400
transform 1 0 9296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_122
timestamp 1669390400
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_123
timestamp 1669390400
transform 1 0 25200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_124
timestamp 1669390400
transform 1 0 33152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_125
timestamp 1669390400
transform 1 0 41104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_126
timestamp 1669390400
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_127
timestamp 1669390400
transform 1 0 13216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_128
timestamp 1669390400
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_129
timestamp 1669390400
transform 1 0 29120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_130
timestamp 1669390400
transform 1 0 37072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_131
timestamp 1669390400
transform 1 0 45024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_132
timestamp 1669390400
transform 1 0 9296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_133
timestamp 1669390400
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_134
timestamp 1669390400
transform 1 0 25200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_135
timestamp 1669390400
transform 1 0 33152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_136
timestamp 1669390400
transform 1 0 41104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_137
timestamp 1669390400
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_138
timestamp 1669390400
transform 1 0 13216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_139
timestamp 1669390400
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_140
timestamp 1669390400
transform 1 0 29120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_141
timestamp 1669390400
transform 1 0 37072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_142
timestamp 1669390400
transform 1 0 45024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_143
timestamp 1669390400
transform 1 0 9296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_144
timestamp 1669390400
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_145
timestamp 1669390400
transform 1 0 25200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_146
timestamp 1669390400
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_147
timestamp 1669390400
transform 1 0 41104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_148
timestamp 1669390400
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_149
timestamp 1669390400
transform 1 0 13216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_150
timestamp 1669390400
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_151
timestamp 1669390400
transform 1 0 29120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_152
timestamp 1669390400
transform 1 0 37072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_153
timestamp 1669390400
transform 1 0 45024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_154
timestamp 1669390400
transform 1 0 9296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_155
timestamp 1669390400
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_156
timestamp 1669390400
transform 1 0 25200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_157
timestamp 1669390400
transform 1 0 33152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_158
timestamp 1669390400
transform 1 0 41104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_159
timestamp 1669390400
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_160
timestamp 1669390400
transform 1 0 13216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_161
timestamp 1669390400
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_162
timestamp 1669390400
transform 1 0 29120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_163
timestamp 1669390400
transform 1 0 37072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_164
timestamp 1669390400
transform 1 0 45024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_165
timestamp 1669390400
transform 1 0 9296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_166
timestamp 1669390400
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_167
timestamp 1669390400
transform 1 0 25200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_168
timestamp 1669390400
transform 1 0 33152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_169
timestamp 1669390400
transform 1 0 41104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_170
timestamp 1669390400
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_171
timestamp 1669390400
transform 1 0 13216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_172
timestamp 1669390400
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_173
timestamp 1669390400
transform 1 0 29120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_174
timestamp 1669390400
transform 1 0 37072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_175
timestamp 1669390400
transform 1 0 45024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_176
timestamp 1669390400
transform 1 0 9296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_177
timestamp 1669390400
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_178
timestamp 1669390400
transform 1 0 25200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_179
timestamp 1669390400
transform 1 0 33152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_180
timestamp 1669390400
transform 1 0 41104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_181
timestamp 1669390400
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_182
timestamp 1669390400
transform 1 0 13216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_183
timestamp 1669390400
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_184
timestamp 1669390400
transform 1 0 29120 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_185
timestamp 1669390400
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_186
timestamp 1669390400
transform 1 0 45024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_187
timestamp 1669390400
transform 1 0 9296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_188
timestamp 1669390400
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_189
timestamp 1669390400
transform 1 0 25200 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_190
timestamp 1669390400
transform 1 0 33152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_191
timestamp 1669390400
transform 1 0 41104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_192
timestamp 1669390400
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_193
timestamp 1669390400
transform 1 0 13216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_194
timestamp 1669390400
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_195
timestamp 1669390400
transform 1 0 29120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_196
timestamp 1669390400
transform 1 0 37072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_197
timestamp 1669390400
transform 1 0 45024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_198
timestamp 1669390400
transform 1 0 9296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_199
timestamp 1669390400
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_200
timestamp 1669390400
transform 1 0 25200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_201
timestamp 1669390400
transform 1 0 33152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_202
timestamp 1669390400
transform 1 0 41104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_203
timestamp 1669390400
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_204
timestamp 1669390400
transform 1 0 13216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_205
timestamp 1669390400
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_206
timestamp 1669390400
transform 1 0 29120 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_207
timestamp 1669390400
transform 1 0 37072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_208
timestamp 1669390400
transform 1 0 45024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_209
timestamp 1669390400
transform 1 0 9296 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_210
timestamp 1669390400
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_211
timestamp 1669390400
transform 1 0 25200 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_212
timestamp 1669390400
transform 1 0 33152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_213
timestamp 1669390400
transform 1 0 41104 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_214
timestamp 1669390400
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_215
timestamp 1669390400
transform 1 0 13216 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_216
timestamp 1669390400
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_217
timestamp 1669390400
transform 1 0 29120 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_218
timestamp 1669390400
transform 1 0 37072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_219
timestamp 1669390400
transform 1 0 45024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_220
timestamp 1669390400
transform 1 0 9296 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_221
timestamp 1669390400
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_222
timestamp 1669390400
transform 1 0 25200 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_223
timestamp 1669390400
transform 1 0 33152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_224
timestamp 1669390400
transform 1 0 41104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_225
timestamp 1669390400
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_226
timestamp 1669390400
transform 1 0 13216 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_227
timestamp 1669390400
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_228
timestamp 1669390400
transform 1 0 29120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_229
timestamp 1669390400
transform 1 0 37072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_230
timestamp 1669390400
transform 1 0 45024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_231
timestamp 1669390400
transform 1 0 9296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_232
timestamp 1669390400
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_233
timestamp 1669390400
transform 1 0 25200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_234
timestamp 1669390400
transform 1 0 33152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_235
timestamp 1669390400
transform 1 0 41104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_236
timestamp 1669390400
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_237
timestamp 1669390400
transform 1 0 13216 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_238
timestamp 1669390400
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_239
timestamp 1669390400
transform 1 0 29120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_240
timestamp 1669390400
transform 1 0 37072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_241
timestamp 1669390400
transform 1 0 45024 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_242
timestamp 1669390400
transform 1 0 9296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_243
timestamp 1669390400
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_244
timestamp 1669390400
transform 1 0 25200 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_245
timestamp 1669390400
transform 1 0 33152 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_246
timestamp 1669390400
transform 1 0 41104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_247
timestamp 1669390400
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_248
timestamp 1669390400
transform 1 0 13216 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_249
timestamp 1669390400
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_250
timestamp 1669390400
transform 1 0 29120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_251
timestamp 1669390400
transform 1 0 37072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_252
timestamp 1669390400
transform 1 0 45024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_253
timestamp 1669390400
transform 1 0 9296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_254
timestamp 1669390400
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_255
timestamp 1669390400
transform 1 0 25200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_256
timestamp 1669390400
transform 1 0 33152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_257
timestamp 1669390400
transform 1 0 41104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_258
timestamp 1669390400
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_259
timestamp 1669390400
transform 1 0 13216 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_260
timestamp 1669390400
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_261
timestamp 1669390400
transform 1 0 29120 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_262
timestamp 1669390400
transform 1 0 37072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_263
timestamp 1669390400
transform 1 0 45024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_264
timestamp 1669390400
transform 1 0 9296 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_265
timestamp 1669390400
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_266
timestamp 1669390400
transform 1 0 25200 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_267
timestamp 1669390400
transform 1 0 33152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_268
timestamp 1669390400
transform 1 0 41104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_269
timestamp 1669390400
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_270
timestamp 1669390400
transform 1 0 13216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_271
timestamp 1669390400
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_272
timestamp 1669390400
transform 1 0 29120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_273
timestamp 1669390400
transform 1 0 37072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_274
timestamp 1669390400
transform 1 0 45024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_275
timestamp 1669390400
transform 1 0 9296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_276
timestamp 1669390400
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_277
timestamp 1669390400
transform 1 0 25200 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_278
timestamp 1669390400
transform 1 0 33152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_279
timestamp 1669390400
transform 1 0 41104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_280
timestamp 1669390400
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_281
timestamp 1669390400
transform 1 0 13216 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_282
timestamp 1669390400
transform 1 0 21168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_283
timestamp 1669390400
transform 1 0 29120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_284
timestamp 1669390400
transform 1 0 37072 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_285
timestamp 1669390400
transform 1 0 45024 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_286
timestamp 1669390400
transform 1 0 9296 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_287
timestamp 1669390400
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_288
timestamp 1669390400
transform 1 0 25200 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_289
timestamp 1669390400
transform 1 0 33152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_290
timestamp 1669390400
transform 1 0 41104 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_291
timestamp 1669390400
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_292
timestamp 1669390400
transform 1 0 13216 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_293
timestamp 1669390400
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_294
timestamp 1669390400
transform 1 0 29120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_295
timestamp 1669390400
transform 1 0 37072 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_296
timestamp 1669390400
transform 1 0 45024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_297
timestamp 1669390400
transform 1 0 9296 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_298
timestamp 1669390400
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_299
timestamp 1669390400
transform 1 0 25200 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_300
timestamp 1669390400
transform 1 0 33152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_301
timestamp 1669390400
transform 1 0 41104 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_302
timestamp 1669390400
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_303
timestamp 1669390400
transform 1 0 13216 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_304
timestamp 1669390400
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_305
timestamp 1669390400
transform 1 0 29120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_306
timestamp 1669390400
transform 1 0 37072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_307
timestamp 1669390400
transform 1 0 45024 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_308
timestamp 1669390400
transform 1 0 9296 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_309
timestamp 1669390400
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_310
timestamp 1669390400
transform 1 0 25200 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_311
timestamp 1669390400
transform 1 0 33152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_312
timestamp 1669390400
transform 1 0 41104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_313
timestamp 1669390400
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_314
timestamp 1669390400
transform 1 0 13216 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_315
timestamp 1669390400
transform 1 0 21168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_316
timestamp 1669390400
transform 1 0 29120 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_317
timestamp 1669390400
transform 1 0 37072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_318
timestamp 1669390400
transform 1 0 45024 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_319
timestamp 1669390400
transform 1 0 9296 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_320
timestamp 1669390400
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_321
timestamp 1669390400
transform 1 0 25200 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_322
timestamp 1669390400
transform 1 0 33152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_323
timestamp 1669390400
transform 1 0 41104 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_324
timestamp 1669390400
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_325
timestamp 1669390400
transform 1 0 13216 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_326
timestamp 1669390400
transform 1 0 21168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_327
timestamp 1669390400
transform 1 0 29120 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_328
timestamp 1669390400
transform 1 0 37072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_329
timestamp 1669390400
transform 1 0 45024 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_330
timestamp 1669390400
transform 1 0 9296 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_331
timestamp 1669390400
transform 1 0 17248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_332
timestamp 1669390400
transform 1 0 25200 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_333
timestamp 1669390400
transform 1 0 33152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_334
timestamp 1669390400
transform 1 0 41104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_335
timestamp 1669390400
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_336
timestamp 1669390400
transform 1 0 13216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_337
timestamp 1669390400
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_338
timestamp 1669390400
transform 1 0 29120 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_339
timestamp 1669390400
transform 1 0 37072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_340
timestamp 1669390400
transform 1 0 45024 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_341
timestamp 1669390400
transform 1 0 9296 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_342
timestamp 1669390400
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_343
timestamp 1669390400
transform 1 0 25200 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_344
timestamp 1669390400
transform 1 0 33152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_345
timestamp 1669390400
transform 1 0 41104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_346
timestamp 1669390400
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_347
timestamp 1669390400
transform 1 0 13216 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_348
timestamp 1669390400
transform 1 0 21168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_349
timestamp 1669390400
transform 1 0 29120 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_350
timestamp 1669390400
transform 1 0 37072 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_351
timestamp 1669390400
transform 1 0 45024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_352
timestamp 1669390400
transform 1 0 9296 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_353
timestamp 1669390400
transform 1 0 17248 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_354
timestamp 1669390400
transform 1 0 25200 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_355
timestamp 1669390400
transform 1 0 33152 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_356
timestamp 1669390400
transform 1 0 41104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_357
timestamp 1669390400
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_358
timestamp 1669390400
transform 1 0 13216 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_359
timestamp 1669390400
transform 1 0 21168 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_360
timestamp 1669390400
transform 1 0 29120 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_361
timestamp 1669390400
transform 1 0 37072 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_362
timestamp 1669390400
transform 1 0 45024 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_363
timestamp 1669390400
transform 1 0 9296 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_364
timestamp 1669390400
transform 1 0 17248 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_365
timestamp 1669390400
transform 1 0 25200 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_366
timestamp 1669390400
transform 1 0 33152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_367
timestamp 1669390400
transform 1 0 41104 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_368
timestamp 1669390400
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_369
timestamp 1669390400
transform 1 0 13216 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_370
timestamp 1669390400
transform 1 0 21168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_371
timestamp 1669390400
transform 1 0 29120 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_372
timestamp 1669390400
transform 1 0 37072 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_373
timestamp 1669390400
transform 1 0 45024 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_374
timestamp 1669390400
transform 1 0 9296 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_375
timestamp 1669390400
transform 1 0 17248 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_376
timestamp 1669390400
transform 1 0 25200 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_377
timestamp 1669390400
transform 1 0 33152 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_378
timestamp 1669390400
transform 1 0 41104 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_379
timestamp 1669390400
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_380
timestamp 1669390400
transform 1 0 13216 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_381
timestamp 1669390400
transform 1 0 21168 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_382
timestamp 1669390400
transform 1 0 29120 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_383
timestamp 1669390400
transform 1 0 37072 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_384
timestamp 1669390400
transform 1 0 45024 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_385
timestamp 1669390400
transform 1 0 9296 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_386
timestamp 1669390400
transform 1 0 17248 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_387
timestamp 1669390400
transform 1 0 25200 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_388
timestamp 1669390400
transform 1 0 33152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_389
timestamp 1669390400
transform 1 0 41104 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_390
timestamp 1669390400
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_391
timestamp 1669390400
transform 1 0 13216 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_392
timestamp 1669390400
transform 1 0 21168 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_393
timestamp 1669390400
transform 1 0 29120 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_394
timestamp 1669390400
transform 1 0 37072 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_395
timestamp 1669390400
transform 1 0 45024 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_396
timestamp 1669390400
transform 1 0 9296 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_397
timestamp 1669390400
transform 1 0 17248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_398
timestamp 1669390400
transform 1 0 25200 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_399
timestamp 1669390400
transform 1 0 33152 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_400
timestamp 1669390400
transform 1 0 41104 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_401
timestamp 1669390400
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_402
timestamp 1669390400
transform 1 0 13216 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_403
timestamp 1669390400
transform 1 0 21168 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_404
timestamp 1669390400
transform 1 0 29120 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_405
timestamp 1669390400
transform 1 0 37072 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_406
timestamp 1669390400
transform 1 0 45024 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_407
timestamp 1669390400
transform 1 0 9296 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_408
timestamp 1669390400
transform 1 0 17248 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_409
timestamp 1669390400
transform 1 0 25200 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_410
timestamp 1669390400
transform 1 0 33152 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_411
timestamp 1669390400
transform 1 0 41104 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_412
timestamp 1669390400
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_413
timestamp 1669390400
transform 1 0 9184 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_414
timestamp 1669390400
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_415
timestamp 1669390400
transform 1 0 17024 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_416
timestamp 1669390400
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_417
timestamp 1669390400
transform 1 0 24864 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_418
timestamp 1669390400
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_419
timestamp 1669390400
transform 1 0 32704 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_420
timestamp 1669390400
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_421
timestamp 1669390400
transform 1 0 40544 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_422
timestamp 1669390400
transform 1 0 44464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _078_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 25648 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _079_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 22400 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _080_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 20384 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _081_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 21392 0 -1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _082_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 38304 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _083_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 39312 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _084_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 35280 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _085_
timestamp 1669390400
transform -1 0 35616 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _086_
timestamp 1669390400
transform -1 0 38192 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _087_
timestamp 1669390400
transform -1 0 38080 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _088_
timestamp 1669390400
transform 1 0 38304 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _089_
timestamp 1669390400
transform -1 0 38528 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _090_
timestamp 1669390400
transform 1 0 39200 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _091_
timestamp 1669390400
transform -1 0 39648 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _092_
timestamp 1669390400
transform 1 0 44016 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _093_
timestamp 1669390400
transform -1 0 47376 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _094_
timestamp 1669390400
transform -1 0 48272 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _095_
timestamp 1669390400
transform -1 0 47376 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _096_
timestamp 1669390400
transform -1 0 47264 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _097_
timestamp 1669390400
transform 1 0 46256 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _098_
timestamp 1669390400
transform -1 0 44016 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _099_
timestamp 1669390400
transform 1 0 45360 0 1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _100_
timestamp 1669390400
transform -1 0 44912 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _101_
timestamp 1669390400
transform 1 0 42224 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _102_
timestamp 1669390400
transform 1 0 45360 0 1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _103_
timestamp 1669390400
transform -1 0 44016 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _104_
timestamp 1669390400
transform 1 0 44128 0 -1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _105_
timestamp 1669390400
transform -1 0 43008 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _106_
timestamp 1669390400
transform -1 0 47040 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _107_
timestamp 1669390400
transform -1 0 48160 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _108_
timestamp 1669390400
transform 1 0 45360 0 1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _109_
timestamp 1669390400
transform -1 0 44912 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _110_
timestamp 1669390400
transform 1 0 43680 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _111_
timestamp 1669390400
transform 1 0 45584 0 1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _112_
timestamp 1669390400
transform 1 0 44240 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _113_
timestamp 1669390400
transform -1 0 47376 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _114_
timestamp 1669390400
transform -1 0 48272 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _115_
timestamp 1669390400
transform 1 0 45696 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _116_
timestamp 1669390400
transform 1 0 44240 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _117_
timestamp 1669390400
transform 1 0 43232 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _118_
timestamp 1669390400
transform -1 0 43120 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _119_
timestamp 1669390400
transform 1 0 39984 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _120_
timestamp 1669390400
transform 1 0 41440 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _121_
timestamp 1669390400
transform 1 0 40880 0 1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _122_
timestamp 1669390400
transform -1 0 38976 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _123_
timestamp 1669390400
transform 1 0 39200 0 -1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _124_
timestamp 1669390400
transform -1 0 38640 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _125_
timestamp 1669390400
transform -1 0 47040 0 1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _126_
timestamp 1669390400
transform -1 0 46816 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _127_
timestamp 1669390400
transform 1 0 45360 0 1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _128_
timestamp 1669390400
transform 1 0 42448 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _129_
timestamp 1669390400
transform 1 0 42896 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _130_
timestamp 1669390400
transform 1 0 45584 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _131_
timestamp 1669390400
transform 1 0 44240 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _132_
timestamp 1669390400
transform 1 0 45696 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _133_
timestamp 1669390400
transform 1 0 44240 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _134_
timestamp 1669390400
transform 1 0 45696 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _135_
timestamp 1669390400
transform 1 0 44240 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _136_
timestamp 1669390400
transform -1 0 47376 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _137_
timestamp 1669390400
transform -1 0 48272 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _138_
timestamp 1669390400
transform -1 0 40992 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _139_
timestamp 1669390400
transform 1 0 41552 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _140_
timestamp 1669390400
transform 1 0 41440 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _141_
timestamp 1669390400
transform 1 0 41440 0 -1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _142_
timestamp 1669390400
transform -1 0 40656 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _143_
timestamp 1669390400
transform 1 0 39648 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _144_
timestamp 1669390400
transform -1 0 38080 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _145_
timestamp 1669390400
transform 1 0 37744 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _146_
timestamp 1669390400
transform -1 0 36176 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _147_
timestamp 1669390400
transform -1 0 39872 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _148_
timestamp 1669390400
transform 1 0 37296 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _149_
timestamp 1669390400
transform 1 0 37408 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _150_
timestamp 1669390400
transform 1 0 35280 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _151_
timestamp 1669390400
transform 1 0 35840 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _152_
timestamp 1669390400
transform 1 0 33488 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _153_
timestamp 1669390400
transform -1 0 32816 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _154_
timestamp 1669390400
transform 1 0 32928 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _155_
timestamp 1669390400
transform -1 0 31024 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _156_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5936 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _157_
timestamp 1669390400
transform 1 0 13216 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _158_
timestamp 1669390400
transform 1 0 22176 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _159_
timestamp 1669390400
transform 1 0 5488 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _160_
timestamp 1669390400
transform 1 0 10864 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _161_
timestamp 1669390400
transform 1 0 16912 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _162_
timestamp 1669390400
transform 1 0 5600 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _163_
timestamp 1669390400
transform 1 0 13552 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _164_
timestamp 1669390400
transform 1 0 19264 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _165_
timestamp 1669390400
transform 1 0 33712 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _166_
timestamp 1669390400
transform 1 0 35280 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _167_
timestamp 1669390400
transform 1 0 37072 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _168_
timestamp 1669390400
transform 1 0 38080 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _169_
timestamp 1669390400
transform -1 0 47824 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _170_
timestamp 1669390400
transform 1 0 44240 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _171_
timestamp 1669390400
transform 1 0 42784 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _172_
timestamp 1669390400
transform 1 0 43680 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _173_
timestamp 1669390400
transform 1 0 41664 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _174_
timestamp 1669390400
transform 1 0 40992 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _175_
timestamp 1669390400
transform -1 0 47264 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _176_
timestamp 1669390400
transform 1 0 43568 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _177_
timestamp 1669390400
transform 1 0 43792 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _178_
timestamp 1669390400
transform 1 0 44464 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _179_
timestamp 1669390400
transform 1 0 44352 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _180_
timestamp 1669390400
transform 1 0 41440 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _181_
timestamp 1669390400
transform 1 0 37408 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _182_
timestamp 1669390400
transform 1 0 36624 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _183_
timestamp 1669390400
transform 1 0 43680 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _184_
timestamp 1669390400
transform 1 0 42672 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _185_
timestamp 1669390400
transform 1 0 43792 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _186_
timestamp 1669390400
transform 1 0 44912 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _187_
timestamp 1669390400
transform 1 0 44128 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _188_
timestamp 1669390400
transform 1 0 44464 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _189_
timestamp 1669390400
transform 1 0 41440 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _190_
timestamp 1669390400
transform 1 0 39200 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _191_
timestamp 1669390400
transform 1 0 35728 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _192_
timestamp 1669390400
transform 1 0 33824 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _193_
timestamp 1669390400
transform 1 0 37408 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _194_
timestamp 1669390400
transform 1 0 35280 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _195_
timestamp 1669390400
transform 1 0 31136 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _196_
timestamp 1669390400
transform 1 0 29456 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _205_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 47824 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _206_
timestamp 1669390400
transform -1 0 3808 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clock dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 26656 0 -1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_0__f_clock
timestamp 1669390400
transform 1 0 34160 0 -1 12544
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_1__f_clock
timestamp 1669390400
transform -1 0 24640 0 -1 12544
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_2__f_clock
timestamp 1669390400
transform 1 0 34160 0 -1 23520
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_3__f_clock
timestamp 1669390400
transform 1 0 30352 0 1 26656
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input1 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1680 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input2
timestamp 1669390400
transform 1 0 1680 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input3
timestamp 1669390400
transform 1 0 1680 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output4
timestamp 1669390400
transform 1 0 44464 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output5 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 44800 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output6
timestamp 1669390400
transform 1 0 43344 0 1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output7
timestamp 1669390400
transform 1 0 45360 0 1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output8
timestamp 1669390400
transform -1 0 46368 0 -1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output9
timestamp 1669390400
transform -1 0 44912 0 1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output10
timestamp 1669390400
transform -1 0 44240 0 -1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output11
timestamp 1669390400
transform 1 0 45360 0 1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output12
timestamp 1669390400
transform 1 0 44912 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output13
timestamp 1669390400
transform 1 0 43344 0 1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output14
timestamp 1669390400
transform -1 0 44912 0 1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output15
timestamp 1669390400
transform 1 0 45360 0 1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output16
timestamp 1669390400
transform 1 0 45360 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output17
timestamp 1669390400
transform -1 0 44240 0 -1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output18
timestamp 1669390400
transform -1 0 44912 0 1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output19
timestamp 1669390400
transform -1 0 46368 0 -1 37632
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output20
timestamp 1669390400
transform 1 0 45360 0 1 37632
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output21
timestamp 1669390400
transform 1 0 44800 0 -1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output22
timestamp 1669390400
transform 1 0 45360 0 1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output23
timestamp 1669390400
transform 1 0 45360 0 1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output24
timestamp 1669390400
transform 1 0 45360 0 1 42336
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output25
timestamp 1669390400
transform 1 0 45360 0 1 43904
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output26
timestamp 1669390400
transform 1 0 44800 0 1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output27
timestamp 1669390400
transform 1 0 43344 0 1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output28
timestamp 1669390400
transform 1 0 44800 0 -1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output29
timestamp 1669390400
transform 1 0 46592 0 1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output30
timestamp 1669390400
transform 1 0 43344 0 1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output31
timestamp 1669390400
transform -1 0 46368 0 -1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output32
timestamp 1669390400
transform -1 0 46928 0 1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output33
timestamp 1669390400
transform 1 0 45360 0 1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output34
timestamp 1669390400
transform -1 0 46368 0 -1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output35
timestamp 1669390400
transform 1 0 46032 0 -1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output36
timestamp 1669390400
transform -1 0 43792 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output37
timestamp 1669390400
transform -1 0 3248 0 1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spi_core_38 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 8960 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spi_core_39
timestamp 1669390400
transform -1 0 14448 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spi_core_40
timestamp 1669390400
transform -1 0 19936 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spi_core_41
timestamp 1669390400
transform -1 0 25648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spi_core_42
timestamp 1669390400
transform -1 0 2128 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spi_core_43
timestamp 1669390400
transform -1 0 2128 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spi_core_44
timestamp 1669390400
transform -1 0 2128 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  spi_core_45 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 2128 0 1 45472
box -86 -86 534 870
<< labels >>
flabel metal2 s 2912 0 3024 800 0 FreeSans 448 90 0 0 clock
port 0 nsew signal input
flabel metal3 s 49200 1568 50000 1680 0 FreeSans 448 0 0 0 clock_out
port 1 nsew signal tristate
flabel metal3 s 49200 3024 50000 3136 0 FreeSans 448 0 0 0 data_out[0]
port 2 nsew signal tristate
flabel metal3 s 49200 17584 50000 17696 0 FreeSans 448 0 0 0 data_out[10]
port 3 nsew signal tristate
flabel metal3 s 49200 19040 50000 19152 0 FreeSans 448 0 0 0 data_out[11]
port 4 nsew signal tristate
flabel metal3 s 49200 20496 50000 20608 0 FreeSans 448 0 0 0 data_out[12]
port 5 nsew signal tristate
flabel metal3 s 49200 21952 50000 22064 0 FreeSans 448 0 0 0 data_out[13]
port 6 nsew signal tristate
flabel metal3 s 49200 23408 50000 23520 0 FreeSans 448 0 0 0 data_out[14]
port 7 nsew signal tristate
flabel metal3 s 49200 24864 50000 24976 0 FreeSans 448 0 0 0 data_out[15]
port 8 nsew signal tristate
flabel metal3 s 49200 26320 50000 26432 0 FreeSans 448 0 0 0 data_out[16]
port 9 nsew signal tristate
flabel metal3 s 49200 27776 50000 27888 0 FreeSans 448 0 0 0 data_out[17]
port 10 nsew signal tristate
flabel metal3 s 49200 29232 50000 29344 0 FreeSans 448 0 0 0 data_out[18]
port 11 nsew signal tristate
flabel metal3 s 49200 30688 50000 30800 0 FreeSans 448 0 0 0 data_out[19]
port 12 nsew signal tristate
flabel metal3 s 49200 4480 50000 4592 0 FreeSans 448 0 0 0 data_out[1]
port 13 nsew signal tristate
flabel metal3 s 49200 32144 50000 32256 0 FreeSans 448 0 0 0 data_out[20]
port 14 nsew signal tristate
flabel metal3 s 49200 33600 50000 33712 0 FreeSans 448 0 0 0 data_out[21]
port 15 nsew signal tristate
flabel metal3 s 49200 35056 50000 35168 0 FreeSans 448 0 0 0 data_out[22]
port 16 nsew signal tristate
flabel metal3 s 49200 36512 50000 36624 0 FreeSans 448 0 0 0 data_out[23]
port 17 nsew signal tristate
flabel metal3 s 49200 37968 50000 38080 0 FreeSans 448 0 0 0 data_out[24]
port 18 nsew signal tristate
flabel metal3 s 49200 39424 50000 39536 0 FreeSans 448 0 0 0 data_out[25]
port 19 nsew signal tristate
flabel metal3 s 49200 40880 50000 40992 0 FreeSans 448 0 0 0 data_out[26]
port 20 nsew signal tristate
flabel metal3 s 49200 42336 50000 42448 0 FreeSans 448 0 0 0 data_out[27]
port 21 nsew signal tristate
flabel metal3 s 49200 43792 50000 43904 0 FreeSans 448 0 0 0 data_out[28]
port 22 nsew signal tristate
flabel metal3 s 49200 45248 50000 45360 0 FreeSans 448 0 0 0 data_out[29]
port 23 nsew signal tristate
flabel metal3 s 49200 5936 50000 6048 0 FreeSans 448 0 0 0 data_out[2]
port 24 nsew signal tristate
flabel metal3 s 49200 46704 50000 46816 0 FreeSans 448 0 0 0 data_out[30]
port 25 nsew signal tristate
flabel metal3 s 49200 48160 50000 48272 0 FreeSans 448 0 0 0 data_out[31]
port 26 nsew signal tristate
flabel metal3 s 49200 7392 50000 7504 0 FreeSans 448 0 0 0 data_out[3]
port 27 nsew signal tristate
flabel metal3 s 49200 8848 50000 8960 0 FreeSans 448 0 0 0 data_out[4]
port 28 nsew signal tristate
flabel metal3 s 49200 10304 50000 10416 0 FreeSans 448 0 0 0 data_out[5]
port 29 nsew signal tristate
flabel metal3 s 49200 11760 50000 11872 0 FreeSans 448 0 0 0 data_out[6]
port 30 nsew signal tristate
flabel metal3 s 49200 13216 50000 13328 0 FreeSans 448 0 0 0 data_out[7]
port 31 nsew signal tristate
flabel metal3 s 49200 14672 50000 14784 0 FreeSans 448 0 0 0 data_out[8]
port 32 nsew signal tristate
flabel metal3 s 49200 16128 50000 16240 0 FreeSans 448 0 0 0 data_out[9]
port 33 nsew signal tristate
flabel metal2 s 30352 0 30464 800 0 FreeSans 448 90 0 0 la_data_in[0]
port 34 nsew signal input
flabel metal2 s 35840 0 35952 800 0 FreeSans 448 90 0 0 la_data_in[1]
port 35 nsew signal input
flabel metal2 s 41328 0 41440 800 0 FreeSans 448 90 0 0 la_data_in[2]
port 36 nsew signal input
flabel metal2 s 46816 0 46928 800 0 FreeSans 448 90 0 0 la_data_in[3]
port 37 nsew signal input
flabel metal2 s 8400 0 8512 800 0 FreeSans 448 90 0 0 la_oenb[0]
port 38 nsew signal tristate
flabel metal2 s 13888 0 14000 800 0 FreeSans 448 90 0 0 la_oenb[1]
port 39 nsew signal tristate
flabel metal2 s 19376 0 19488 800 0 FreeSans 448 90 0 0 la_oenb[2]
port 40 nsew signal tristate
flabel metal2 s 24864 0 24976 800 0 FreeSans 448 90 0 0 la_oenb[3]
port 41 nsew signal tristate
flabel metal3 s 0 40320 800 40432 0 FreeSans 448 0 0 0 miso
port 42 nsew signal tristate
flabel metal3 s 0 46480 800 46592 0 FreeSans 448 0 0 0 miso_oeb
port 43 nsew signal tristate
flabel metal3 s 0 15680 800 15792 0 FreeSans 448 0 0 0 mosi
port 44 nsew signal input
flabel metal3 s 0 21840 800 21952 0 FreeSans 448 0 0 0 mosi_oeb
port 45 nsew signal tristate
flabel metal3 s 0 3360 800 3472 0 FreeSans 448 0 0 0 sclk
port 46 nsew signal input
flabel metal3 s 0 9520 800 9632 0 FreeSans 448 0 0 0 sclk_oeb
port 47 nsew signal tristate
flabel metal3 s 0 28000 800 28112 0 FreeSans 448 0 0 0 ss_n
port 48 nsew signal input
flabel metal3 s 0 34160 800 34272 0 FreeSans 448 0 0 0 ss_n_oeb
port 49 nsew signal tristate
flabel metal4 s 4448 3076 4768 46316 0 FreeSans 1280 90 0 0 vdd
port 50 nsew power bidirectional
flabel metal4 s 35168 3076 35488 46316 0 FreeSans 1280 90 0 0 vdd
port 50 nsew power bidirectional
flabel metal4 s 19808 3076 20128 46316 0 FreeSans 1280 90 0 0 vss
port 51 nsew ground bidirectional
rlabel metal1 24976 46256 24976 46256 0 vdd
rlabel metal1 24976 45472 24976 45472 0 vss
rlabel metal2 34664 5600 34664 5600 0 _000_
rlabel metal3 36904 4424 36904 4424 0 _001_
rlabel metal2 38024 7784 38024 7784 0 _002_
rlabel metal2 39088 9912 39088 9912 0 _003_
rlabel metal3 47320 5992 47320 5992 0 _004_
rlabel metal3 45976 9128 45976 9128 0 _005_
rlabel metal2 43736 10920 43736 10920 0 _006_
rlabel metal2 44408 11648 44408 11648 0 _007_
rlabel metal2 43512 14168 43512 14168 0 _008_
rlabel metal3 42224 15512 42224 15512 0 _009_
rlabel metal3 46984 16968 46984 16968 0 _010_
rlabel metal2 44464 18536 44464 18536 0 _011_
rlabel metal2 44744 21056 44744 21056 0 _012_
rlabel metal3 46592 22120 46592 22120 0 _013_
rlabel metal2 45304 25032 45304 25032 0 _014_
rlabel metal2 42616 25760 42616 25760 0 _015_
rlabel metal2 38416 26488 38416 26488 0 _016_
rlabel metal2 37576 28168 37576 28168 0 _017_
rlabel metal3 45528 28056 45528 28056 0 _018_
rlabel metal2 43624 28000 43624 28000 0 _019_
rlabel metal2 44744 31304 44744 31304 0 _020_
rlabel metal3 45304 34216 45304 34216 0 _021_
rlabel metal2 45080 35896 45080 35896 0 _022_
rlabel metal2 45416 33376 45416 33376 0 _023_
rlabel metal3 42168 34216 42168 34216 0 _024_
rlabel metal2 40152 35392 40152 35392 0 _025_
rlabel metal3 37128 34776 37128 34776 0 _026_
rlabel metal3 35224 34216 35224 34216 0 _027_
rlabel metal2 38136 33208 38136 33208 0 _028_
rlabel metal2 36288 31640 36288 31640 0 _029_
rlabel metal2 32312 32984 32312 32984 0 _030_
rlabel metal2 30464 34328 30464 34328 0 _031_
rlabel metal3 45192 17864 45192 17864 0 _032_
rlabel metal3 45416 20664 45416 20664 0 _033_
rlabel metal3 45192 20776 45192 20776 0 _034_
rlabel metal2 47544 22344 47544 22344 0 _035_
rlabel metal2 45976 24472 45976 24472 0 _036_
rlabel metal2 43512 24304 43512 24304 0 _037_
rlabel metal2 40824 25536 40824 25536 0 _038_
rlabel metal2 46200 27720 46200 27720 0 _039_
rlabel metal2 38808 26712 38808 26712 0 _040_
rlabel metal2 39480 26600 39480 26600 0 _041_
rlabel metal2 46704 27272 46704 27272 0 _042_
rlabel metal2 42616 28560 42616 28560 0 _043_
rlabel metal3 46984 30072 46984 30072 0 _044_
rlabel metal3 45136 30184 45136 30184 0 _045_
rlabel metal3 45192 33544 45192 33544 0 _046_
rlabel metal3 45360 35112 45360 35112 0 _047_
rlabel metal3 47544 35672 47544 35672 0 _048_
rlabel metal2 40432 36344 40432 36344 0 _049_
rlabel metal2 41776 35672 41776 35672 0 _050_
rlabel metal2 40544 35784 40544 35784 0 _051_
rlabel metal2 37912 35560 37912 35560 0 _052_
rlabel metal2 35896 35112 35896 35112 0 _053_
rlabel metal3 38864 34104 38864 34104 0 _054_
rlabel metal2 37688 31836 37688 31836 0 _055_
rlabel metal2 35728 32312 35728 32312 0 _056_
rlabel metal2 32648 33824 32648 33824 0 _057_
rlabel metal2 33208 34440 33208 34440 0 _058_
rlabel metal2 34888 7336 34888 7336 0 _059_
rlabel metal2 22064 14728 22064 14728 0 _060_
rlabel metal2 21000 14504 21000 14504 0 _061_
rlabel metal2 40152 22624 40152 22624 0 _062_
rlabel metal2 44184 9408 44184 9408 0 _063_
rlabel metal3 39816 6664 39816 6664 0 _064_
rlabel metal2 35504 5992 35504 5992 0 _065_
rlabel metal2 37912 5376 37912 5376 0 _066_
rlabel metal2 38584 7504 38584 7504 0 _067_
rlabel metal2 39480 9464 39480 9464 0 _068_
rlabel metal2 46312 7448 46312 7448 0 _069_
rlabel metal2 47544 6664 47544 6664 0 _070_
rlabel metal2 47096 8736 47096 8736 0 _071_
rlabel metal3 45192 10808 45192 10808 0 _072_
rlabel metal3 45192 11256 45192 11256 0 _073_
rlabel metal2 46200 17640 46200 17640 0 _074_
rlabel metal3 44744 13832 44744 13832 0 _075_
rlabel metal3 43624 15288 43624 15288 0 _076_
rlabel metal2 46760 16688 46760 16688 0 _077_
rlabel metal2 30128 26936 30128 26936 0 clknet_0_clock
rlabel metal3 44128 7448 44128 7448 0 clknet_2_0__leaf_clock
rlabel metal2 21728 7672 21728 7672 0 clknet_2_1__leaf_clock
rlabel metal2 44632 23912 44632 23912 0 clknet_2_2__leaf_clock
rlabel metal2 5768 23072 5768 23072 0 clknet_2_3__leaf_clock
rlabel metal2 2968 2478 2968 2478 0 clock
rlabel metal2 45024 4424 45024 4424 0 clock_out
rlabel metal3 47698 3080 47698 3080 0 data_out[0]
rlabel metal3 46970 17640 46970 17640 0 data_out[10]
rlabel metal3 47978 19096 47978 19096 0 data_out[11]
rlabel metal3 47306 20552 47306 20552 0 data_out[12]
rlabel metal2 44072 22232 44072 22232 0 data_out[13]
rlabel metal3 47768 23184 47768 23184 0 data_out[14]
rlabel metal3 47978 24920 47978 24920 0 data_out[15]
rlabel metal3 47754 26376 47754 26376 0 data_out[16]
rlabel metal3 46970 27832 46970 27832 0 data_out[17]
rlabel metal2 44072 29792 44072 29792 0 data_out[18]
rlabel metal3 47978 30744 47978 30744 0 data_out[19]
rlabel metal3 48650 4536 48650 4536 0 data_out[1]
rlabel metal2 43288 32312 43288 32312 0 data_out[20]
rlabel metal2 44072 33544 44072 33544 0 data_out[21]
rlabel metal2 45304 36176 45304 36176 0 data_out[22]
rlabel metal3 47978 36568 47978 36568 0 data_out[23]
rlabel metal2 46088 38360 46088 38360 0 data_out[24]
rlabel metal3 47978 39480 47978 39480 0 data_out[25]
rlabel metal3 47978 40936 47978 40936 0 data_out[26]
rlabel metal3 47978 42392 47978 42392 0 data_out[27]
rlabel metal3 47978 43848 47978 43848 0 data_out[28]
rlabel metal3 47698 45304 47698 45304 0 data_out[29]
rlabel metal3 48650 5992 48650 5992 0 data_out[2]
rlabel metal2 45976 45864 45976 45864 0 data_out[30]
rlabel metal2 47880 47096 47880 47096 0 data_out[31]
rlabel metal3 46970 7448 46970 7448 0 data_out[3]
rlabel metal3 47306 8904 47306 8904 0 data_out[4]
rlabel metal2 46088 10136 46088 10136 0 data_out[5]
rlabel metal3 47978 11816 47978 11816 0 data_out[6]
rlabel metal2 45304 13440 45304 13440 0 data_out[7]
rlabel metal2 47320 14952 47320 14952 0 data_out[8]
rlabel metal3 49336 15680 49336 15680 0 data_out[9]
rlabel metal3 1358 40376 1358 40376 0 miso
rlabel metal2 1848 15624 1848 15624 0 mosi
rlabel metal2 9016 12936 9016 12936 0 mosi_reg\[0\]
rlabel metal2 26040 7952 26040 7952 0 mosi_reg\[1\]
rlabel metal2 25536 8344 25536 8344 0 mosi_reg\[2\]
rlabel metal3 5152 13832 5152 13832 0 net1
rlabel metal2 46312 24360 46312 24360 0 net10
rlabel metal2 44520 26544 44520 26544 0 net11
rlabel metal2 45080 26544 45080 26544 0 net12
rlabel metal2 45640 27608 45640 27608 0 net13
rlabel metal2 46760 29400 46760 29400 0 net14
rlabel metal2 46760 30184 46760 30184 0 net15
rlabel metal3 44912 5096 44912 5096 0 net16
rlabel metal2 46200 30464 46200 30464 0 net17
rlabel metal3 45528 33320 45528 33320 0 net18
rlabel metal2 46200 36792 46200 36792 0 net19
rlabel metal2 3360 3640 3360 3640 0 net2
rlabel metal2 48104 36008 48104 36008 0 net20
rlabel metal2 44968 37856 44968 37856 0 net21
rlabel metal2 44744 38416 44744 38416 0 net22
rlabel metal3 45136 41160 45136 41160 0 net23
rlabel metal2 44688 42504 44688 42504 0 net24
rlabel metal3 45136 44296 45136 44296 0 net25
rlabel metal2 44576 45864 44576 45864 0 net26
rlabel metal3 41832 7336 41832 7336 0 net27
rlabel metal2 44464 44968 44464 44968 0 net28
rlabel metal2 46536 44968 46536 44968 0 net29
rlabel metal2 6440 25088 6440 25088 0 net3
rlabel metal2 45976 6720 45976 6720 0 net30
rlabel metal3 45752 6776 45752 6776 0 net31
rlabel metal2 47376 7336 47376 7336 0 net32
rlabel metal2 45808 10472 45808 10472 0 net33
rlabel metal2 46368 13720 46368 13720 0 net34
rlabel metal2 45864 15400 45864 15400 0 net35
rlabel metal2 44072 16240 44072 16240 0 net36
rlabel metal2 3304 40880 3304 40880 0 net37
rlabel metal2 8456 2030 8456 2030 0 net38
rlabel metal2 13944 2030 13944 2030 0 net39
rlabel metal3 45976 4536 45976 4536 0 net4
rlabel metal2 19432 2030 19432 2030 0 net40
rlabel metal2 24920 2030 24920 2030 0 net41
rlabel metal3 1302 21896 1302 21896 0 net42
rlabel metal3 1302 9576 1302 9576 0 net43
rlabel metal3 1302 34216 1302 34216 0 net44
rlabel metal2 1848 46312 1848 46312 0 net45
rlabel metal3 44632 3528 44632 3528 0 net5
rlabel metal2 44184 17192 44184 17192 0 net6
rlabel metal2 46760 20412 46760 20412 0 net7
rlabel metal2 46200 21616 46200 21616 0 net8
rlabel metal3 45752 22344 45752 22344 0 net9
rlabel metal3 1358 3416 1358 3416 0 sclk
rlabel metal2 8680 5096 8680 5096 0 sclk_reg\[0\]
rlabel metal2 21000 15120 21000 15120 0 sclk_reg\[1\]
rlabel metal2 22288 13608 22288 13608 0 sclk_reg\[2\]
rlabel metal3 1302 28056 1302 28056 0 ss_n
rlabel metal2 8568 22736 8568 22736 0 ss_n_reg\[0\]
rlabel metal2 17864 14000 17864 14000 0 ss_n_reg\[1\]
rlabel metal2 19992 14504 19992 14504 0 ss_n_reg\[2\]
<< properties >>
string FIXED_BBOX 0 0 50000 50000
<< end >>

// This is the unpowered netlist.
module controller_core (clock,
    io_control_trigger_in,
    io_control_trigger_oeb,
    io_latch_data_in,
    io_latch_data_oeb,
    io_reset_n_in,
    io_reset_n_oeb,
    io_update_cycle_complete_oeb,
    io_update_cycle_complete_out,
    output_active_left,
    output_active_right,
    spi_data_clock,
    clock_out,
    col_select_left,
    col_select_right,
    data_out_left,
    data_out_right,
    inverter_select,
    io_driver_io_oeb,
    la_data_in,
    la_oenb,
    mem_address_left,
    mem_address_right,
    mem_write_n,
    row_col_select,
    row_select_left,
    row_select_right,
    spi_data);
 input clock;
 input io_control_trigger_in;
 output io_control_trigger_oeb;
 input io_latch_data_in;
 output io_latch_data_oeb;
 input io_reset_n_in;
 output io_reset_n_oeb;
 output io_update_cycle_complete_oeb;
 output io_update_cycle_complete_out;
 output output_active_left;
 output output_active_right;
 input spi_data_clock;
 output [9:0] clock_out;
 output [5:0] col_select_left;
 output [5:0] col_select_right;
 output [15:0] data_out_left;
 output [15:0] data_out_right;
 output [9:0] inverter_select;
 output [19:0] io_driver_io_oeb;
 input [17:0] la_data_in;
 input [17:0] la_oenb;
 output [9:0] mem_address_left;
 output [9:0] mem_address_right;
 output [9:0] mem_write_n;
 output [9:0] row_col_select;
 output [5:0] row_select_left;
 output [5:0] row_select_right;
 input [31:0] spi_data;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire control_trigger;
 wire \control_trigger_sync[0] ;
 wire \control_trigger_sync[1] ;
 wire latch_data;
 wire \latch_data_sync[0] ;
 wire \latch_data_sync[1] ;
 wire reset_n;
 wire \reset_n_sync[0] ;
 wire \reset_n_sync[1] ;
 wire \spi_data_crossing[0].A ;
 wire \spi_data_crossing[0].data_sync ;
 wire \spi_data_crossing[10].A ;
 wire \spi_data_crossing[10].data_sync ;
 wire \spi_data_crossing[11].A ;
 wire \spi_data_crossing[11].data_sync ;
 wire \spi_data_crossing[12].A ;
 wire \spi_data_crossing[12].data_sync ;
 wire \spi_data_crossing[13].A ;
 wire \spi_data_crossing[13].data_sync ;
 wire \spi_data_crossing[14].A ;
 wire \spi_data_crossing[14].data_sync ;
 wire \spi_data_crossing[15].A ;
 wire \spi_data_crossing[15].data_sync ;
 wire \spi_data_crossing[16].A ;
 wire \spi_data_crossing[16].data_sync ;
 wire \spi_data_crossing[17].A ;
 wire \spi_data_crossing[17].data_sync ;
 wire \spi_data_crossing[18].A ;
 wire \spi_data_crossing[18].data_sync ;
 wire \spi_data_crossing[19].A ;
 wire \spi_data_crossing[19].data_sync ;
 wire \spi_data_crossing[1].A ;
 wire \spi_data_crossing[1].data_sync ;
 wire \spi_data_crossing[20].A ;
 wire \spi_data_crossing[20].data_sync ;
 wire \spi_data_crossing[21].A ;
 wire \spi_data_crossing[21].data_sync ;
 wire \spi_data_crossing[22].A ;
 wire \spi_data_crossing[22].data_sync ;
 wire \spi_data_crossing[23].A ;
 wire \spi_data_crossing[23].data_sync ;
 wire \spi_data_crossing[24].A ;
 wire \spi_data_crossing[24].data_sync ;
 wire \spi_data_crossing[25].A ;
 wire \spi_data_crossing[25].data_sync ;
 wire \spi_data_crossing[26].A ;
 wire \spi_data_crossing[26].data_sync ;
 wire \spi_data_crossing[27].A ;
 wire \spi_data_crossing[27].data_sync ;
 wire \spi_data_crossing[28].A ;
 wire \spi_data_crossing[28].data_sync ;
 wire \spi_data_crossing[29].A ;
 wire \spi_data_crossing[29].data_sync ;
 wire \spi_data_crossing[2].A ;
 wire \spi_data_crossing[2].data_sync ;
 wire \spi_data_crossing[30].A ;
 wire \spi_data_crossing[30].data_sync ;
 wire \spi_data_crossing[31].A ;
 wire \spi_data_crossing[31].data_sync ;
 wire \spi_data_crossing[3].A ;
 wire \spi_data_crossing[3].data_sync ;
 wire \spi_data_crossing[4].A ;
 wire \spi_data_crossing[4].data_sync ;
 wire \spi_data_crossing[5].A ;
 wire \spi_data_crossing[5].data_sync ;
 wire \spi_data_crossing[6].A ;
 wire \spi_data_crossing[6].data_sync ;
 wire \spi_data_crossing[7].A ;
 wire \spi_data_crossing[7].data_sync ;
 wire \spi_data_crossing[8].A ;
 wire \spi_data_crossing[8].data_sync ;
 wire \spi_data_crossing[9].A ;
 wire \spi_data_crossing[9].data_sync ;
 wire \u0.cmd[0] ;
 wire \u0.cmd[10] ;
 wire \u0.cmd[11] ;
 wire \u0.cmd[12] ;
 wire \u0.cmd[13] ;
 wire \u0.cmd[14] ;
 wire \u0.cmd[15] ;
 wire \u0.cmd[16] ;
 wire \u0.cmd[17] ;
 wire \u0.cmd[18] ;
 wire \u0.cmd[19] ;
 wire \u0.cmd[1] ;
 wire \u0.cmd[20] ;
 wire \u0.cmd[21] ;
 wire \u0.cmd[22] ;
 wire \u0.cmd[23] ;
 wire \u0.cmd[24] ;
 wire \u0.cmd[25] ;
 wire \u0.cmd[26] ;
 wire \u0.cmd[27] ;
 wire \u0.cmd[28] ;
 wire \u0.cmd[29] ;
 wire \u0.cmd[2] ;
 wire \u0.cmd[30] ;
 wire \u0.cmd[31] ;
 wire \u0.cmd[3] ;
 wire \u0.cmd[4] ;
 wire \u0.cmd[5] ;
 wire \u0.cmd[6] ;
 wire \u0.cmd[7] ;
 wire \u0.cmd[8] ;
 wire \u0.cmd[9] ;
 wire \u0.latch_cmd ;
 wire \u0.mem_write_n[0] ;
 wire \u0.mem_write_n[1] ;
 wire \u0.mem_write_n[2] ;
 wire \u0.mem_write_n[3] ;
 wire \u0.mem_write_n[4] ;
 wire \u0.mem_write_n[5] ;
 wire \u0.mem_write_n[6] ;
 wire \u0.mem_write_n[7] ;
 wire \u0.mem_write_n[8] ;
 wire \u0.mem_write_n[9] ;
 wire \u0.run_state[0] ;
 wire \u0.run_state[1] ;
 wire \u0.run_state[2] ;
 wire \u0.run_state[3] ;
 wire \u0.run_state[4] ;
 wire \u0.run_state[5] ;
 wire \u0.run_state[6] ;
 wire \u0.timer_enable ;
 wire \u0.u11.impulse_gen[0] ;
 wire \u0.u11.impulse_gen[1] ;
 wire \u0.update_cmd ;
 wire \u0.write_config_n ;
 wire \u1.ccr0[0] ;
 wire \u1.ccr0[10] ;
 wire \u1.ccr0[11] ;
 wire \u1.ccr0[12] ;
 wire \u1.ccr0[13] ;
 wire \u1.ccr0[14] ;
 wire \u1.ccr0[15] ;
 wire \u1.ccr0[16] ;
 wire \u1.ccr0[17] ;
 wire \u1.ccr0[18] ;
 wire \u1.ccr0[19] ;
 wire \u1.ccr0[1] ;
 wire \u1.ccr0[20] ;
 wire \u1.ccr0[21] ;
 wire \u1.ccr0[22] ;
 wire \u1.ccr0[23] ;
 wire \u1.ccr0[24] ;
 wire \u1.ccr0[25] ;
 wire \u1.ccr0[26] ;
 wire \u1.ccr0[27] ;
 wire \u1.ccr0[28] ;
 wire \u1.ccr0[29] ;
 wire \u1.ccr0[2] ;
 wire \u1.ccr0[30] ;
 wire \u1.ccr0[31] ;
 wire \u1.ccr0[3] ;
 wire \u1.ccr0[4] ;
 wire \u1.ccr0[5] ;
 wire \u1.ccr0[6] ;
 wire \u1.ccr0[7] ;
 wire \u1.ccr0[8] ;
 wire \u1.ccr0[9] ;
 wire \u1.ccr1[0] ;
 wire \u1.ccr1[10] ;
 wire \u1.ccr1[11] ;
 wire \u1.ccr1[12] ;
 wire \u1.ccr1[13] ;
 wire \u1.ccr1[14] ;
 wire \u1.ccr1[15] ;
 wire \u1.ccr1[16] ;
 wire \u1.ccr1[17] ;
 wire \u1.ccr1[18] ;
 wire \u1.ccr1[19] ;
 wire \u1.ccr1[1] ;
 wire \u1.ccr1[20] ;
 wire \u1.ccr1[21] ;
 wire \u1.ccr1[22] ;
 wire \u1.ccr1[23] ;
 wire \u1.ccr1[24] ;
 wire \u1.ccr1[25] ;
 wire \u1.ccr1[26] ;
 wire \u1.ccr1[27] ;
 wire \u1.ccr1[28] ;
 wire \u1.ccr1[29] ;
 wire \u1.ccr1[2] ;
 wire \u1.ccr1[30] ;
 wire \u1.ccr1[31] ;
 wire \u1.ccr1[3] ;
 wire \u1.ccr1[4] ;
 wire \u1.ccr1[5] ;
 wire \u1.ccr1[6] ;
 wire \u1.ccr1[7] ;
 wire \u1.ccr1[8] ;
 wire \u1.ccr1[9] ;
 wire \u1.ccr1_flag ;
 wire \u1.col_limit[0] ;
 wire \u1.col_limit[1] ;
 wire \u1.col_limit[2] ;
 wire \u1.col_limit[3] ;
 wire \u1.col_limit[4] ;
 wire \u1.col_limit[5] ;
 wire \u1.col_limit[6] ;
 wire \u1.col_sel[0] ;
 wire \u1.col_sel[1] ;
 wire \u1.col_sel[2] ;
 wire \u1.col_sel[3] ;
 wire \u1.col_sel[4] ;
 wire \u1.col_sel[5] ;
 wire \u1.col_sel[6] ;
 wire \u1.inverter_select[0] ;
 wire \u1.inverter_select[1] ;
 wire \u1.inverter_select[2] ;
 wire \u1.inverter_select[3] ;
 wire \u1.inverter_select[4] ;
 wire \u1.inverter_select[5] ;
 wire \u1.inverter_select[6] ;
 wire \u1.inverter_select[7] ;
 wire \u1.inverter_select[8] ;
 wire \u1.inverter_select[9] ;
 wire \u1.ordering_complete[0] ;
 wire \u1.ordering_complete[10] ;
 wire \u1.ordering_complete[11] ;
 wire \u1.ordering_complete[12] ;
 wire \u1.ordering_complete[13] ;
 wire \u1.ordering_complete[14] ;
 wire \u1.ordering_complete[15] ;
 wire \u1.ordering_complete[16] ;
 wire \u1.ordering_complete[17] ;
 wire \u1.ordering_complete[18] ;
 wire \u1.ordering_complete[19] ;
 wire \u1.ordering_complete[1] ;
 wire \u1.ordering_complete[20] ;
 wire \u1.ordering_complete[21] ;
 wire \u1.ordering_complete[22] ;
 wire \u1.ordering_complete[23] ;
 wire \u1.ordering_complete[24] ;
 wire \u1.ordering_complete[25] ;
 wire \u1.ordering_complete[26] ;
 wire \u1.ordering_complete[27] ;
 wire \u1.ordering_complete[28] ;
 wire \u1.ordering_complete[29] ;
 wire \u1.ordering_complete[2] ;
 wire \u1.ordering_complete[30] ;
 wire \u1.ordering_complete[31] ;
 wire \u1.ordering_complete[3] ;
 wire \u1.ordering_complete[4] ;
 wire \u1.ordering_complete[5] ;
 wire \u1.ordering_complete[6] ;
 wire \u1.ordering_complete[7] ;
 wire \u1.ordering_complete[8] ;
 wire \u1.ordering_complete[9] ;
 wire \u1.ordering_timer[0] ;
 wire \u1.ordering_timer[10] ;
 wire \u1.ordering_timer[11] ;
 wire \u1.ordering_timer[12] ;
 wire \u1.ordering_timer[13] ;
 wire \u1.ordering_timer[14] ;
 wire \u1.ordering_timer[15] ;
 wire \u1.ordering_timer[16] ;
 wire \u1.ordering_timer[17] ;
 wire \u1.ordering_timer[18] ;
 wire \u1.ordering_timer[19] ;
 wire \u1.ordering_timer[1] ;
 wire \u1.ordering_timer[20] ;
 wire \u1.ordering_timer[21] ;
 wire \u1.ordering_timer[22] ;
 wire \u1.ordering_timer[23] ;
 wire \u1.ordering_timer[24] ;
 wire \u1.ordering_timer[25] ;
 wire \u1.ordering_timer[26] ;
 wire \u1.ordering_timer[27] ;
 wire \u1.ordering_timer[28] ;
 wire \u1.ordering_timer[29] ;
 wire \u1.ordering_timer[2] ;
 wire \u1.ordering_timer[30] ;
 wire \u1.ordering_timer[31] ;
 wire \u1.ordering_timer[3] ;
 wire \u1.ordering_timer[4] ;
 wire \u1.ordering_timer[5] ;
 wire \u1.ordering_timer[6] ;
 wire \u1.ordering_timer[7] ;
 wire \u1.ordering_timer[8] ;
 wire \u1.ordering_timer[9] ;
 wire \u1.output_active ;
 wire \u1.row_col_select[0] ;
 wire \u1.row_col_select[1] ;
 wire \u1.row_col_select[2] ;
 wire \u1.row_col_select[3] ;
 wire \u1.row_col_select[4] ;
 wire \u1.row_col_select[5] ;
 wire \u1.row_col_select[6] ;
 wire \u1.row_col_select[7] ;
 wire \u1.row_col_select[8] ;
 wire \u1.row_col_select[9] ;
 wire \u1.row_limit[0] ;
 wire \u1.row_limit[1] ;
 wire \u1.row_limit[2] ;
 wire \u1.row_limit[3] ;
 wire \u1.row_limit[4] ;
 wire \u1.row_limit[5] ;
 wire \u1.row_limit[6] ;
 wire \u1.row_sel[0] ;
 wire \u1.row_sel[1] ;
 wire \u1.row_sel[2] ;
 wire \u1.row_sel[3] ;
 wire \u1.row_sel[4] ;
 wire \u1.row_sel[5] ;
 wire \u1.row_sel[6] ;
 wire \u1.timer[0] ;
 wire \u1.timer[10] ;
 wire \u1.timer[11] ;
 wire \u1.timer[12] ;
 wire \u1.timer[13] ;
 wire \u1.timer[14] ;
 wire \u1.timer[15] ;
 wire \u1.timer[16] ;
 wire \u1.timer[17] ;
 wire \u1.timer[18] ;
 wire \u1.timer[19] ;
 wire \u1.timer[1] ;
 wire \u1.timer[20] ;
 wire \u1.timer[21] ;
 wire \u1.timer[22] ;
 wire \u1.timer[23] ;
 wire \u1.timer[24] ;
 wire \u1.timer[25] ;
 wire \u1.timer[26] ;
 wire \u1.timer[27] ;
 wire \u1.timer[28] ;
 wire \u1.timer[29] ;
 wire \u1.timer[2] ;
 wire \u1.timer[30] ;
 wire \u1.timer[31] ;
 wire \u1.timer[3] ;
 wire \u1.timer[4] ;
 wire \u1.timer[5] ;
 wire \u1.timer[6] ;
 wire \u1.timer[7] ;
 wire \u1.timer[8] ;
 wire \u1.timer[9] ;
 wire \u1.u1.impulse_gen[0] ;
 wire \u1.u1.impulse_gen[1] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire clknet_leaf_0_clock;
 wire clknet_leaf_1_clock;
 wire clknet_leaf_2_clock;
 wire clknet_leaf_3_clock;
 wire clknet_leaf_4_clock;
 wire clknet_leaf_5_clock;
 wire clknet_leaf_6_clock;
 wire clknet_leaf_7_clock;
 wire clknet_leaf_8_clock;
 wire clknet_leaf_9_clock;
 wire clknet_leaf_10_clock;
 wire clknet_leaf_11_clock;
 wire clknet_leaf_12_clock;
 wire clknet_leaf_13_clock;
 wire clknet_leaf_14_clock;
 wire clknet_leaf_15_clock;
 wire clknet_leaf_16_clock;
 wire clknet_leaf_17_clock;
 wire clknet_leaf_18_clock;
 wire clknet_leaf_19_clock;
 wire clknet_leaf_20_clock;
 wire clknet_leaf_21_clock;
 wire clknet_leaf_22_clock;
 wire clknet_leaf_23_clock;
 wire clknet_leaf_24_clock;
 wire clknet_leaf_25_clock;
 wire clknet_leaf_26_clock;
 wire clknet_leaf_27_clock;
 wire clknet_leaf_28_clock;
 wire clknet_leaf_29_clock;
 wire clknet_leaf_30_clock;
 wire clknet_leaf_31_clock;
 wire clknet_leaf_32_clock;
 wire clknet_leaf_33_clock;
 wire clknet_leaf_34_clock;
 wire clknet_leaf_35_clock;
 wire clknet_leaf_36_clock;
 wire clknet_0_clock;
 wire clknet_2_0__leaf_clock;
 wire clknet_2_1__leaf_clock;
 wire clknet_2_2__leaf_clock;
 wire clknet_2_3__leaf_clock;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;

 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1415_ (.I(\u0.cmd[31] ),
    .Z(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1416_ (.A1(\reset_n_sync[1] ),
    .A2(\reset_n_sync[0] ),
    .A3(reset_n),
    .Z(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1417_ (.I(_1041_),
    .Z(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1418_ (.A1(_1040_),
    .A2(\u0.cmd[30] ),
    .A3(_1042_),
    .ZN(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1419_ (.A1(\control_trigger_sync[0] ),
    .A2(control_trigger),
    .A3(\control_trigger_sync[1] ),
    .Z(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1420_ (.A1(\u0.cmd[26] ),
    .A2(_1044_),
    .ZN(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1421_ (.I(\u1.ordering_timer[23] ),
    .ZN(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1422_ (.I(\u1.ordering_timer[22] ),
    .ZN(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1423_ (.A1(_1046_),
    .A2(\u1.ordering_complete[23] ),
    .B1(_1047_),
    .B2(\u1.ordering_complete[22] ),
    .ZN(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1424_ (.I(\u1.ordering_timer[21] ),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1425_ (.I(\u1.ordering_timer[20] ),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1426_ (.A1(_1049_),
    .A2(\u1.ordering_complete[21] ),
    .B1(_1050_),
    .B2(\u1.ordering_complete[20] ),
    .ZN(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1427_ (.A1(_1048_),
    .A2(_1051_),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1428_ (.A1(_1047_),
    .A2(\u1.ordering_complete[22] ),
    .B1(_1049_),
    .B2(\u1.ordering_complete[21] ),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1429_ (.I(\u1.ordering_complete[23] ),
    .ZN(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1430_ (.A1(\u1.ordering_timer[23] ),
    .A2(_1054_),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1431_ (.A1(_1050_),
    .A2(\u1.ordering_complete[20] ),
    .B(_1055_),
    .ZN(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1432_ (.A1(_1052_),
    .A2(_1053_),
    .A3(_1056_),
    .ZN(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1433_ (.I(\u1.ordering_complete[19] ),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1434_ (.I(\u1.ordering_timer[16] ),
    .Z(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1435_ (.I(\u1.ordering_complete[16] ),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1436_ (.I(\u1.ordering_complete[17] ),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1437_ (.A1(\u1.ordering_timer[17] ),
    .A2(_1061_),
    .B1(\u1.ordering_timer[16] ),
    .B2(_1060_),
    .ZN(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _1438_ (.A1(\u1.ordering_timer[19] ),
    .A2(_1058_),
    .B1(_1059_),
    .B2(_1060_),
    .C(_1062_),
    .ZN(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1439_ (.I(\u1.ordering_timer[19] ),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1440_ (.I(\u1.ordering_timer[18] ),
    .ZN(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _1441_ (.A1(_1064_),
    .A2(\u1.ordering_complete[19] ),
    .B1(_1065_),
    .B2(\u1.ordering_complete[18] ),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1442_ (.I(\u1.ordering_complete[18] ),
    .ZN(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1443_ (.I(\u1.ordering_timer[17] ),
    .Z(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _1444_ (.A1(\u1.ordering_timer[18] ),
    .A2(_1067_),
    .B1(_1068_),
    .B2(_1061_),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1445_ (.A1(_1057_),
    .A2(_1063_),
    .A3(_1066_),
    .A4(_1069_),
    .ZN(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1446_ (.I(\u1.ordering_timer[28] ),
    .ZN(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1447_ (.I(\u1.ordering_timer[27] ),
    .ZN(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1448_ (.I(\u1.ordering_complete[31] ),
    .ZN(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1449_ (.A1(\u1.ordering_timer[31] ),
    .A2(_1073_),
    .ZN(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _1450_ (.A1(_1071_),
    .A2(\u1.ordering_complete[28] ),
    .B1(_1072_),
    .B2(\u1.ordering_complete[27] ),
    .C(_1074_),
    .ZN(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1451_ (.I(\u1.ordering_timer[29] ),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1452_ (.A1(_1076_),
    .A2(\u1.ordering_complete[29] ),
    .B1(_1071_),
    .B2(\u1.ordering_complete[28] ),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1453_ (.I(\u1.ordering_complete[30] ),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1454_ (.I(\u1.ordering_complete[29] ),
    .ZN(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1455_ (.A1(\u1.ordering_timer[30] ),
    .A2(_1078_),
    .B1(\u1.ordering_timer[29] ),
    .B2(_1079_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1456_ (.A1(_1077_),
    .A2(_1080_),
    .ZN(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1457_ (.I(\u1.ordering_timer[30] ),
    .Z(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1458_ (.A1(\u1.ordering_timer[31] ),
    .A2(_1073_),
    .B1(_1082_),
    .B2(_1078_),
    .ZN(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1459_ (.A1(_1075_),
    .A2(_1081_),
    .A3(_1083_),
    .ZN(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1460_ (.I(\u1.ordering_timer[24] ),
    .Z(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1461_ (.I(\u1.ordering_complete[24] ),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1462_ (.I(\u1.ordering_timer[26] ),
    .ZN(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1463_ (.I(\u1.ordering_timer[25] ),
    .ZN(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1464_ (.A1(_1087_),
    .A2(\u1.ordering_complete[26] ),
    .B1(_1088_),
    .B2(\u1.ordering_complete[25] ),
    .ZN(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1465_ (.A1(_1085_),
    .A2(_1086_),
    .B(_1089_),
    .ZN(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1466_ (.A1(\u1.ordering_timer[24] ),
    .A2(_1086_),
    .ZN(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1467_ (.A1(_1088_),
    .A2(\u1.ordering_complete[25] ),
    .B(_1091_),
    .ZN(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1468_ (.I(_1072_),
    .Z(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _1469_ (.A1(_1093_),
    .A2(\u1.ordering_complete[27] ),
    .B1(_1087_),
    .B2(\u1.ordering_complete[26] ),
    .ZN(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1470_ (.A1(_1084_),
    .A2(_1090_),
    .A3(_1092_),
    .A4(_1094_),
    .ZN(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1471_ (.I(\u1.ordering_timer[15] ),
    .Z(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1472_ (.I(\u1.ordering_complete[15] ),
    .ZN(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1473_ (.I(\u1.ordering_complete[14] ),
    .ZN(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1474_ (.A1(_1096_),
    .A2(_1097_),
    .B1(\u1.ordering_timer[14] ),
    .B2(_1098_),
    .ZN(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1475_ (.I(\u1.ordering_timer[14] ),
    .ZN(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1476_ (.I(\u1.ordering_timer[13] ),
    .ZN(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1477_ (.A1(_1100_),
    .A2(\u1.ordering_complete[14] ),
    .B1(_1101_),
    .B2(\u1.ordering_complete[13] ),
    .ZN(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1478_ (.I(\u1.ordering_timer[12] ),
    .ZN(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1479_ (.I(\u1.ordering_complete[11] ),
    .ZN(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1480_ (.A1(\u1.ordering_timer[15] ),
    .A2(_1097_),
    .B1(\u1.ordering_timer[11] ),
    .B2(_1104_),
    .ZN(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1481_ (.A1(_1101_),
    .A2(\u1.ordering_complete[13] ),
    .B1(_1103_),
    .B2(\u1.ordering_complete[12] ),
    .ZN(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1482_ (.A1(_1103_),
    .A2(\u1.ordering_complete[12] ),
    .B(_1105_),
    .C(_1106_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1483_ (.A1(_1099_),
    .A2(_1102_),
    .A3(_1107_),
    .ZN(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1484_ (.I(\u1.ordering_timer[9] ),
    .ZN(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1485_ (.I(\u1.ordering_complete[9] ),
    .Z(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1486_ (.I(\u1.ordering_timer[8] ),
    .ZN(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1487_ (.I(\u1.ordering_complete[8] ),
    .Z(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1488_ (.I(\u1.ordering_complete[10] ),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1489_ (.A1(\u1.ordering_timer[11] ),
    .A2(_1104_),
    .B1(\u1.ordering_timer[10] ),
    .B2(_1113_),
    .ZN(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _1490_ (.A1(_1109_),
    .A2(_1110_),
    .B1(_1111_),
    .B2(_1112_),
    .C(_1114_),
    .ZN(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1491_ (.I(\u1.ordering_timer[10] ),
    .ZN(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1492_ (.A1(_1116_),
    .A2(\u1.ordering_complete[10] ),
    .B1(_1109_),
    .B2(\u1.ordering_complete[9] ),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1493_ (.A1(_1111_),
    .A2(_1112_),
    .ZN(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1494_ (.A1(_1117_),
    .A2(_1118_),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1495_ (.A1(_1108_),
    .A2(_1115_),
    .A3(_1119_),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1496_ (.I(\u1.ordering_timer[5] ),
    .ZN(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1497_ (.I(\u1.ordering_timer[4] ),
    .ZN(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1498_ (.A1(_1121_),
    .A2(\u1.ordering_complete[5] ),
    .B1(_1122_),
    .B2(\u1.ordering_complete[4] ),
    .ZN(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1499_ (.I(\u1.ordering_timer[7] ),
    .ZN(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1500_ (.I(\u1.ordering_timer[6] ),
    .ZN(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1501_ (.A1(_1124_),
    .A2(\u1.ordering_complete[7] ),
    .B1(_1125_),
    .B2(\u1.ordering_complete[6] ),
    .ZN(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1502_ (.A1(_1123_),
    .A2(_1126_),
    .ZN(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1503_ (.I(\u1.ordering_timer[3] ),
    .ZN(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1504_ (.A1(_1124_),
    .A2(\u1.ordering_complete[7] ),
    .Z(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _1505_ (.A1(_1128_),
    .A2(\u1.ordering_complete[3] ),
    .B1(_1122_),
    .B2(\u1.ordering_complete[4] ),
    .C(_1129_),
    .ZN(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1506_ (.A1(_1125_),
    .A2(\u1.ordering_complete[6] ),
    .B1(_1121_),
    .B2(\u1.ordering_complete[5] ),
    .ZN(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1507_ (.A1(_1127_),
    .A2(_1130_),
    .A3(_1131_),
    .ZN(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1508_ (.I(\u1.ordering_complete[0] ),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1509_ (.I(\u1.ordering_complete[1] ),
    .ZN(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _1510_ (.A1(\u1.ordering_timer[0] ),
    .A2(_1133_),
    .B1(\u1.ordering_timer[1] ),
    .B2(_1134_),
    .ZN(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1511_ (.I(\u1.ordering_timer[2] ),
    .ZN(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _1512_ (.A1(_1128_),
    .A2(\u1.ordering_complete[3] ),
    .B1(_1136_),
    .B2(\u1.ordering_complete[2] ),
    .ZN(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1513_ (.I(\u1.ordering_timer[0] ),
    .Z(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1514_ (.I(_1138_),
    .ZN(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1515_ (.A1(\u1.ordering_timer[1] ),
    .A2(_1134_),
    .ZN(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1516_ (.A1(_1136_),
    .A2(\u1.ordering_complete[2] ),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1517_ (.A1(_1139_),
    .A2(\u1.ordering_complete[0] ),
    .B(_1140_),
    .C(_1141_),
    .ZN(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1518_ (.A1(_1132_),
    .A2(_1135_),
    .A3(_1137_),
    .A4(_1142_),
    .ZN(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _1519_ (.A1(_1070_),
    .A2(_1095_),
    .A3(_1120_),
    .A4(_1143_),
    .ZN(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1520_ (.I(_1144_),
    .ZN(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1521_ (.A1(\u0.run_state[6] ),
    .A2(_1045_),
    .B1(_1145_),
    .B2(\u0.run_state[3] ),
    .ZN(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1522_ (.A1(_1043_),
    .A2(_1146_),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1523_ (.A1(\control_trigger_sync[0] ),
    .A2(control_trigger),
    .A3(\control_trigger_sync[1] ),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1524_ (.A1(\u0.cmd[28] ),
    .A2(\u0.run_state[2] ),
    .B1(_1147_),
    .B2(\u0.run_state[5] ),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1525_ (.A1(_1043_),
    .A2(_1148_),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1526_ (.I(\u0.cmd[27] ),
    .ZN(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1527_ (.A1(\u0.run_state[5] ),
    .A2(_1044_),
    .B(\u0.run_state[1] ),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1528_ (.A1(_1149_),
    .A2(_1150_),
    .ZN(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1529_ (.A1(\u0.run_state[4] ),
    .A2(_1151_),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1530_ (.A1(_1043_),
    .A2(_1152_),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1531_ (.I(\u0.cmd[29] ),
    .Z(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1532_ (.I(\u0.run_state[0] ),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1533_ (.A1(_1040_),
    .A2(\u0.cmd[30] ),
    .A3(_1042_),
    .Z(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1534_ (.A1(_1153_),
    .A2(_1154_),
    .B(_1155_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1535_ (.I(\u0.u11.impulse_gen[0] ),
    .ZN(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1536_ (.A1(_1156_),
    .A2(\u0.u11.impulse_gen[1] ),
    .ZN(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1537_ (.I(_1157_),
    .Z(\u0.latch_cmd ));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1538_ (.A1(\u0.run_state[3] ),
    .A2(\u0.run_state[4] ),
    .Z(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1539_ (.I(_1158_),
    .Z(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1540_ (.I(\u0.run_state[6] ),
    .ZN(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1541_ (.I(\u0.cmd[27] ),
    .Z(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1542_ (.A1(_1159_),
    .A2(_1045_),
    .B1(_1150_),
    .B2(_1160_),
    .ZN(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1543_ (.A1(\u0.run_state[3] ),
    .A2(_1144_),
    .B(_1161_),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1544_ (.A1(_1043_),
    .A2(_1162_),
    .ZN(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1545_ (.I(\u1.timer[25] ),
    .ZN(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1546_ (.I(_1163_),
    .Z(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1547_ (.I(\u1.timer[24] ),
    .ZN(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1548_ (.I(_1165_),
    .Z(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1549_ (.I(\u1.timer[30] ),
    .ZN(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1550_ (.I(\u1.timer[29] ),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1551_ (.A1(\u1.ccr1[30] ),
    .A2(_1167_),
    .B1(\u1.ccr1[29] ),
    .B2(_1168_),
    .ZN(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _1552_ (.A1(\u1.ccr1[25] ),
    .A2(_1164_),
    .B1(\u1.ccr1[24] ),
    .B2(_1166_),
    .C(_1169_),
    .ZN(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1553_ (.I(\u1.timer[31] ),
    .ZN(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1554_ (.A1(\u1.ccr1[31] ),
    .A2(_1171_),
    .B1(\u1.ccr1[30] ),
    .B2(_1167_),
    .ZN(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1555_ (.I(\u1.timer[28] ),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1556_ (.A1(\u1.ccr1[29] ),
    .A2(_1168_),
    .B1(\u1.ccr1[28] ),
    .B2(_1173_),
    .ZN(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1557_ (.A1(_1172_),
    .A2(_1174_),
    .Z(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1558_ (.I(\u1.ccr1[27] ),
    .ZN(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1559_ (.I(\u1.timer[27] ),
    .Z(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1560_ (.I(\u1.ccr1[26] ),
    .ZN(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1561_ (.A1(_1176_),
    .A2(\u1.timer[27] ),
    .B1(_1178_),
    .B2(\u1.timer[26] ),
    .ZN(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1562_ (.I(\u1.timer[26] ),
    .ZN(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1563_ (.A1(\u1.ccr1[26] ),
    .A2(_1180_),
    .ZN(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1564_ (.A1(_1176_),
    .A2(_1177_),
    .B(_1179_),
    .C(_1181_),
    .ZN(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1565_ (.A1(\u1.ccr1[25] ),
    .A2(_1163_),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1566_ (.A1(\u1.ccr1[28] ),
    .A2(_1173_),
    .B1(\u1.ccr1[24] ),
    .B2(_1165_),
    .ZN(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1567_ (.A1(\u1.ccr1[31] ),
    .A2(_1171_),
    .ZN(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1568_ (.A1(_1183_),
    .A2(_1184_),
    .A3(_1185_),
    .ZN(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1569_ (.A1(_1170_),
    .A2(_1175_),
    .A3(_1182_),
    .A4(_1186_),
    .ZN(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1570_ (.I(\u1.timer[6] ),
    .Z(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1571_ (.I(_1188_),
    .ZN(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1572_ (.I(\u1.timer[5] ),
    .Z(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1573_ (.I(_1190_),
    .ZN(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1574_ (.A1(\u1.ccr1[6] ),
    .A2(_1189_),
    .B1(\u1.ccr1[5] ),
    .B2(_1191_),
    .ZN(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1575_ (.I(\u1.timer[7] ),
    .ZN(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1576_ (.I(\u1.timer[4] ),
    .ZN(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1577_ (.A1(\u1.ccr1[7] ),
    .A2(_1193_),
    .B1(\u1.ccr1[4] ),
    .B2(_1194_),
    .ZN(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1578_ (.I(\u1.ccr1[5] ),
    .ZN(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1579_ (.I(\u1.ccr1[4] ),
    .ZN(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1580_ (.A1(_1196_),
    .A2(_1190_),
    .B1(_1197_),
    .B2(\u1.timer[4] ),
    .ZN(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1581_ (.I(\u1.ccr1[7] ),
    .ZN(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1582_ (.I(\u1.ccr1[6] ),
    .ZN(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1583_ (.A1(_1199_),
    .A2(\u1.timer[7] ),
    .B1(_1200_),
    .B2(_1188_),
    .ZN(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _1584_ (.A1(_1192_),
    .A2(_1195_),
    .A3(_1198_),
    .A4(_1201_),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1585_ (.I(\u1.timer[2] ),
    .Z(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1586_ (.I(_1203_),
    .ZN(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1587_ (.A1(\u1.ccr1[2] ),
    .A2(_1204_),
    .ZN(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1588_ (.I(\u1.timer[0] ),
    .Z(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1589_ (.I(_1206_),
    .ZN(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1590_ (.I(\u1.timer[1] ),
    .Z(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1591_ (.I(_1208_),
    .ZN(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1592_ (.A1(_1207_),
    .A2(\u1.ccr1[0] ),
    .B1(\u1.ccr1[1] ),
    .B2(_1209_),
    .ZN(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1593_ (.A1(_1205_),
    .A2(_1210_),
    .ZN(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1594_ (.I(\u0.timer_enable ),
    .Z(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1595_ (.I(\u1.ccr1[3] ),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1596_ (.I(\u1.timer[3] ),
    .Z(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1597_ (.I(\u1.ccr1[2] ),
    .ZN(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1598_ (.A1(_1213_),
    .A2(_1214_),
    .B1(_1215_),
    .B2(_1203_),
    .ZN(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1599_ (.A1(_1207_),
    .A2(\u1.ccr1[0] ),
    .Z(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1600_ (.A1(\u1.ccr1[1] ),
    .A2(_1209_),
    .ZN(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1601_ (.A1(_1213_),
    .A2(\u1.timer[3] ),
    .ZN(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1602_ (.A1(_1218_),
    .A2(_1219_),
    .ZN(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1603_ (.A1(_1212_),
    .A2(_1216_),
    .A3(_1217_),
    .A4(_1220_),
    .ZN(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1604_ (.A1(_1202_),
    .A2(_1211_),
    .A3(_1221_),
    .ZN(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1605_ (.I(\u1.timer[20] ),
    .ZN(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1606_ (.I(_1223_),
    .Z(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1607_ (.I(\u1.ccr1[23] ),
    .ZN(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1608_ (.I(\u1.ccr1[22] ),
    .ZN(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1609_ (.A1(_1225_),
    .A2(\u1.timer[23] ),
    .B1(_1226_),
    .B2(\u1.timer[22] ),
    .ZN(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1610_ (.I(\u1.timer[23] ),
    .ZN(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1611_ (.I(\u1.timer[22] ),
    .ZN(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1612_ (.I(\u1.timer[21] ),
    .ZN(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _1613_ (.A1(\u1.ccr1[23] ),
    .A2(_1228_),
    .B1(\u1.ccr1[22] ),
    .B2(_1229_),
    .C1(\u1.ccr1[21] ),
    .C2(_1230_),
    .ZN(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1614_ (.A1(_1227_),
    .A2(_1231_),
    .ZN(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1615_ (.I(_1230_),
    .Z(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1616_ (.A1(\u1.ccr1[21] ),
    .A2(_1233_),
    .B1(\u1.ccr1[20] ),
    .B2(_1223_),
    .ZN(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1617_ (.A1(\u1.ccr1[20] ),
    .A2(_1224_),
    .B(_1232_),
    .C(_1234_),
    .ZN(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1618_ (.I(\u1.timer[17] ),
    .ZN(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1619_ (.I(\u1.timer[16] ),
    .ZN(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1620_ (.A1(\u1.ccr1[17] ),
    .A2(_1236_),
    .B1(\u1.ccr1[16] ),
    .B2(_1237_),
    .ZN(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1621_ (.A1(\u1.ccr1[19] ),
    .A2(\u1.timer[19] ),
    .Z(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1622_ (.A1(\u1.ccr1[18] ),
    .A2(\u1.timer[18] ),
    .Z(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1623_ (.A1(_1239_),
    .A2(_1240_),
    .ZN(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1624_ (.A1(\u1.ccr1[17] ),
    .A2(_1236_),
    .ZN(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1625_ (.A1(\u1.ccr1[16] ),
    .A2(_1237_),
    .ZN(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1626_ (.A1(_1241_),
    .A2(_1242_),
    .A3(_1243_),
    .ZN(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1627_ (.A1(_1238_),
    .A2(_1244_),
    .ZN(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1628_ (.A1(_1235_),
    .A2(_1245_),
    .ZN(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1629_ (.I(\u1.ccr1[9] ),
    .ZN(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1630_ (.I(\u1.timer[9] ),
    .Z(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1631_ (.I(\u1.ccr1[8] ),
    .ZN(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1632_ (.I(\u1.timer[8] ),
    .Z(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1633_ (.A1(_1247_),
    .A2(_1248_),
    .B1(_1249_),
    .B2(_1250_),
    .ZN(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1634_ (.I(\u1.ccr1[15] ),
    .ZN(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1635_ (.I(\u1.ccr1[14] ),
    .ZN(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1636_ (.I(\u1.timer[14] ),
    .Z(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1637_ (.A1(_1252_),
    .A2(\u1.timer[15] ),
    .B1(_1253_),
    .B2(_1254_),
    .ZN(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1638_ (.I(\u1.timer[15] ),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1639_ (.I(\u1.timer[14] ),
    .ZN(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1640_ (.I(\u1.timer[13] ),
    .ZN(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _1641_ (.A1(\u1.ccr1[15] ),
    .A2(_1256_),
    .B1(\u1.ccr1[14] ),
    .B2(_1257_),
    .C1(\u1.ccr1[13] ),
    .C2(_1258_),
    .ZN(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1642_ (.A1(_1255_),
    .A2(_1259_),
    .ZN(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1643_ (.I(\u1.ccr1[12] ),
    .ZN(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1644_ (.I(\u1.timer[12] ),
    .Z(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1645_ (.I(\u1.ccr1[13] ),
    .ZN(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1646_ (.A1(_1263_),
    .A2(\u1.timer[13] ),
    .B1(_1261_),
    .B2(\u1.timer[12] ),
    .ZN(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1647_ (.A1(_1261_),
    .A2(_1262_),
    .B(_1264_),
    .ZN(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1648_ (.A1(_1260_),
    .A2(_1265_),
    .ZN(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1649_ (.I(\u1.timer[8] ),
    .ZN(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1650_ (.I(\u1.timer[10] ),
    .ZN(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1651_ (.I(\u1.timer[11] ),
    .ZN(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1652_ (.A1(\u1.ccr1[11] ),
    .A2(_1269_),
    .ZN(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1653_ (.I(\u1.ccr1[11] ),
    .ZN(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1654_ (.I(\u1.timer[11] ),
    .Z(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1655_ (.A1(_1271_),
    .A2(_1272_),
    .B1(\u1.ccr1[10] ),
    .B2(_1268_),
    .ZN(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1656_ (.A1(\u1.ccr1[10] ),
    .A2(_1268_),
    .B(_1270_),
    .C(_1273_),
    .ZN(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1657_ (.A1(_1247_),
    .A2(_1248_),
    .ZN(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1658_ (.A1(\u1.ccr1[8] ),
    .A2(_1267_),
    .B(_1274_),
    .C(_1275_),
    .ZN(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1659_ (.A1(_1251_),
    .A2(_1266_),
    .A3(_1276_),
    .ZN(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1660_ (.A1(_1246_),
    .A2(_1277_),
    .ZN(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1661_ (.A1(_1187_),
    .A2(_1222_),
    .A3(_1278_),
    .ZN(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1662_ (.I(_1279_),
    .ZN(\u1.ccr1_flag ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1663_ (.I(_1188_),
    .Z(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1664_ (.I(\u1.ccr0[6] ),
    .ZN(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1665_ (.I(\u1.ccr0[5] ),
    .ZN(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1666_ (.I(_1190_),
    .Z(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1667_ (.A1(_1280_),
    .A2(_1281_),
    .B1(_1282_),
    .B2(_1283_),
    .ZN(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1668_ (.A1(_1193_),
    .A2(\u1.ccr0[7] ),
    .B1(\u1.ccr0[4] ),
    .B2(_1194_),
    .C(_1284_),
    .ZN(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1669_ (.I(\u1.ccr0[4] ),
    .ZN(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1670_ (.I(\u1.timer[4] ),
    .Z(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1671_ (.A1(_1283_),
    .A2(_1282_),
    .B1(_1286_),
    .B2(_1287_),
    .ZN(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1672_ (.I(\u1.timer[7] ),
    .Z(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1673_ (.I(\u1.ccr0[7] ),
    .ZN(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1674_ (.A1(_1289_),
    .A2(_1290_),
    .B1(_1281_),
    .B2(_1280_),
    .ZN(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1675_ (.A1(_1285_),
    .A2(_1288_),
    .A3(_1291_),
    .Z(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1676_ (.I(\u1.timer[9] ),
    .ZN(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _1677_ (.A1(_1269_),
    .A2(\u1.ccr0[11] ),
    .B1(\u1.ccr0[10] ),
    .B2(_1268_),
    .ZN(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1678_ (.I(\u1.timer[10] ),
    .Z(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1679_ (.I(\u1.ccr0[10] ),
    .ZN(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1680_ (.A1(_1269_),
    .A2(\u1.ccr0[11] ),
    .ZN(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1681_ (.A1(_1295_),
    .A2(_1296_),
    .B(_1297_),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1682_ (.A1(_1293_),
    .A2(\u1.ccr0[9] ),
    .B(_1294_),
    .C(_1298_),
    .ZN(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1683_ (.I(\u1.timer[13] ),
    .Z(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1684_ (.I(\u1.ccr0[13] ),
    .ZN(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1685_ (.A1(_1300_),
    .A2(_1301_),
    .ZN(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1686_ (.I(\u1.timer[15] ),
    .Z(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1687_ (.I(\u1.ccr0[15] ),
    .ZN(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1688_ (.I(\u1.ccr0[14] ),
    .ZN(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1689_ (.A1(_1303_),
    .A2(_1304_),
    .B1(_1305_),
    .B2(_1254_),
    .ZN(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1690_ (.A1(_1256_),
    .A2(\u1.ccr0[15] ),
    .B1(\u1.ccr0[14] ),
    .B2(_1257_),
    .ZN(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1691_ (.A1(_1306_),
    .A2(_1307_),
    .ZN(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1692_ (.A1(_1293_),
    .A2(\u1.ccr0[9] ),
    .B1(\u1.ccr0[8] ),
    .B2(_1267_),
    .ZN(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1693_ (.I(\u1.ccr0[12] ),
    .ZN(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1694_ (.I(_1262_),
    .Z(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1695_ (.A1(_1300_),
    .A2(_1301_),
    .B1(_1310_),
    .B2(_1311_),
    .ZN(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1696_ (.A1(_1262_),
    .A2(_1310_),
    .ZN(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1697_ (.A1(_1267_),
    .A2(\u1.ccr0[8] ),
    .B(_1313_),
    .ZN(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1698_ (.A1(_1312_),
    .A2(_1314_),
    .ZN(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _1699_ (.A1(_1302_),
    .A2(_1308_),
    .A3(_1309_),
    .A4(_1315_),
    .ZN(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1700_ (.A1(_1299_),
    .A2(_1316_),
    .ZN(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1701_ (.I(\u1.timer[19] ),
    .Z(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1702_ (.I(\u1.ccr0[19] ),
    .ZN(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1703_ (.I(\u1.ccr0[18] ),
    .ZN(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1704_ (.I(\u1.timer[18] ),
    .Z(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1705_ (.I(_1321_),
    .Z(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1706_ (.A1(_1318_),
    .A2(_1319_),
    .B1(_1320_),
    .B2(_1322_),
    .ZN(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1707_ (.A1(_1321_),
    .A2(_1320_),
    .ZN(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1708_ (.A1(_1318_),
    .A2(_1319_),
    .ZN(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1709_ (.A1(_1324_),
    .A2(_1325_),
    .ZN(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1710_ (.I(\u1.timer[23] ),
    .Z(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1711_ (.I(\u1.ccr0[23] ),
    .ZN(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1712_ (.I(\u1.ccr0[22] ),
    .ZN(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1713_ (.A1(_1327_),
    .A2(_1328_),
    .B1(_1329_),
    .B2(\u1.timer[22] ),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1714_ (.A1(_1327_),
    .A2(_1328_),
    .ZN(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1715_ (.A1(_1229_),
    .A2(\u1.ccr0[22] ),
    .B(_1331_),
    .ZN(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1716_ (.A1(_1330_),
    .A2(_1332_),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1717_ (.A1(_1236_),
    .A2(\u1.ccr0[17] ),
    .B1(\u1.ccr0[16] ),
    .B2(_1237_),
    .ZN(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1718_ (.A1(_1233_),
    .A2(\u1.ccr0[21] ),
    .B1(\u1.ccr0[20] ),
    .B2(_1224_),
    .ZN(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1719_ (.A1(_1236_),
    .A2(\u1.ccr0[17] ),
    .ZN(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1720_ (.A1(_1233_),
    .A2(\u1.ccr0[21] ),
    .ZN(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1721_ (.A1(_1224_),
    .A2(\u1.ccr0[20] ),
    .ZN(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1722_ (.A1(_1237_),
    .A2(\u1.ccr0[16] ),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1723_ (.A1(_1336_),
    .A2(_1337_),
    .A3(_1338_),
    .A4(_1339_),
    .ZN(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1724_ (.A1(_1333_),
    .A2(_1334_),
    .A3(_1335_),
    .A4(_1340_),
    .ZN(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1725_ (.A1(_1323_),
    .A2(_1326_),
    .A3(_1341_),
    .ZN(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1726_ (.I(\u1.ccr0[27] ),
    .ZN(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1727_ (.I(\u1.ccr0[26] ),
    .ZN(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1728_ (.I(\u1.timer[26] ),
    .Z(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1729_ (.A1(_1177_),
    .A2(_1343_),
    .B1(_1344_),
    .B2(_1345_),
    .ZN(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _1730_ (.A1(_1164_),
    .A2(\u1.ccr0[25] ),
    .B1(\u1.ccr0[24] ),
    .B2(_1166_),
    .C(_1346_),
    .ZN(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1731_ (.A1(_1180_),
    .A2(\u1.ccr0[26] ),
    .B1(\u1.ccr0[25] ),
    .B2(_1164_),
    .ZN(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1732_ (.I(_1177_),
    .ZN(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1733_ (.A1(_1173_),
    .A2(\u1.ccr0[28] ),
    .B1(\u1.ccr0[27] ),
    .B2(_1349_),
    .ZN(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1734_ (.I(\u1.timer[31] ),
    .Z(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1735_ (.I(\u1.ccr0[31] ),
    .ZN(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1736_ (.I(\u1.ccr0[30] ),
    .ZN(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1737_ (.A1(_1351_),
    .A2(_1352_),
    .B1(_1353_),
    .B2(\u1.timer[30] ),
    .ZN(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1738_ (.A1(_1171_),
    .A2(\u1.ccr0[31] ),
    .B1(\u1.ccr0[24] ),
    .B2(_1166_),
    .ZN(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1739_ (.A1(_1348_),
    .A2(_1350_),
    .A3(_1354_),
    .A4(_1355_),
    .ZN(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1740_ (.I(\u1.ccr0[29] ),
    .ZN(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1741_ (.I(\u1.ccr0[28] ),
    .ZN(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1742_ (.A1(\u1.timer[29] ),
    .A2(_1357_),
    .B1(_1358_),
    .B2(\u1.timer[28] ),
    .ZN(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1743_ (.A1(_1167_),
    .A2(\u1.ccr0[30] ),
    .B1(\u1.ccr0[29] ),
    .B2(_1168_),
    .ZN(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1744_ (.A1(_1359_),
    .A2(_1360_),
    .ZN(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1745_ (.A1(_1347_),
    .A2(_1356_),
    .A3(_1361_),
    .ZN(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1746_ (.I(_1209_),
    .Z(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1747_ (.I(_1207_),
    .Z(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1748_ (.A1(_1363_),
    .A2(\u1.ccr0[1] ),
    .B1(\u1.ccr0[0] ),
    .B2(_1364_),
    .ZN(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1749_ (.A1(_1363_),
    .A2(\u1.ccr0[1] ),
    .B(_1365_),
    .ZN(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1750_ (.I(_1214_),
    .ZN(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1751_ (.A1(_1367_),
    .A2(\u1.ccr0[3] ),
    .B1(\u1.ccr0[2] ),
    .B2(_1204_),
    .ZN(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1752_ (.A1(_1367_),
    .A2(\u1.ccr0[3] ),
    .ZN(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1753_ (.A1(_1204_),
    .A2(\u1.ccr0[2] ),
    .ZN(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1754_ (.A1(_1364_),
    .A2(\u1.ccr0[0] ),
    .B(_1369_),
    .C(_1370_),
    .ZN(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1755_ (.A1(_1366_),
    .A2(_1368_),
    .A3(_1371_),
    .ZN(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1756_ (.A1(_1362_),
    .A2(_1372_),
    .ZN(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1757_ (.A1(_1317_),
    .A2(_1342_),
    .A3(_1373_),
    .ZN(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1758_ (.A1(_1299_),
    .A2(_1316_),
    .Z(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1759_ (.A1(_1363_),
    .A2(\u1.ccr0[1] ),
    .B(_1366_),
    .ZN(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1760_ (.A1(_1370_),
    .A2(_1376_),
    .B(_1368_),
    .ZN(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1761_ (.A1(_1292_),
    .A2(_1369_),
    .ZN(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1762_ (.A1(_1284_),
    .A2(_1288_),
    .B(_1291_),
    .ZN(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1763_ (.A1(_1289_),
    .A2(_1290_),
    .B(_1379_),
    .ZN(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1764_ (.A1(_1377_),
    .A2(_1378_),
    .B(_1380_),
    .ZN(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1765_ (.A1(_1294_),
    .A2(_1297_),
    .B1(_1299_),
    .B2(_1309_),
    .ZN(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1766_ (.A1(_1313_),
    .A2(_1382_),
    .B(_1312_),
    .ZN(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1767_ (.A1(_1302_),
    .A2(_1308_),
    .ZN(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1768_ (.A1(_1256_),
    .A2(\u1.ccr0[15] ),
    .B(_1306_),
    .ZN(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _1769_ (.A1(_1375_),
    .A2(_1381_),
    .B1(_1383_),
    .B2(_1384_),
    .C(_1385_),
    .ZN(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1770_ (.A1(_1323_),
    .A2(_1326_),
    .ZN(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1771_ (.A1(_1336_),
    .A2(_1334_),
    .ZN(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1772_ (.A1(_1323_),
    .A2(_1325_),
    .B1(_1387_),
    .B2(_1388_),
    .ZN(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1773_ (.A1(_1338_),
    .A2(_1389_),
    .B(_1335_),
    .ZN(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1774_ (.A1(_1333_),
    .A2(_1390_),
    .ZN(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1775_ (.A1(_1337_),
    .A2(_1391_),
    .ZN(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1776_ (.A1(_1330_),
    .A2(_1331_),
    .B1(_1342_),
    .B2(_1386_),
    .C(_1392_),
    .ZN(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1777_ (.I(_1177_),
    .Z(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1778_ (.A1(_1394_),
    .A2(_1343_),
    .B1(_1344_),
    .B2(_1345_),
    .C(_1348_),
    .ZN(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1779_ (.A1(_1350_),
    .A2(_1347_),
    .ZN(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1780_ (.A1(_1395_),
    .A2(_1396_),
    .B(_1359_),
    .ZN(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1781_ (.A1(_1360_),
    .A2(_1397_),
    .ZN(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1782_ (.A1(_1171_),
    .A2(\u1.ccr0[31] ),
    .B1(_1354_),
    .B2(_1398_),
    .ZN(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1783_ (.A1(_1362_),
    .A2(_1393_),
    .B(_1399_),
    .ZN(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1784_ (.A1(_1292_),
    .A2(_1374_),
    .B(_1400_),
    .ZN(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1785_ (.I(_1212_),
    .Z(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1786_ (.A1(_1402_),
    .A2(_1144_),
    .ZN(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1787_ (.I(_1311_),
    .ZN(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1788_ (.A1(_1256_),
    .A2(_1257_),
    .A3(_1258_),
    .A4(_1404_),
    .ZN(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1789_ (.A1(_1289_),
    .A2(_1280_),
    .A3(_1283_),
    .A4(_1287_),
    .ZN(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1790_ (.A1(_1206_),
    .A2(_1208_),
    .A3(_1214_),
    .A4(_1203_),
    .ZN(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1791_ (.A1(_1272_),
    .A2(_1295_),
    .A3(_1248_),
    .A4(_1250_),
    .ZN(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1792_ (.A1(_1406_),
    .A2(_1407_),
    .A3(_1408_),
    .ZN(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1793_ (.I(_1345_),
    .Z(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1794_ (.I(\u1.timer[25] ),
    .Z(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1795_ (.A1(_1394_),
    .A2(_1410_),
    .A3(_1411_),
    .A4(\u1.timer[24] ),
    .ZN(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1796_ (.I(\u1.timer[28] ),
    .Z(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1797_ (.A1(_1351_),
    .A2(\u1.timer[30] ),
    .A3(\u1.timer[29] ),
    .A4(_1413_),
    .ZN(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1798_ (.A1(_1412_),
    .A2(_1414_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1799_ (.I(_1318_),
    .Z(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1800_ (.I(\u1.timer[17] ),
    .Z(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1801_ (.I(\u1.timer[16] ),
    .Z(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1802_ (.A1(_0281_),
    .A2(_1322_),
    .A3(_0282_),
    .A4(_0283_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1803_ (.I(_1327_),
    .Z(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1804_ (.I(\u1.timer[22] ),
    .Z(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1805_ (.A1(_0285_),
    .A2(_0286_),
    .A3(\u1.timer[21] ),
    .A4(\u1.timer[20] ),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1806_ (.A1(_0284_),
    .A2(_0287_),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1807_ (.A1(_1405_),
    .A2(_1409_),
    .A3(_0280_),
    .A4(_0288_),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1808_ (.A1(_1401_),
    .A2(_1403_),
    .A3(_0289_),
    .ZN(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1809_ (.I0(net16),
    .I1(net3),
    .S(net34),
    .Z(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1810_ (.I(_0290_),
    .Z(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1811_ (.I0(net17),
    .I1(net2),
    .S(net35),
    .Z(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1812_ (.I(_0291_),
    .Z(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1813_ (.I0(net18),
    .I1(net1),
    .S(net36),
    .Z(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1814_ (.I(_0292_),
    .Z(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1815_ (.A1(net19),
    .A2(net37),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1816_ (.A1(net37),
    .A2(_1144_),
    .B(_0293_),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1817_ (.A1(_1153_),
    .A2(\u0.run_state[0] ),
    .A3(_1155_),
    .Z(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1818_ (.I(_0294_),
    .Z(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1819_ (.I(\u0.cmd[30] ),
    .ZN(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1820_ (.A1(_1040_),
    .A2(_0295_),
    .A3(\u0.update_cmd ),
    .ZN(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1821_ (.A1(\u0.cmd[28] ),
    .A2(\u0.cmd[29] ),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1822_ (.A1(_0295_),
    .A2(\u0.update_cmd ),
    .ZN(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1823_ (.A1(\u0.cmd[31] ),
    .A2(\u0.cmd[26] ),
    .A3(\u0.cmd[27] ),
    .A4(_0297_),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1824_ (.A1(_0296_),
    .A2(_0298_),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1825_ (.I(\u0.cmd[26] ),
    .Z(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1826_ (.A1(\u0.cmd[31] ),
    .A2(_0297_),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1827_ (.A1(_0299_),
    .A2(_1149_),
    .A3(_0300_),
    .Z(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1828_ (.A1(_0296_),
    .A2(_0301_),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1829_ (.I(_0300_),
    .Z(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1830_ (.A1(\u0.cmd[26] ),
    .A2(_1149_),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1831_ (.A1(_0296_),
    .A2(_0302_),
    .A3(_0303_),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1832_ (.A1(_0299_),
    .A2(_1160_),
    .A3(_0296_),
    .A4(_0302_),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1833_ (.I(\u0.cmd[28] ),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1834_ (.A1(_0304_),
    .A2(\u0.cmd[29] ),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1835_ (.A1(_0298_),
    .A2(_0305_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1836_ (.A1(_0301_),
    .A2(_0305_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1837_ (.A1(_0302_),
    .A2(_0303_),
    .A3(_0305_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1838_ (.A1(_0299_),
    .A2(_1160_),
    .A3(_0302_),
    .A4(_0305_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1839_ (.A1(_0304_),
    .A2(_1153_),
    .A3(_0298_),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1840_ (.A1(_0304_),
    .A2(_1153_),
    .A3(_0301_),
    .ZN(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1841_ (.A1(_0304_),
    .A2(\u0.run_state[2] ),
    .A3(_1155_),
    .Z(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1842_ (.I(_0306_),
    .Z(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1843_ (.I(net15),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1844_ (.A1(_0307_),
    .A2(net33),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1845_ (.I(\u1.u1.impulse_gen[1] ),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1846_ (.A1(\u1.u1.impulse_gen[0] ),
    .A2(_0308_),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1847_ (.I(\u1.col_limit[6] ),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1848_ (.I(\u1.col_sel[5] ),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1849_ (.A1(_0311_),
    .A2(\u1.col_limit[5] ),
    .Z(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1850_ (.I(\u1.col_sel[3] ),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1851_ (.I(\u1.col_sel[4] ),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1852_ (.A1(_0313_),
    .A2(\u1.col_limit[3] ),
    .B1(_0314_),
    .B2(\u1.col_limit[4] ),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1853_ (.I(\u1.col_sel[2] ),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1854_ (.I(\u1.col_sel[1] ),
    .Z(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1855_ (.I(\u1.col_limit[1] ),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1856_ (.I(\u1.col_limit[2] ),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1857_ (.A1(_0317_),
    .A2(_0318_),
    .B1(net225),
    .B2(_0319_),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1858_ (.I(\u1.col_limit[0] ),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1859_ (.A1(net226),
    .A2(_0321_),
    .B1(\u1.col_sel[1] ),
    .B2(_0318_),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _1860_ (.A1(_0313_),
    .A2(\u1.col_limit[3] ),
    .B1(_0316_),
    .B2(\u1.col_limit[2] ),
    .C1(_0320_),
    .C2(_0322_),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1861_ (.A1(_0311_),
    .A2(\u1.col_limit[5] ),
    .B1(_0314_),
    .B2(\u1.col_limit[4] ),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1862_ (.A1(_0315_),
    .A2(_0323_),
    .B(_0324_),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1863_ (.A1(\u1.col_sel[6] ),
    .A2(\u1.col_limit[6] ),
    .Z(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1864_ (.A1(_0312_),
    .A2(_0325_),
    .B(_0326_),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1865_ (.A1(\u1.col_sel[6] ),
    .A2(_0310_),
    .B(_0327_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1866_ (.I(_1402_),
    .Z(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1867_ (.A1(_0309_),
    .A2(_0328_),
    .B(_0329_),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1868_ (.I(_0330_),
    .Z(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1869_ (.A1(\u0.timer_enable ),
    .A2(_0309_),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1870_ (.A1(net226),
    .A2(_0332_),
    .Z(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1871_ (.A1(net226),
    .A2(_0332_),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1872_ (.A1(_0331_),
    .A2(_0333_),
    .A3(_0334_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1873_ (.A1(_0317_),
    .A2(_0333_),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1874_ (.A1(_0331_),
    .A2(_0335_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1875_ (.A1(_0317_),
    .A2(net225),
    .A3(_0333_),
    .Z(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1876_ (.A1(_0317_),
    .A2(_0333_),
    .B(net225),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1877_ (.A1(_0330_),
    .A2(_0336_),
    .A3(_0337_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1878_ (.A1(\u1.col_sel[3] ),
    .A2(_0336_),
    .Z(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1879_ (.A1(\u1.col_sel[3] ),
    .A2(_0336_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1880_ (.A1(_0330_),
    .A2(_0338_),
    .A3(_0339_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1881_ (.A1(\u1.col_sel[4] ),
    .A2(_0338_),
    .Z(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1882_ (.A1(\u1.col_sel[4] ),
    .A2(_0338_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1883_ (.A1(_0330_),
    .A2(_0340_),
    .A3(_0341_),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1884_ (.A1(_0311_),
    .A2(_0340_),
    .Z(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1885_ (.A1(_0331_),
    .A2(_0342_),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1886_ (.A1(\u1.col_sel[5] ),
    .A2(_0340_),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1887_ (.A1(\u1.col_sel[6] ),
    .A2(_0343_),
    .Z(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1888_ (.A1(_0331_),
    .A2(_0344_),
    .ZN(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1889_ (.I(\u0.cmd[0] ),
    .Z(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1890_ (.I(_0345_),
    .Z(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1891_ (.I(\u0.cmd[16] ),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1892_ (.I(\u0.cmd[17] ),
    .Z(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1893_ (.I(net218),
    .ZN(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1894_ (.A1(\u0.write_config_n ),
    .A2(\u0.cmd[18] ),
    .A3(\u0.cmd[21] ),
    .A4(\u0.cmd[20] ),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1895_ (.A1(_0349_),
    .A2(_0350_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1896_ (.A1(_0347_),
    .A2(_0348_),
    .A3(_0351_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1897_ (.I(_0352_),
    .Z(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1898_ (.I(_0353_),
    .Z(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1899_ (.I0(\u1.ccr0[16] ),
    .I1(_0346_),
    .S(_0354_),
    .Z(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1900_ (.I(_0355_),
    .Z(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1901_ (.I(\u0.cmd[1] ),
    .Z(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1902_ (.I(_0356_),
    .Z(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1903_ (.I0(\u1.ccr0[17] ),
    .I1(_0357_),
    .S(_0354_),
    .Z(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1904_ (.I(_0358_),
    .Z(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1905_ (.I(_0352_),
    .Z(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1906_ (.I(_0359_),
    .Z(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1907_ (.I(\u0.cmd[2] ),
    .Z(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1908_ (.I(_0353_),
    .Z(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1909_ (.A1(_0361_),
    .A2(_0362_),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1910_ (.A1(_1320_),
    .A2(_0360_),
    .B(_0363_),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1911_ (.I(\u0.cmd[3] ),
    .Z(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1912_ (.A1(_0364_),
    .A2(_0362_),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1913_ (.A1(_1319_),
    .A2(_0360_),
    .B(_0365_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1914_ (.I(\u0.cmd[4] ),
    .Z(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1915_ (.I0(\u1.ccr0[20] ),
    .I1(_0366_),
    .S(_0354_),
    .Z(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1916_ (.I(_0367_),
    .Z(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1917_ (.I(\u0.cmd[5] ),
    .Z(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1918_ (.I0(\u1.ccr0[21] ),
    .I1(_0368_),
    .S(_0354_),
    .Z(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1919_ (.I(_0369_),
    .Z(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1920_ (.I(\u0.cmd[6] ),
    .Z(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1921_ (.I(_0353_),
    .Z(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1922_ (.A1(_0370_),
    .A2(_0371_),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1923_ (.A1(_1329_),
    .A2(_0360_),
    .B(_0372_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1924_ (.I(\u0.cmd[7] ),
    .Z(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1925_ (.A1(_0373_),
    .A2(_0371_),
    .ZN(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1926_ (.A1(_1328_),
    .A2(_0360_),
    .B(_0374_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1927_ (.I(\u0.cmd[8] ),
    .Z(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1928_ (.I0(\u1.ccr0[24] ),
    .I1(_0375_),
    .S(_0359_),
    .Z(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1929_ (.I(_0376_),
    .Z(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1930_ (.I(\u0.cmd[9] ),
    .Z(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1931_ (.I0(\u1.ccr0[25] ),
    .I1(_0377_),
    .S(_0359_),
    .Z(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1932_ (.I(_0378_),
    .Z(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1933_ (.I(_0359_),
    .Z(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1934_ (.I(net224),
    .Z(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1935_ (.A1(_0380_),
    .A2(_0371_),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1936_ (.A1(_1344_),
    .A2(_0379_),
    .B(_0381_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1937_ (.I(net223),
    .Z(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1938_ (.A1(_0382_),
    .A2(_0371_),
    .ZN(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1939_ (.A1(_1343_),
    .A2(_0379_),
    .B(_0383_),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1940_ (.I(_0353_),
    .Z(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1941_ (.A1(net222),
    .A2(_0384_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1942_ (.A1(_1358_),
    .A2(_0379_),
    .B(_0385_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1943_ (.I(net221),
    .Z(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1944_ (.A1(_0386_),
    .A2(_0384_),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1945_ (.A1(_1357_),
    .A2(_0379_),
    .B(_0387_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1946_ (.I(net220),
    .Z(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1947_ (.A1(_0388_),
    .A2(_0384_),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1948_ (.A1(_1353_),
    .A2(_0362_),
    .B(_0389_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1949_ (.I(net219),
    .Z(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1950_ (.A1(_0390_),
    .A2(_0384_),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1951_ (.A1(_1352_),
    .A2(_0362_),
    .B(_0391_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1952_ (.I(\u0.cmd[0] ),
    .Z(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1953_ (.I(\u0.cmd[16] ),
    .Z(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1954_ (.I(\u0.cmd[17] ),
    .Z(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1955_ (.I(_0394_),
    .ZN(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1956_ (.A1(_0393_),
    .A2(_0395_),
    .A3(_0351_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1957_ (.I(_0396_),
    .Z(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1958_ (.I(_0397_),
    .Z(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1959_ (.I0(\u1.ccr1[0] ),
    .I1(_0392_),
    .S(_0398_),
    .Z(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1960_ (.I(_0399_),
    .Z(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1961_ (.I(\u0.cmd[1] ),
    .Z(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1962_ (.I0(\u1.ccr1[1] ),
    .I1(_0400_),
    .S(_0398_),
    .Z(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1963_ (.I(_0401_),
    .Z(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1964_ (.I(_0397_),
    .Z(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1965_ (.I(_0402_),
    .Z(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1966_ (.I(\u0.cmd[2] ),
    .Z(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1967_ (.I(_0396_),
    .Z(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1968_ (.A1(_0404_),
    .A2(_0405_),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1969_ (.A1(_1215_),
    .A2(_0403_),
    .B(_0406_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1970_ (.I(\u0.cmd[3] ),
    .Z(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1971_ (.A1(_0407_),
    .A2(_0405_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1972_ (.A1(_1213_),
    .A2(_0403_),
    .B(_0408_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1973_ (.I(\u0.cmd[4] ),
    .Z(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1974_ (.A1(_0409_),
    .A2(_0405_),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1975_ (.A1(_1197_),
    .A2(_0403_),
    .B(_0410_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1976_ (.I(\u0.cmd[5] ),
    .Z(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1977_ (.I(_0397_),
    .Z(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1978_ (.A1(_0411_),
    .A2(_0412_),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1979_ (.A1(_1196_),
    .A2(_0403_),
    .B(_0413_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1980_ (.I(_0402_),
    .Z(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1981_ (.A1(_0370_),
    .A2(_0412_),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1982_ (.A1(_1200_),
    .A2(_0414_),
    .B(_0415_),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1983_ (.A1(_0373_),
    .A2(_0412_),
    .ZN(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1984_ (.A1(_1199_),
    .A2(_0414_),
    .B(_0416_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1985_ (.A1(\u0.cmd[8] ),
    .A2(_0412_),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1986_ (.A1(_1249_),
    .A2(_0414_),
    .B(_0417_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1987_ (.I(_0397_),
    .Z(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1988_ (.A1(\u0.cmd[9] ),
    .A2(_0418_),
    .ZN(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1989_ (.A1(_1247_),
    .A2(_0414_),
    .B(_0419_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1990_ (.I0(\u1.ccr1[10] ),
    .I1(_0380_),
    .S(_0402_),
    .Z(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1991_ (.I(_0420_),
    .Z(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1992_ (.I(_0402_),
    .Z(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1993_ (.A1(_0382_),
    .A2(_0418_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1994_ (.A1(_1271_),
    .A2(_0421_),
    .B(_0422_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1995_ (.A1(net222),
    .A2(_0418_),
    .ZN(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1996_ (.A1(_1261_),
    .A2(_0421_),
    .B(_0423_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1997_ (.A1(net221),
    .A2(_0418_),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1998_ (.A1(_1263_),
    .A2(_0421_),
    .B(_0424_),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1999_ (.A1(_0388_),
    .A2(_0398_),
    .ZN(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2000_ (.A1(_1253_),
    .A2(_0421_),
    .B(_0425_),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2001_ (.A1(_0390_),
    .A2(_0398_),
    .ZN(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2002_ (.A1(_1252_),
    .A2(_0405_),
    .B(_0426_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2003_ (.A1(_0347_),
    .A2(_0395_),
    .A3(_0351_),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2004_ (.I(_0427_),
    .Z(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2005_ (.I0(\u1.ccr1[16] ),
    .I1(_0392_),
    .S(_0428_),
    .Z(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2006_ (.I(_0429_),
    .Z(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2007_ (.I0(\u1.ccr1[17] ),
    .I1(_0400_),
    .S(_0428_),
    .Z(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2008_ (.I(_0430_),
    .Z(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2009_ (.I(_0427_),
    .Z(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2010_ (.I(_0431_),
    .Z(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2011_ (.I0(\u1.ccr1[18] ),
    .I1(_0361_),
    .S(_0432_),
    .Z(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2012_ (.I(_0433_),
    .Z(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2013_ (.I(\u1.ccr1[19] ),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2014_ (.I(_0431_),
    .Z(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2015_ (.I(_0427_),
    .Z(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2016_ (.A1(_0407_),
    .A2(_0436_),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2017_ (.A1(_0434_),
    .A2(_0435_),
    .B(_0437_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2018_ (.I0(\u1.ccr1[20] ),
    .I1(_0366_),
    .S(_0432_),
    .Z(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2019_ (.I(_0438_),
    .Z(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2020_ (.I0(\u1.ccr1[21] ),
    .I1(_0368_),
    .S(_0432_),
    .Z(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2021_ (.I(_0439_),
    .Z(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2022_ (.A1(_0370_),
    .A2(_0436_),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2023_ (.A1(_1226_),
    .A2(_0435_),
    .B(_0440_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2024_ (.A1(_0373_),
    .A2(_0436_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2025_ (.A1(_1225_),
    .A2(_0435_),
    .B(_0441_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2026_ (.I0(\u1.ccr1[24] ),
    .I1(_0375_),
    .S(_0432_),
    .Z(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2027_ (.I(_0442_),
    .Z(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2028_ (.I(_0431_),
    .Z(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2029_ (.I0(\u1.ccr1[25] ),
    .I1(_0377_),
    .S(_0443_),
    .Z(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2030_ (.I(_0444_),
    .Z(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2031_ (.A1(_0380_),
    .A2(_0428_),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2032_ (.A1(_1178_),
    .A2(_0435_),
    .B(_0445_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2033_ (.A1(_0382_),
    .A2(_0428_),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2034_ (.A1(_1176_),
    .A2(_0436_),
    .B(_0446_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2035_ (.I(net222),
    .Z(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2036_ (.I0(\u1.ccr1[28] ),
    .I1(_0447_),
    .S(_0443_),
    .Z(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2037_ (.I(_0448_),
    .Z(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2038_ (.I0(\u1.ccr1[29] ),
    .I1(_0386_),
    .S(_0443_),
    .Z(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2039_ (.I(_0449_),
    .Z(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2040_ (.I0(\u1.ccr1[30] ),
    .I1(_0388_),
    .S(_0443_),
    .Z(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2041_ (.I(_0450_),
    .Z(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2042_ (.I0(\u1.ccr1[31] ),
    .I1(_0390_),
    .S(_0431_),
    .Z(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2043_ (.I(_0451_),
    .Z(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2044_ (.A1(\u0.cmd[16] ),
    .A2(_0394_),
    .ZN(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2045_ (.A1(\u0.cmd[18] ),
    .A2(_0349_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2046_ (.A1(\u0.write_config_n ),
    .A2(\u0.cmd[21] ),
    .A3(\u0.cmd[20] ),
    .A4(_0453_),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2047_ (.A1(_0452_),
    .A2(_0454_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2048_ (.I(_0455_),
    .Z(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2049_ (.I(_0456_),
    .Z(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2050_ (.I(_0456_),
    .Z(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2051_ (.A1(_0345_),
    .A2(_0458_),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2052_ (.A1(_1133_),
    .A2(_0457_),
    .B(_0459_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2053_ (.A1(_0356_),
    .A2(_0458_),
    .ZN(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2054_ (.A1(_1134_),
    .A2(_0457_),
    .B(_0460_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2055_ (.I(_0404_),
    .Z(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2056_ (.I(_0455_),
    .Z(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2057_ (.I0(_0461_),
    .I1(\u1.ordering_complete[2] ),
    .S(_0462_),
    .Z(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2058_ (.I(_0463_),
    .Z(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2059_ (.I(_0407_),
    .Z(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2060_ (.I0(_0464_),
    .I1(\u1.ordering_complete[3] ),
    .S(_0462_),
    .Z(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2061_ (.I(_0465_),
    .Z(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2062_ (.I(_0409_),
    .Z(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2063_ (.I0(_0466_),
    .I1(\u1.ordering_complete[4] ),
    .S(_0462_),
    .Z(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2064_ (.I(_0467_),
    .Z(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2065_ (.I(_0411_),
    .Z(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2066_ (.I0(_0468_),
    .I1(\u1.ordering_complete[5] ),
    .S(_0462_),
    .Z(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2067_ (.I(_0469_),
    .Z(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2068_ (.I(\u0.cmd[6] ),
    .Z(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2069_ (.I(_0470_),
    .Z(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2070_ (.I(_0455_),
    .Z(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2071_ (.I0(_0471_),
    .I1(\u1.ordering_complete[6] ),
    .S(_0472_),
    .Z(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2072_ (.I(_0473_),
    .Z(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2073_ (.I(\u0.cmd[7] ),
    .Z(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2074_ (.I0(_0474_),
    .I1(\u1.ordering_complete[7] ),
    .S(_0472_),
    .Z(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2075_ (.I(_0475_),
    .Z(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2076_ (.I(\u0.cmd[8] ),
    .Z(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2077_ (.I0(_0476_),
    .I1(_1112_),
    .S(_0472_),
    .Z(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2078_ (.I(_0477_),
    .Z(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2079_ (.I(\u0.cmd[9] ),
    .Z(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2080_ (.I0(_0478_),
    .I1(_1110_),
    .S(_0472_),
    .Z(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2081_ (.I(_0479_),
    .Z(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2082_ (.I(_0455_),
    .Z(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2083_ (.A1(net224),
    .A2(_0480_),
    .ZN(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2084_ (.A1(_1113_),
    .A2(_0457_),
    .B(_0481_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2085_ (.A1(net223),
    .A2(_0480_),
    .ZN(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2086_ (.A1(_1104_),
    .A2(_0457_),
    .B(_0482_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2087_ (.I0(_0447_),
    .I1(\u1.ordering_complete[12] ),
    .S(_0456_),
    .Z(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2088_ (.I(_0483_),
    .Z(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2089_ (.I0(_0386_),
    .I1(\u1.ordering_complete[13] ),
    .S(_0456_),
    .Z(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2090_ (.I(_0484_),
    .Z(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2091_ (.A1(net220),
    .A2(_0480_),
    .ZN(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2092_ (.A1(_1098_),
    .A2(_0458_),
    .B(_0485_),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2093_ (.A1(net219),
    .A2(_0480_),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2094_ (.A1(_1097_),
    .A2(_0458_),
    .B(_0486_),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2095_ (.A1(_0347_),
    .A2(_0394_),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2096_ (.A1(_0487_),
    .A2(_0454_),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2097_ (.I(_0488_),
    .Z(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2098_ (.I(_0489_),
    .Z(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2099_ (.I(_0488_),
    .Z(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2100_ (.I(_0491_),
    .Z(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2101_ (.A1(_0345_),
    .A2(_0492_),
    .ZN(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2102_ (.A1(_1060_),
    .A2(_0490_),
    .B(_0493_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2103_ (.A1(_0356_),
    .A2(_0492_),
    .ZN(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2104_ (.A1(_1061_),
    .A2(_0490_),
    .B(_0494_),
    .ZN(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2105_ (.I(_0491_),
    .Z(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2106_ (.A1(_0404_),
    .A2(_0495_),
    .ZN(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2107_ (.A1(_1067_),
    .A2(_0490_),
    .B(_0496_),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2108_ (.A1(_0407_),
    .A2(_0495_),
    .ZN(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2109_ (.A1(_1058_),
    .A2(_0490_),
    .B(_0497_),
    .ZN(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2110_ (.I(_0491_),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2111_ (.I0(_0466_),
    .I1(\u1.ordering_complete[20] ),
    .S(_0498_),
    .Z(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2112_ (.I(_0499_),
    .Z(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2113_ (.I0(_0468_),
    .I1(\u1.ordering_complete[21] ),
    .S(_0498_),
    .Z(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2114_ (.I(_0500_),
    .Z(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2115_ (.I0(_0471_),
    .I1(\u1.ordering_complete[22] ),
    .S(_0498_),
    .Z(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2116_ (.I(_0501_),
    .Z(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2117_ (.I(_0489_),
    .Z(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2118_ (.A1(\u0.cmd[7] ),
    .A2(_0495_),
    .ZN(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2119_ (.A1(_1054_),
    .A2(_0502_),
    .B(_0503_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2120_ (.I0(_0476_),
    .I1(\u1.ordering_complete[24] ),
    .S(_0498_),
    .Z(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2121_ (.I(_0504_),
    .Z(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2122_ (.I0(_0478_),
    .I1(\u1.ordering_complete[25] ),
    .S(_0489_),
    .Z(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2123_ (.I(_0505_),
    .Z(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2124_ (.I(\u1.ordering_complete[26] ),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2125_ (.A1(\u0.cmd[10] ),
    .A2(_0495_),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2126_ (.A1(_0506_),
    .A2(_0502_),
    .B(_0507_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2127_ (.I(\u1.ordering_complete[27] ),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2128_ (.I(_0491_),
    .Z(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2129_ (.A1(\u0.cmd[11] ),
    .A2(_0509_),
    .ZN(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2130_ (.A1(_0508_),
    .A2(_0502_),
    .B(_0510_),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2131_ (.I0(_0447_),
    .I1(\u1.ordering_complete[28] ),
    .S(_0489_),
    .Z(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2132_ (.I(_0511_),
    .Z(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2133_ (.A1(\u0.cmd[13] ),
    .A2(_0509_),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2134_ (.A1(_1079_),
    .A2(_0502_),
    .B(_0512_),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2135_ (.A1(\u0.cmd[14] ),
    .A2(_0509_),
    .ZN(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2136_ (.A1(_1078_),
    .A2(_0492_),
    .B(_0513_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2137_ (.A1(\u0.cmd[15] ),
    .A2(_0509_),
    .ZN(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2138_ (.A1(_1073_),
    .A2(_0492_),
    .B(_0514_),
    .ZN(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2139_ (.A1(_0347_),
    .A2(_0348_),
    .A3(_0454_),
    .ZN(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2140_ (.I(_0515_),
    .Z(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2141_ (.I0(_0346_),
    .I1(\u1.row_limit[0] ),
    .S(_0516_),
    .Z(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2142_ (.I(_0517_),
    .Z(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2143_ (.I0(_0357_),
    .I1(\u1.row_limit[1] ),
    .S(_0516_),
    .Z(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2144_ (.I(_0518_),
    .Z(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2145_ (.I0(_0461_),
    .I1(\u1.row_limit[2] ),
    .S(_0515_),
    .Z(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2146_ (.I(_0519_),
    .Z(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2147_ (.I0(_0464_),
    .I1(\u1.row_limit[3] ),
    .S(_0515_),
    .Z(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2148_ (.I(_0520_),
    .Z(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2149_ (.I(\u1.row_limit[4] ),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2150_ (.I(_0515_),
    .Z(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2151_ (.A1(_0409_),
    .A2(_0522_),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2152_ (.A1(_0521_),
    .A2(_0522_),
    .B(_0523_),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2153_ (.I(\u1.row_limit[5] ),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2154_ (.A1(_0411_),
    .A2(_0516_),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2155_ (.A1(_0524_),
    .A2(_0522_),
    .B(_0525_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2156_ (.I(\u1.row_limit[6] ),
    .ZN(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2157_ (.A1(_0470_),
    .A2(_0516_),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2158_ (.A1(_0526_),
    .A2(_0522_),
    .B(_0527_),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2159_ (.A1(_0393_),
    .A2(_0348_),
    .A3(_0454_),
    .ZN(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2160_ (.I(_0528_),
    .Z(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2161_ (.I(_0529_),
    .Z(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2162_ (.I(_0528_),
    .Z(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2163_ (.A1(_0345_),
    .A2(_0531_),
    .ZN(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2164_ (.A1(_0321_),
    .A2(_0530_),
    .B(_0532_),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2165_ (.A1(_0356_),
    .A2(_0531_),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2166_ (.A1(_0318_),
    .A2(_0530_),
    .B(_0533_),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2167_ (.A1(_0404_),
    .A2(_0531_),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2168_ (.A1(_0319_),
    .A2(_0530_),
    .B(_0534_),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2169_ (.I0(_0464_),
    .I1(\u1.col_limit[3] ),
    .S(_0529_),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2170_ (.I(_0535_),
    .Z(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2171_ (.I0(_0466_),
    .I1(\u1.col_limit[4] ),
    .S(_0529_),
    .Z(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2172_ (.I(_0536_),
    .Z(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2173_ (.I0(_0468_),
    .I1(\u1.col_limit[5] ),
    .S(_0529_),
    .Z(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2174_ (.I(_0537_),
    .Z(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2175_ (.A1(_0470_),
    .A2(_0531_),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2176_ (.A1(_0310_),
    .A2(_0530_),
    .B(_0538_),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _2177_ (.A1(net218),
    .A2(_0350_),
    .A3(_0452_),
    .ZN(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2178_ (.I(_0539_),
    .Z(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2179_ (.I0(_0346_),
    .I1(\u1.inverter_select[0] ),
    .S(_0540_),
    .Z(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2180_ (.I(_0541_),
    .Z(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2181_ (.I0(_0357_),
    .I1(\u1.inverter_select[1] ),
    .S(_0540_),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2182_ (.I(_0542_),
    .Z(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2183_ (.I0(_0461_),
    .I1(\u1.inverter_select[2] ),
    .S(_0540_),
    .Z(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2184_ (.I(_0543_),
    .Z(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2185_ (.I0(_0464_),
    .I1(\u1.inverter_select[3] ),
    .S(_0540_),
    .Z(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2186_ (.I(_0544_),
    .Z(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2187_ (.I(_0539_),
    .Z(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2188_ (.I0(_0466_),
    .I1(\u1.inverter_select[4] ),
    .S(_0545_),
    .Z(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2189_ (.I(_0546_),
    .Z(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2190_ (.I0(_0468_),
    .I1(\u1.inverter_select[5] ),
    .S(_0545_),
    .Z(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2191_ (.I(_0547_),
    .Z(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2192_ (.I0(_0471_),
    .I1(\u1.inverter_select[6] ),
    .S(_0545_),
    .Z(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2193_ (.I(_0548_),
    .Z(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2194_ (.I0(_0474_),
    .I1(\u1.inverter_select[7] ),
    .S(_0545_),
    .Z(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2195_ (.I(_0549_),
    .Z(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2196_ (.I0(_0476_),
    .I1(\u1.inverter_select[8] ),
    .S(_0539_),
    .Z(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2197_ (.I(_0550_),
    .Z(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2198_ (.I0(_0478_),
    .I1(\u1.inverter_select[9] ),
    .S(_0539_),
    .Z(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2199_ (.I(_0551_),
    .Z(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _2200_ (.A1(\u0.cmd[19] ),
    .A2(_0487_),
    .A3(_0350_),
    .ZN(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2201_ (.I(_0552_),
    .Z(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2202_ (.I0(_0346_),
    .I1(\u1.row_col_select[0] ),
    .S(_0553_),
    .Z(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2203_ (.I(_0554_),
    .Z(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2204_ (.I0(_0357_),
    .I1(\u1.row_col_select[1] ),
    .S(_0553_),
    .Z(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2205_ (.I(_0555_),
    .Z(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2206_ (.I0(_0461_),
    .I1(\u1.row_col_select[2] ),
    .S(_0553_),
    .Z(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2207_ (.I(_0556_),
    .Z(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2208_ (.I0(_0364_),
    .I1(\u1.row_col_select[3] ),
    .S(_0553_),
    .Z(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2209_ (.I(_0557_),
    .Z(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2210_ (.I(_0552_),
    .Z(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2211_ (.I0(_0366_),
    .I1(\u1.row_col_select[4] ),
    .S(_0558_),
    .Z(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2212_ (.I(_0559_),
    .Z(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2213_ (.I0(_0368_),
    .I1(\u1.row_col_select[5] ),
    .S(_0558_),
    .Z(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2214_ (.I(_0560_),
    .Z(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2215_ (.I0(_0471_),
    .I1(\u1.row_col_select[6] ),
    .S(_0558_),
    .Z(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2216_ (.I(_0561_),
    .Z(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2217_ (.I0(_0474_),
    .I1(\u1.row_col_select[7] ),
    .S(_0558_),
    .Z(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2218_ (.I(_0562_),
    .Z(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2219_ (.I0(_0476_),
    .I1(\u1.row_col_select[8] ),
    .S(_0552_),
    .Z(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2220_ (.I(_0563_),
    .Z(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2221_ (.I0(_0478_),
    .I1(\u1.row_col_select[9] ),
    .S(_0552_),
    .Z(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2222_ (.I(_0564_),
    .Z(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2223_ (.I(_1402_),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2224_ (.A1(_1070_),
    .A2(_1095_),
    .ZN(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2225_ (.A1(_1135_),
    .A2(_1140_),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2226_ (.A1(_1141_),
    .A2(_0567_),
    .B(_1137_),
    .ZN(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2227_ (.A1(_1123_),
    .A2(_1131_),
    .B(_1126_),
    .ZN(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2228_ (.A1(_1132_),
    .A2(_0568_),
    .B1(_0569_),
    .B2(_1129_),
    .ZN(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2229_ (.I(_1096_),
    .ZN(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2230_ (.A1(_1102_),
    .A2(_1106_),
    .ZN(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2231_ (.A1(_0571_),
    .A2(\u1.ordering_complete[15] ),
    .B1(_1099_),
    .B2(_0572_),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2232_ (.A1(_1109_),
    .A2(_1110_),
    .B1(_1111_),
    .B2(\u1.ordering_complete[8] ),
    .ZN(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2233_ (.A1(_1117_),
    .A2(_0574_),
    .ZN(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2234_ (.A1(_1114_),
    .A2(_0575_),
    .B(_1108_),
    .ZN(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2235_ (.A1(_1120_),
    .A2(_0570_),
    .B(_0573_),
    .C(_0576_),
    .ZN(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2236_ (.A1(_0566_),
    .A2(_0577_),
    .Z(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2237_ (.A1(_1187_),
    .A2(_1235_),
    .A3(_1245_),
    .ZN(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2238_ (.A1(_1205_),
    .A2(_1216_),
    .A3(_1217_),
    .A4(_1220_),
    .Z(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2239_ (.A1(_1210_),
    .A2(_0580_),
    .ZN(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _2240_ (.A1(_1202_),
    .A2(_1277_),
    .A3(_0579_),
    .A4(_0581_),
    .ZN(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2241_ (.I(\u1.ordering_timer[19] ),
    .Z(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2242_ (.A1(_0583_),
    .A2(_1058_),
    .ZN(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2243_ (.A1(_1062_),
    .A2(_1069_),
    .ZN(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2244_ (.A1(_1066_),
    .A2(_0585_),
    .ZN(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2245_ (.A1(_1051_),
    .A2(_1053_),
    .B(_1048_),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2246_ (.A1(_1057_),
    .A2(_0584_),
    .A3(_0586_),
    .B1(_0587_),
    .B2(_1055_),
    .ZN(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2247_ (.A1(\u1.ordering_timer[27] ),
    .A2(_0508_),
    .B1(\u1.ordering_timer[26] ),
    .B2(_0506_),
    .C1(_1089_),
    .C2(_1092_),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2248_ (.A1(_1084_),
    .A2(_0589_),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2249_ (.I(_1080_),
    .ZN(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2250_ (.A1(_1077_),
    .A2(_0591_),
    .ZN(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2251_ (.A1(_1083_),
    .A2(_0592_),
    .B(_1074_),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2252_ (.A1(_1095_),
    .A2(_0588_),
    .B(_0590_),
    .C(_0593_),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2253_ (.A1(_1212_),
    .A2(_0578_),
    .A3(_0582_),
    .A4(_0594_),
    .Z(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2254_ (.I(_0595_),
    .Z(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2255_ (.I(_0596_),
    .Z(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2256_ (.A1(_1139_),
    .A2(_0597_),
    .Z(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2257_ (.A1(_0565_),
    .A2(_0598_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2258_ (.I(\u1.ordering_timer[1] ),
    .Z(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2259_ (.A1(_1403_),
    .A2(_0595_),
    .ZN(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2260_ (.I(_0600_),
    .Z(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2261_ (.I(_0601_),
    .Z(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2262_ (.A1(_0565_),
    .A2(_0600_),
    .ZN(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2263_ (.I(_0603_),
    .Z(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2264_ (.I(_0604_),
    .Z(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2265_ (.A1(_1138_),
    .A2(_0599_),
    .Z(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2266_ (.I(_0595_),
    .Z(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2267_ (.I(_0607_),
    .Z(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2268_ (.I(_0608_),
    .Z(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2269_ (.I0(\u1.ordering_complete[1] ),
    .I1(_0606_),
    .S(_0609_),
    .Z(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2270_ (.A1(_0599_),
    .A2(_0602_),
    .B1(_0605_),
    .B2(_0610_),
    .ZN(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2271_ (.I(_0611_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2272_ (.I(_0607_),
    .Z(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2273_ (.I(_0612_),
    .Z(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2274_ (.A1(_1138_),
    .A2(_0599_),
    .A3(\u1.ordering_timer[2] ),
    .ZN(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2275_ (.A1(_1138_),
    .A2(_0599_),
    .ZN(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2276_ (.A1(_1136_),
    .A2(_0615_),
    .ZN(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2277_ (.A1(_0614_),
    .A2(_0616_),
    .ZN(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2278_ (.A1(\u1.ordering_complete[2] ),
    .A2(_0597_),
    .ZN(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2279_ (.A1(_0613_),
    .A2(_0617_),
    .B(_0618_),
    .ZN(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2280_ (.A1(\u1.ordering_timer[2] ),
    .A2(_0602_),
    .B1(_0605_),
    .B2(_0619_),
    .ZN(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2281_ (.I(_0620_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2282_ (.A1(\u1.ordering_timer[3] ),
    .A2(_0614_),
    .Z(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2283_ (.A1(\u1.ordering_complete[3] ),
    .A2(_0597_),
    .ZN(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2284_ (.A1(_0613_),
    .A2(_0621_),
    .B(_0622_),
    .ZN(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2285_ (.A1(\u1.ordering_timer[3] ),
    .A2(_0602_),
    .B1(_0605_),
    .B2(_0623_),
    .ZN(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2286_ (.I(_0624_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2287_ (.I(\u1.ordering_timer[4] ),
    .Z(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2288_ (.I(_0600_),
    .Z(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2289_ (.I(_0626_),
    .Z(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2290_ (.A1(\u1.ordering_timer[0] ),
    .A2(\u1.ordering_timer[1] ),
    .A3(\u1.ordering_timer[3] ),
    .A4(\u1.ordering_timer[2] ),
    .Z(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2291_ (.A1(_1122_),
    .A2(_0628_),
    .Z(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2292_ (.I(_0608_),
    .Z(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2293_ (.A1(\u1.ordering_complete[4] ),
    .A2(_0630_),
    .ZN(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2294_ (.A1(_0613_),
    .A2(_0629_),
    .B(_0631_),
    .ZN(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2295_ (.A1(_0625_),
    .A2(_0627_),
    .B1(_0605_),
    .B2(_0632_),
    .ZN(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2296_ (.I(_0633_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2297_ (.I(_0603_),
    .Z(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2298_ (.I(_0634_),
    .Z(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2299_ (.A1(\u1.ordering_timer[5] ),
    .A2(_0625_),
    .A3(_0628_),
    .ZN(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2300_ (.A1(_0625_),
    .A2(_0628_),
    .ZN(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2301_ (.A1(_1121_),
    .A2(_0637_),
    .ZN(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2302_ (.A1(_0636_),
    .A2(_0638_),
    .ZN(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2303_ (.A1(\u1.ordering_complete[5] ),
    .A2(_0630_),
    .ZN(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2304_ (.A1(_0613_),
    .A2(_0639_),
    .B(_0640_),
    .ZN(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2305_ (.A1(\u1.ordering_timer[5] ),
    .A2(_0627_),
    .B1(_0635_),
    .B2(_0641_),
    .ZN(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2306_ (.I(_0642_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2307_ (.I(_0612_),
    .Z(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2308_ (.A1(\u1.ordering_timer[6] ),
    .A2(_0636_),
    .Z(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2309_ (.A1(\u1.ordering_complete[6] ),
    .A2(_0630_),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2310_ (.A1(_0643_),
    .A2(_0644_),
    .B(_0645_),
    .ZN(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2311_ (.A1(\u1.ordering_timer[6] ),
    .A2(_0627_),
    .B1(_0635_),
    .B2(_0646_),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2312_ (.I(_0647_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2313_ (.I(\u1.ordering_timer[7] ),
    .Z(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2314_ (.A1(\u1.ordering_timer[6] ),
    .A2(\u1.ordering_timer[5] ),
    .A3(_0625_),
    .A4(_0628_),
    .Z(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2315_ (.A1(_1124_),
    .A2(_0649_),
    .Z(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2316_ (.A1(\u1.ordering_complete[7] ),
    .A2(_0630_),
    .ZN(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2317_ (.A1(_0643_),
    .A2(_0650_),
    .B(_0651_),
    .ZN(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2318_ (.A1(_0648_),
    .A2(_0627_),
    .B1(_0635_),
    .B2(_0652_),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2319_ (.I(_0653_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2320_ (.I(\u1.ordering_timer[8] ),
    .Z(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2321_ (.I(_0626_),
    .Z(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2322_ (.A1(_0648_),
    .A2(_0649_),
    .Z(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2323_ (.A1(_1111_),
    .A2(_0656_),
    .Z(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2324_ (.I(_0596_),
    .Z(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2325_ (.A1(_1112_),
    .A2(_0658_),
    .ZN(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2326_ (.A1(_0643_),
    .A2(_0657_),
    .B(_0659_),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2327_ (.A1(_0654_),
    .A2(_0655_),
    .B1(_0635_),
    .B2(_0660_),
    .ZN(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2328_ (.I(_0661_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2329_ (.I(_0634_),
    .Z(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2330_ (.A1(_0654_),
    .A2(_0656_),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2331_ (.A1(_1109_),
    .A2(_0663_),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2332_ (.A1(_0648_),
    .A2(\u1.ordering_timer[9] ),
    .A3(_0654_),
    .A4(_0649_),
    .ZN(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2333_ (.A1(_0664_),
    .A2(_0665_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2334_ (.A1(_1110_),
    .A2(_0658_),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2335_ (.A1(_0643_),
    .A2(_0666_),
    .B(_0667_),
    .ZN(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2336_ (.A1(\u1.ordering_timer[9] ),
    .A2(_0655_),
    .B1(_0662_),
    .B2(_0668_),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2337_ (.I(_0669_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2338_ (.I(_0612_),
    .Z(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2339_ (.A1(\u1.ordering_timer[10] ),
    .A2(_0665_),
    .Z(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2340_ (.A1(\u1.ordering_complete[10] ),
    .A2(_0658_),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2341_ (.A1(_0670_),
    .A2(_0671_),
    .B(_0672_),
    .ZN(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2342_ (.A1(\u1.ordering_timer[10] ),
    .A2(_0655_),
    .B1(_0662_),
    .B2(_0673_),
    .ZN(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2343_ (.I(_0674_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2344_ (.I(\u1.ordering_timer[11] ),
    .Z(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2345_ (.I(_0675_),
    .ZN(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2346_ (.A1(_1116_),
    .A2(_0665_),
    .ZN(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2347_ (.A1(_0676_),
    .A2(_0677_),
    .Z(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2348_ (.A1(\u1.ordering_complete[11] ),
    .A2(_0658_),
    .ZN(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2349_ (.A1(_0670_),
    .A2(_0678_),
    .B(_0679_),
    .ZN(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2350_ (.A1(_0675_),
    .A2(_0655_),
    .B1(_0662_),
    .B2(_0680_),
    .ZN(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2351_ (.I(_0681_),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2352_ (.I(_0626_),
    .Z(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2353_ (.A1(_0675_),
    .A2(_0677_),
    .ZN(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2354_ (.A1(_1103_),
    .A2(_0683_),
    .ZN(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2355_ (.A1(\u1.ordering_timer[12] ),
    .A2(_0675_),
    .A3(_0677_),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2356_ (.A1(_0684_),
    .A2(_0685_),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2357_ (.I(_0596_),
    .Z(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2358_ (.A1(\u1.ordering_complete[12] ),
    .A2(_0687_),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2359_ (.A1(_0670_),
    .A2(_0686_),
    .B(_0688_),
    .ZN(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2360_ (.A1(\u1.ordering_timer[12] ),
    .A2(_0682_),
    .B1(_0662_),
    .B2(_0689_),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2361_ (.I(_0690_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2362_ (.I(_0634_),
    .Z(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2363_ (.A1(\u1.ordering_timer[13] ),
    .A2(\u1.ordering_timer[12] ),
    .ZN(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _2364_ (.A1(_0676_),
    .A2(_1116_),
    .A3(_0665_),
    .A4(_0692_),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2365_ (.I(_0693_),
    .Z(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2366_ (.A1(_1101_),
    .A2(_0685_),
    .B(_0694_),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2367_ (.I0(\u1.ordering_complete[13] ),
    .I1(_0695_),
    .S(_0609_),
    .Z(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2368_ (.A1(\u1.ordering_timer[13] ),
    .A2(_0682_),
    .B1(_0691_),
    .B2(_0696_),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2369_ (.I(_0697_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2370_ (.I(\u1.ordering_timer[14] ),
    .Z(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2371_ (.A1(_1100_),
    .A2(_0694_),
    .Z(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2372_ (.A1(\u1.ordering_complete[14] ),
    .A2(_0687_),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2373_ (.A1(_0670_),
    .A2(_0699_),
    .B(_0700_),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2374_ (.A1(_0698_),
    .A2(_0682_),
    .B1(_0691_),
    .B2(_0701_),
    .ZN(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2375_ (.I(_0702_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2376_ (.I(_1096_),
    .Z(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2377_ (.A1(_0698_),
    .A2(_0694_),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2378_ (.A1(_0703_),
    .A2(_0704_),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2379_ (.I0(\u1.ordering_complete[15] ),
    .I1(_0705_),
    .S(_0609_),
    .Z(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2380_ (.A1(_0703_),
    .A2(_0682_),
    .B1(_0691_),
    .B2(_0706_),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2381_ (.I(_0707_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2382_ (.I(_1059_),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2383_ (.I(_0601_),
    .ZN(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2384_ (.I(_0709_),
    .Z(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2385_ (.I(_0608_),
    .Z(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2386_ (.A1(_0703_),
    .A2(_0698_),
    .A3(_0694_),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2387_ (.A1(_1059_),
    .A2(_0712_),
    .Z(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2388_ (.I(_0607_),
    .Z(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2389_ (.A1(\u1.ordering_complete[16] ),
    .A2(_0714_),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2390_ (.I(_0601_),
    .Z(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2391_ (.A1(_0711_),
    .A2(_0713_),
    .B(_0715_),
    .C(_0716_),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2392_ (.A1(_0329_),
    .A2(_0717_),
    .ZN(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2393_ (.A1(_0708_),
    .A2(_0710_),
    .B(_0718_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2394_ (.I(_0626_),
    .Z(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2395_ (.I(_0612_),
    .Z(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2396_ (.A1(_0708_),
    .A2(_0712_),
    .ZN(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2397_ (.A1(_1068_),
    .A2(_1059_),
    .Z(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2398_ (.A1(_1096_),
    .A2(\u1.ordering_timer[14] ),
    .A3(_0693_),
    .A4(_0722_),
    .Z(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2399_ (.I(_0723_),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2400_ (.A1(_1068_),
    .A2(_0721_),
    .B(_0724_),
    .C(_0714_),
    .ZN(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2401_ (.A1(_1061_),
    .A2(_0720_),
    .B(_0725_),
    .ZN(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2402_ (.A1(_1068_),
    .A2(_0719_),
    .B1(_0691_),
    .B2(_0726_),
    .ZN(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2403_ (.I(_0727_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2404_ (.I(_1065_),
    .Z(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2405_ (.A1(_0728_),
    .A2(_0723_),
    .Z(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2406_ (.A1(\u1.ordering_complete[18] ),
    .A2(_0714_),
    .ZN(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2407_ (.A1(_0711_),
    .A2(_0729_),
    .B(_0730_),
    .C(_0716_),
    .ZN(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2408_ (.A1(_0329_),
    .A2(_0731_),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2409_ (.A1(_0728_),
    .A2(_0710_),
    .B(_0732_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2410_ (.I(_0634_),
    .Z(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2411_ (.I(_0608_),
    .Z(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2412_ (.A1(\u1.ordering_timer[18] ),
    .A2(_0723_),
    .B(_0583_),
    .ZN(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2413_ (.A1(_1064_),
    .A2(_0728_),
    .A3(_0724_),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2414_ (.A1(_0735_),
    .A2(_0736_),
    .Z(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2415_ (.A1(\u1.ordering_complete[19] ),
    .A2(_0687_),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2416_ (.A1(_0734_),
    .A2(_0737_),
    .B(_0738_),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2417_ (.A1(_0583_),
    .A2(_0719_),
    .B1(_0733_),
    .B2(_0739_),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2418_ (.I(_0740_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2419_ (.A1(_1050_),
    .A2(_0736_),
    .Z(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2420_ (.A1(\u1.ordering_complete[20] ),
    .A2(_0687_),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2421_ (.A1(_0734_),
    .A2(_0741_),
    .B(_0742_),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2422_ (.A1(\u1.ordering_timer[20] ),
    .A2(_0719_),
    .B1(_0733_),
    .B2(_0743_),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2423_ (.I(_0744_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2424_ (.A1(\u1.ordering_timer[20] ),
    .A2(_0736_),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2425_ (.A1(\u1.ordering_timer[21] ),
    .A2(\u1.ordering_timer[20] ),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2426_ (.I(_0746_),
    .ZN(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2427_ (.A1(_0583_),
    .A2(\u1.ordering_timer[18] ),
    .A3(_0723_),
    .A4(_0747_),
    .Z(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2428_ (.I(_0748_),
    .Z(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2429_ (.A1(_1049_),
    .A2(_0745_),
    .B(_0749_),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2430_ (.I0(\u1.ordering_complete[21] ),
    .I1(_0750_),
    .S(_0609_),
    .Z(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2431_ (.A1(\u1.ordering_timer[21] ),
    .A2(_0719_),
    .B1(_0733_),
    .B2(_0751_),
    .ZN(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2432_ (.I(_0752_),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2433_ (.I(\u1.ordering_timer[22] ),
    .Z(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2434_ (.I(_0601_),
    .Z(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2435_ (.A1(_1047_),
    .A2(_0749_),
    .Z(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2436_ (.I(_0596_),
    .Z(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2437_ (.A1(\u1.ordering_complete[22] ),
    .A2(_0756_),
    .ZN(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2438_ (.A1(_0734_),
    .A2(_0755_),
    .B(_0757_),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2439_ (.A1(_0753_),
    .A2(_0754_),
    .B1(_0733_),
    .B2(_0758_),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2440_ (.I(_0759_),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2441_ (.I(\u1.ordering_timer[23] ),
    .Z(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2442_ (.I(_0603_),
    .Z(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2443_ (.A1(_0753_),
    .A2(_0749_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2444_ (.A1(_1046_),
    .A2(_0762_),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2445_ (.A1(_0760_),
    .A2(_0753_),
    .A3(_0749_),
    .ZN(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2446_ (.A1(_0756_),
    .A2(_0763_),
    .A3(_0764_),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2447_ (.A1(_1054_),
    .A2(_0720_),
    .B(_0765_),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2448_ (.A1(_0760_),
    .A2(_0754_),
    .B1(_0761_),
    .B2(_0766_),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2449_ (.I(_0767_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2450_ (.I(_1085_),
    .Z(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2451_ (.A1(_0768_),
    .A2(_0764_),
    .Z(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2452_ (.A1(\u1.ordering_complete[24] ),
    .A2(_0756_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2453_ (.A1(_0734_),
    .A2(_0769_),
    .B(_0770_),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2454_ (.A1(_0768_),
    .A2(_0754_),
    .B1(_0761_),
    .B2(_0771_),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2455_ (.I(_0772_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2456_ (.I(\u1.ordering_timer[25] ),
    .Z(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2457_ (.A1(_0648_),
    .A2(\u1.ordering_timer[9] ),
    .A3(_0654_),
    .A4(_0649_),
    .ZN(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _2458_ (.A1(_0676_),
    .A2(_1116_),
    .A3(_0774_),
    .A4(_0692_),
    .ZN(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2459_ (.A1(_0703_),
    .A2(_0698_),
    .A3(_0775_),
    .A4(_0722_),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _2460_ (.A1(_1064_),
    .A2(_0728_),
    .A3(_0776_),
    .A4(_0746_),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2461_ (.A1(_1085_),
    .A2(_0760_),
    .A3(_0753_),
    .A4(_0777_),
    .Z(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2462_ (.A1(_0773_),
    .A2(_0778_),
    .Z(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2463_ (.I(_0607_),
    .Z(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2464_ (.I0(\u1.ordering_complete[25] ),
    .I1(_0779_),
    .S(_0780_),
    .Z(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2465_ (.A1(_0773_),
    .A2(_0754_),
    .B1(_0761_),
    .B2(_0781_),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2466_ (.I(_0782_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2467_ (.I(\u1.ordering_timer[26] ),
    .Z(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2468_ (.A1(_0773_),
    .A2(_0760_),
    .A3(\u1.ordering_timer[22] ),
    .A4(_0748_),
    .Z(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2469_ (.A1(_0768_),
    .A2(_0784_),
    .Z(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2470_ (.A1(_1087_),
    .A2(_0785_),
    .Z(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2471_ (.A1(\u1.ordering_complete[26] ),
    .A2(_0756_),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2472_ (.A1(_0711_),
    .A2(_0786_),
    .B(_0787_),
    .ZN(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2473_ (.A1(_0783_),
    .A2(_0716_),
    .B1(_0761_),
    .B2(_0788_),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2474_ (.I(_0789_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2475_ (.A1(_0783_),
    .A2(_0773_),
    .A3(_0778_),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2476_ (.A1(\u1.ordering_timer[27] ),
    .A2(_0783_),
    .A3(_1085_),
    .A4(_0784_),
    .Z(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2477_ (.I(_0780_),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2478_ (.A1(_1093_),
    .A2(_0790_),
    .B(_0791_),
    .C(_0792_),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2479_ (.A1(_0508_),
    .A2(_0711_),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2480_ (.A1(_0793_),
    .A2(_0794_),
    .B(_0604_),
    .ZN(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2481_ (.A1(_1093_),
    .A2(_0710_),
    .B(_0795_),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2482_ (.I(_1071_),
    .Z(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2483_ (.A1(_0796_),
    .A2(_0791_),
    .Z(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2484_ (.A1(_0597_),
    .A2(_0797_),
    .ZN(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2485_ (.A1(\u1.ordering_complete[28] ),
    .A2(_0720_),
    .B(_0604_),
    .C(_0798_),
    .ZN(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2486_ (.A1(_0796_),
    .A2(_0710_),
    .B(_0799_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2487_ (.A1(\u1.ordering_timer[28] ),
    .A2(_0791_),
    .B(\u1.ordering_timer[29] ),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _2488_ (.A1(_1076_),
    .A2(_0796_),
    .A3(_1093_),
    .A4(_0790_),
    .ZN(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2489_ (.A1(_0800_),
    .A2(_0801_),
    .B(_0714_),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2490_ (.A1(\u1.ordering_complete[29] ),
    .A2(_0720_),
    .B(_0709_),
    .C(_0802_),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2491_ (.A1(_1076_),
    .A2(_0709_),
    .B1(_0803_),
    .B2(_0565_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2492_ (.A1(\u1.ordering_complete[30] ),
    .A2(_0792_),
    .ZN(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2493_ (.A1(_1082_),
    .A2(\u1.ordering_timer[29] ),
    .ZN(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2494_ (.A1(\u1.ordering_timer[28] ),
    .A2(_0791_),
    .ZN(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2495_ (.A1(_1082_),
    .A2(_0801_),
    .B1(_0805_),
    .B2(_0806_),
    .C(_0780_),
    .ZN(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2496_ (.A1(_0804_),
    .A2(_0807_),
    .Z(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2497_ (.A1(_1082_),
    .A2(_0716_),
    .ZN(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2498_ (.A1(_0565_),
    .A2(_0602_),
    .A3(_0808_),
    .B(_0809_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2499_ (.I(\u1.ordering_timer[31] ),
    .ZN(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2500_ (.A1(\u1.ordering_timer[27] ),
    .A2(_0783_),
    .A3(_0768_),
    .A4(_0784_),
    .ZN(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2501_ (.A1(_0796_),
    .A2(_0811_),
    .A3(_0805_),
    .B(_0810_),
    .ZN(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2502_ (.I0(\u1.ordering_complete[31] ),
    .I1(_0812_),
    .S(_0780_),
    .Z(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2503_ (.A1(_0604_),
    .A2(_0813_),
    .ZN(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2504_ (.A1(_0810_),
    .A2(_0709_),
    .B(_0814_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2505_ (.I(_1041_),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2506_ (.A1(_0815_),
    .A2(\u0.latch_cmd ),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2507_ (.I(_0816_),
    .Z(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2508_ (.I(_0817_),
    .Z(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2509_ (.A1(_1042_),
    .A2(\u0.latch_cmd ),
    .Z(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2510_ (.I(_0819_),
    .Z(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2511_ (.I(_0820_),
    .Z(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2512_ (.A1(_0392_),
    .A2(_0818_),
    .B1(_0821_),
    .B2(\spi_data_crossing[0].data_sync ),
    .ZN(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2513_ (.I(_0822_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2514_ (.A1(_0400_),
    .A2(_0818_),
    .B1(_0821_),
    .B2(\spi_data_crossing[1].data_sync ),
    .ZN(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2515_ (.I(_0823_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2516_ (.A1(_0361_),
    .A2(_0818_),
    .B1(_0821_),
    .B2(\spi_data_crossing[2].data_sync ),
    .ZN(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2517_ (.I(_0824_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2518_ (.A1(_0364_),
    .A2(_0818_),
    .B1(_0821_),
    .B2(\spi_data_crossing[3].data_sync ),
    .ZN(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2519_ (.I(_0825_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2520_ (.I(_0817_),
    .Z(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2521_ (.I(_0820_),
    .Z(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2522_ (.A1(_0366_),
    .A2(_0826_),
    .B1(_0827_),
    .B2(\spi_data_crossing[4].data_sync ),
    .ZN(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2523_ (.I(_0828_),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2524_ (.A1(_0368_),
    .A2(_0826_),
    .B1(_0827_),
    .B2(\spi_data_crossing[5].data_sync ),
    .ZN(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2525_ (.I(_0829_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2526_ (.A1(_0370_),
    .A2(_0826_),
    .B1(_0827_),
    .B2(\spi_data_crossing[6].data_sync ),
    .ZN(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2527_ (.I(_0830_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2528_ (.A1(_0474_),
    .A2(_0826_),
    .B1(_0827_),
    .B2(\spi_data_crossing[7].data_sync ),
    .ZN(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2529_ (.I(_0831_),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2530_ (.I(_0817_),
    .Z(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2531_ (.I(_0820_),
    .Z(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2532_ (.A1(_0375_),
    .A2(_0832_),
    .B1(_0833_),
    .B2(\spi_data_crossing[8].data_sync ),
    .ZN(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2533_ (.I(_0834_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2534_ (.A1(_0377_),
    .A2(_0832_),
    .B1(_0833_),
    .B2(\spi_data_crossing[9].data_sync ),
    .ZN(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2535_ (.I(_0835_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2536_ (.A1(_0380_),
    .A2(_0832_),
    .B1(_0833_),
    .B2(\spi_data_crossing[10].data_sync ),
    .ZN(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2537_ (.I(_0836_),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2538_ (.A1(_0382_),
    .A2(_0832_),
    .B1(_0833_),
    .B2(\spi_data_crossing[11].data_sync ),
    .ZN(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2539_ (.I(_0837_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2540_ (.I(_0817_),
    .Z(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2541_ (.I(_0820_),
    .Z(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2542_ (.A1(_0447_),
    .A2(_0838_),
    .B1(_0839_),
    .B2(\spi_data_crossing[12].data_sync ),
    .ZN(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2543_ (.I(_0840_),
    .ZN(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2544_ (.A1(_0386_),
    .A2(_0838_),
    .B1(_0839_),
    .B2(\spi_data_crossing[13].data_sync ),
    .ZN(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2545_ (.I(_0841_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2546_ (.A1(_0388_),
    .A2(_0838_),
    .B1(_0839_),
    .B2(\spi_data_crossing[14].data_sync ),
    .ZN(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2547_ (.I(_0842_),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2548_ (.A1(_0390_),
    .A2(_0838_),
    .B1(_0839_),
    .B2(\spi_data_crossing[15].data_sync ),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2549_ (.I(_0843_),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2550_ (.I(_0816_),
    .Z(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2551_ (.I(_0844_),
    .Z(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2552_ (.I(_0819_),
    .Z(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2553_ (.I(_0846_),
    .Z(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2554_ (.A1(_0393_),
    .A2(_0845_),
    .B1(_0847_),
    .B2(\spi_data_crossing[16].data_sync ),
    .ZN(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2555_ (.I(_0848_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2556_ (.A1(_0348_),
    .A2(_0845_),
    .B1(_0847_),
    .B2(\spi_data_crossing[17].data_sync ),
    .ZN(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2557_ (.I(_0849_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2558_ (.A1(\u0.cmd[18] ),
    .A2(_0845_),
    .B1(_0847_),
    .B2(\spi_data_crossing[18].data_sync ),
    .ZN(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2559_ (.I(_0850_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2560_ (.A1(net218),
    .A2(_0845_),
    .B1(_0847_),
    .B2(\spi_data_crossing[19].data_sync ),
    .ZN(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2561_ (.I(_0851_),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2562_ (.I(_0844_),
    .Z(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2563_ (.I(_0846_),
    .Z(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2564_ (.A1(\u0.cmd[20] ),
    .A2(_0852_),
    .B1(_0853_),
    .B2(\spi_data_crossing[20].data_sync ),
    .ZN(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2565_ (.I(_0854_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2566_ (.A1(\u0.cmd[21] ),
    .A2(_0852_),
    .B1(_0853_),
    .B2(\spi_data_crossing[21].data_sync ),
    .ZN(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2567_ (.I(_0855_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2568_ (.A1(\u0.cmd[22] ),
    .A2(_0852_),
    .B1(_0853_),
    .B2(\spi_data_crossing[22].data_sync ),
    .ZN(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2569_ (.I(_0856_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2570_ (.A1(\u0.cmd[23] ),
    .A2(_0852_),
    .B1(_0853_),
    .B2(\spi_data_crossing[23].data_sync ),
    .ZN(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2571_ (.I(_0857_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2572_ (.I(_0844_),
    .Z(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2573_ (.I(_0846_),
    .Z(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2574_ (.A1(\u0.cmd[24] ),
    .A2(_0858_),
    .B1(_0859_),
    .B2(\spi_data_crossing[24].data_sync ),
    .ZN(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2575_ (.I(_0860_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2576_ (.A1(\u0.cmd[25] ),
    .A2(_0858_),
    .B1(_0859_),
    .B2(\spi_data_crossing[25].data_sync ),
    .ZN(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2577_ (.I(_0861_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2578_ (.A1(_0299_),
    .A2(_0858_),
    .B1(_0859_),
    .B2(\spi_data_crossing[26].data_sync ),
    .ZN(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2579_ (.I(_0862_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2580_ (.A1(_1160_),
    .A2(_0858_),
    .B1(_0859_),
    .B2(\spi_data_crossing[27].data_sync ),
    .ZN(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2581_ (.I(_0863_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2582_ (.I(_0844_),
    .Z(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2583_ (.I(_0846_),
    .Z(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2584_ (.A1(\u0.cmd[28] ),
    .A2(_0864_),
    .B1(_0865_),
    .B2(\spi_data_crossing[28].data_sync ),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2585_ (.I(_0866_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2586_ (.A1(\u0.cmd[29] ),
    .A2(_0864_),
    .B1(_0865_),
    .B2(\spi_data_crossing[29].data_sync ),
    .ZN(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2587_ (.I(_0867_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2588_ (.A1(\u0.cmd[30] ),
    .A2(_0864_),
    .B1(_0865_),
    .B2(\spi_data_crossing[30].data_sync ),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2589_ (.I(_0868_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2590_ (.A1(_1040_),
    .A2(_0864_),
    .B1(_0865_),
    .B2(\spi_data_crossing[31].data_sync ),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2591_ (.I(_0869_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2592_ (.A1(net226),
    .A2(_0321_),
    .ZN(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2593_ (.A1(_0312_),
    .A2(_0324_),
    .A3(_0870_),
    .ZN(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2594_ (.A1(_0322_),
    .A2(_0326_),
    .A3(_0871_),
    .ZN(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2595_ (.A1(_0313_),
    .A2(\u1.col_limit[3] ),
    .B1(_0316_),
    .B2(\u1.col_limit[2] ),
    .C(_0315_),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2596_ (.A1(_0320_),
    .A2(_0872_),
    .A3(_0873_),
    .ZN(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2597_ (.A1(_0309_),
    .A2(_0874_),
    .B(_1212_),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2598_ (.I(net217),
    .ZN(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2599_ (.I(\u1.row_sel[3] ),
    .ZN(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2600_ (.I(\u1.row_sel[1] ),
    .ZN(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2601_ (.I(\u1.row_sel[0] ),
    .ZN(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2602_ (.A1(\u1.row_limit[1] ),
    .A2(_0878_),
    .B(\u1.row_limit[0] ),
    .C(_0879_),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2603_ (.I(\u1.row_sel[2] ),
    .ZN(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2604_ (.A1(\u1.row_limit[2] ),
    .A2(_0881_),
    .B1(\u1.row_limit[1] ),
    .B2(_0878_),
    .ZN(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2605_ (.A1(\u1.row_limit[3] ),
    .A2(_0877_),
    .B1(\u1.row_limit[2] ),
    .B2(_0881_),
    .ZN(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2606_ (.A1(_0880_),
    .A2(_0882_),
    .B(_0883_),
    .ZN(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2607_ (.A1(\u1.row_limit[4] ),
    .A2(_0876_),
    .B1(\u1.row_limit[3] ),
    .B2(_0877_),
    .C(_0884_),
    .ZN(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2608_ (.A1(_0524_),
    .A2(net216),
    .B1(_0521_),
    .B2(net217),
    .C(_0885_),
    .ZN(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2609_ (.A1(\u1.row_sel[6] ),
    .A2(_0526_),
    .B1(_0524_),
    .B2(net216),
    .ZN(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2610_ (.A1(\u1.row_sel[6] ),
    .A2(_0526_),
    .ZN(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2611_ (.A1(_0886_),
    .A2(_0887_),
    .B(_0888_),
    .C(_0329_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2612_ (.A1(_0875_),
    .A2(_0889_),
    .Z(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2613_ (.I(_0890_),
    .Z(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2614_ (.A1(\u1.row_sel[0] ),
    .A2(_0875_),
    .Z(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2615_ (.A1(\u1.row_sel[0] ),
    .A2(_0875_),
    .ZN(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2616_ (.A1(_0891_),
    .A2(_0892_),
    .A3(_0893_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2617_ (.A1(_0878_),
    .A2(_0892_),
    .Z(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2618_ (.A1(_0891_),
    .A2(_0894_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2619_ (.A1(\u1.row_sel[2] ),
    .A2(\u1.row_sel[1] ),
    .A3(_0892_),
    .Z(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2620_ (.A1(\u1.row_sel[1] ),
    .A2(_0892_),
    .B(\u1.row_sel[2] ),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2621_ (.A1(_0890_),
    .A2(_0895_),
    .A3(_0896_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2622_ (.A1(\u1.row_sel[3] ),
    .A2(_0895_),
    .Z(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2623_ (.A1(\u1.row_sel[3] ),
    .A2(_0895_),
    .ZN(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2624_ (.A1(_0890_),
    .A2(_0897_),
    .A3(_0898_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2625_ (.A1(net217),
    .A2(_0897_),
    .ZN(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2626_ (.A1(net217),
    .A2(_0897_),
    .Z(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2627_ (.A1(_0890_),
    .A2(_0899_),
    .A3(_0900_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2628_ (.I(net216),
    .ZN(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2629_ (.A1(_0901_),
    .A2(_0900_),
    .Z(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2630_ (.A1(_0891_),
    .A2(_0902_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2631_ (.A1(net216),
    .A2(_0900_),
    .B(\u1.row_sel[6] ),
    .ZN(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2632_ (.A1(_0891_),
    .A2(_0903_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2633_ (.A1(\latch_data_sync[0] ),
    .A2(latch_data),
    .A3(\latch_data_sync[1] ),
    .A4(_1042_),
    .Z(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2634_ (.I(_0904_),
    .Z(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2635_ (.A1(_1156_),
    .A2(_0815_),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2636_ (.I(net20),
    .ZN(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2637_ (.A1(_0905_),
    .A2(net38),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2638_ (.A1(\u1.ccr1[11] ),
    .A2(_1269_),
    .B1(\u1.ccr1[10] ),
    .B2(_1268_),
    .ZN(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2639_ (.A1(_0906_),
    .A2(_1270_),
    .ZN(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2640_ (.A1(_1274_),
    .A2(_1251_),
    .A3(_1275_),
    .B(_0907_),
    .ZN(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2641_ (.A1(_1252_),
    .A2(_1303_),
    .ZN(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2642_ (.A1(_1255_),
    .A2(_0909_),
    .B1(_1260_),
    .B2(_1264_),
    .ZN(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2643_ (.A1(\u1.ccr1[7] ),
    .A2(_1193_),
    .ZN(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2644_ (.A1(_1200_),
    .A2(_1188_),
    .B1(_1196_),
    .B2(_1190_),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2645_ (.A1(_0912_),
    .A2(_1198_),
    .B(_1201_),
    .ZN(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2646_ (.A1(_1210_),
    .A2(_1218_),
    .B(_1205_),
    .ZN(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2647_ (.A1(_1216_),
    .A2(_0914_),
    .B(_1219_),
    .C(_1202_),
    .ZN(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2648_ (.A1(_0911_),
    .A2(_0913_),
    .B(_0915_),
    .ZN(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2649_ (.A1(_1277_),
    .A2(_0916_),
    .ZN(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2650_ (.A1(_1266_),
    .A2(_0908_),
    .B(_0910_),
    .C(_0917_),
    .ZN(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2651_ (.A1(_1227_),
    .A2(_1231_),
    .Z(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2652_ (.A1(_0434_),
    .A2(_1318_),
    .B(_1321_),
    .ZN(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2653_ (.A1(_1241_),
    .A2(_1238_),
    .A3(_1242_),
    .ZN(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2654_ (.A1(_0434_),
    .A2(\u1.timer[19] ),
    .ZN(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2655_ (.A1(\u1.ccr1[18] ),
    .A2(_0920_),
    .B(_0921_),
    .C(_0922_),
    .ZN(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2656_ (.A1(\u1.ccr1[23] ),
    .A2(_1228_),
    .B(_1227_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2657_ (.A1(_0919_),
    .A2(_1234_),
    .B1(_1235_),
    .B2(_0923_),
    .C(_0924_),
    .ZN(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2658_ (.A1(_1246_),
    .A2(_0918_),
    .B(_0925_),
    .ZN(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2659_ (.A1(_1187_),
    .A2(_0926_),
    .ZN(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2660_ (.A1(\u1.ccr1[25] ),
    .A2(_1164_),
    .B1(\u1.ccr1[24] ),
    .B2(_1166_),
    .ZN(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2661_ (.A1(_0928_),
    .A2(_1181_),
    .A3(_1183_),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2662_ (.A1(\u1.ccr1[28] ),
    .A2(_1173_),
    .B1(\u1.ccr1[27] ),
    .B2(_1349_),
    .C1(_1179_),
    .C2(_0929_),
    .ZN(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2663_ (.A1(_1169_),
    .A2(_1172_),
    .B1(_1175_),
    .B2(_0930_),
    .C(_1185_),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2664_ (.A1(_1402_),
    .A2(_0927_),
    .A3(_0931_),
    .ZN(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2665_ (.A1(_1279_),
    .A2(_0932_),
    .Z(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2666_ (.I(_0933_),
    .Z(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2667_ (.I(_0934_),
    .Z(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2668_ (.A1(_1206_),
    .A2(_0935_),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2669_ (.A1(_1364_),
    .A2(_1208_),
    .Z(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2670_ (.A1(_0935_),
    .A2(_0936_),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2671_ (.I(_0933_),
    .Z(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2672_ (.A1(_1364_),
    .A2(_1363_),
    .A3(_1204_),
    .ZN(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2673_ (.A1(_1206_),
    .A2(_1208_),
    .B(_1203_),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2674_ (.A1(_0937_),
    .A2(_0938_),
    .A3(_0939_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2675_ (.A1(_1214_),
    .A2(_0938_),
    .ZN(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2676_ (.A1(\u1.timer[0] ),
    .A2(\u1.timer[1] ),
    .A3(\u1.timer[3] ),
    .A4(\u1.timer[2] ),
    .Z(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2677_ (.A1(_0937_),
    .A2(_0940_),
    .A3(_0941_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2678_ (.A1(_1287_),
    .A2(_0941_),
    .Z(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2679_ (.A1(_1287_),
    .A2(_0941_),
    .ZN(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2680_ (.A1(_0937_),
    .A2(_0942_),
    .A3(_0943_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2681_ (.A1(_1191_),
    .A2(_0942_),
    .Z(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2682_ (.A1(_0935_),
    .A2(_0944_),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2683_ (.I(_0933_),
    .Z(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2684_ (.I(_0945_),
    .Z(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2685_ (.A1(\u1.timer[6] ),
    .A2(\u1.timer[5] ),
    .Z(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2686_ (.A1(_0942_),
    .A2(_0947_),
    .Z(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2687_ (.A1(_1283_),
    .A2(_0942_),
    .B(_1280_),
    .ZN(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2688_ (.A1(_0946_),
    .A2(_0948_),
    .A3(_0949_),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2689_ (.A1(\u1.timer[7] ),
    .A2(\u1.timer[4] ),
    .A3(_0941_),
    .A4(_0947_),
    .Z(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2690_ (.I(_0950_),
    .Z(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2691_ (.A1(_1289_),
    .A2(_0948_),
    .ZN(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2692_ (.A1(_0946_),
    .A2(_0951_),
    .A3(_0952_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2693_ (.A1(_1250_),
    .A2(_0951_),
    .ZN(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2694_ (.A1(_1250_),
    .A2(_0951_),
    .Z(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2695_ (.A1(_0946_),
    .A2(_0953_),
    .A3(_0954_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2696_ (.A1(_1293_),
    .A2(_1267_),
    .ZN(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2697_ (.A1(_0951_),
    .A2(_0955_),
    .Z(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2698_ (.A1(_1248_),
    .A2(_0954_),
    .ZN(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2699_ (.A1(_0946_),
    .A2(_0956_),
    .A3(_0957_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2700_ (.I(_0945_),
    .Z(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2701_ (.A1(_1295_),
    .A2(_0956_),
    .Z(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2702_ (.A1(_1295_),
    .A2(_0956_),
    .ZN(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2703_ (.A1(_0958_),
    .A2(_0959_),
    .A3(_0960_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2704_ (.A1(_1272_),
    .A2(\u1.timer[10] ),
    .A3(_0950_),
    .A4(_0955_),
    .Z(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2705_ (.A1(_1272_),
    .A2(_0959_),
    .ZN(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2706_ (.A1(_0958_),
    .A2(_0961_),
    .A3(_0962_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2707_ (.A1(_1311_),
    .A2(_0961_),
    .Z(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2708_ (.A1(_1311_),
    .A2(_0961_),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2709_ (.A1(_0958_),
    .A2(_0963_),
    .A3(_0964_),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2710_ (.A1(_1258_),
    .A2(_0963_),
    .Z(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2711_ (.A1(_0935_),
    .A2(_0965_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2712_ (.A1(_1254_),
    .A2(_1300_),
    .A3(_1262_),
    .A4(_0961_),
    .Z(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2713_ (.A1(_1300_),
    .A2(_0963_),
    .B(_1254_),
    .ZN(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2714_ (.A1(_0958_),
    .A2(_0966_),
    .A3(_0967_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2715_ (.I(_0945_),
    .Z(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2716_ (.A1(_1303_),
    .A2(_0966_),
    .ZN(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2717_ (.A1(_1303_),
    .A2(_0966_),
    .Z(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2718_ (.I(_0970_),
    .Z(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2719_ (.A1(_0968_),
    .A2(_0969_),
    .A3(_0971_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2720_ (.A1(_0283_),
    .A2(_0971_),
    .ZN(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2721_ (.A1(_1279_),
    .A2(_0932_),
    .B1(_0971_),
    .B2(_0283_),
    .C(_0972_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2722_ (.A1(_0283_),
    .A2(_0971_),
    .B(_0282_),
    .ZN(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2723_ (.A1(_0282_),
    .A2(\u1.timer[16] ),
    .A3(_0970_),
    .Z(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2724_ (.A1(_0968_),
    .A2(_0973_),
    .A3(_0974_),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2725_ (.A1(_1322_),
    .A2(_0974_),
    .ZN(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2726_ (.A1(_1321_),
    .A2(_0282_),
    .A3(\u1.timer[16] ),
    .A4(_0970_),
    .Z(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2727_ (.A1(_0968_),
    .A2(_0975_),
    .A3(_0976_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2728_ (.A1(_0281_),
    .A2(_0976_),
    .ZN(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2729_ (.A1(_0281_),
    .A2(_1322_),
    .A3(_0974_),
    .Z(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2730_ (.A1(_0968_),
    .A2(_0977_),
    .A3(_0978_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2731_ (.A1(_1224_),
    .A2(_0978_),
    .Z(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2732_ (.A1(_0937_),
    .A2(_0979_),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2733_ (.A1(\u1.timer[20] ),
    .A2(_0978_),
    .ZN(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2734_ (.A1(\u1.timer[21] ),
    .A2(\u1.timer[20] ),
    .A3(_0281_),
    .A4(_0976_),
    .Z(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2735_ (.I(_0945_),
    .Z(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2736_ (.A1(_1233_),
    .A2(_0980_),
    .B(_0981_),
    .C(_0982_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2737_ (.I(_0933_),
    .Z(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2738_ (.A1(_0286_),
    .A2(_0981_),
    .ZN(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2739_ (.A1(_0286_),
    .A2(_0981_),
    .Z(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2740_ (.A1(_0983_),
    .A2(_0984_),
    .A3(_0985_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2741_ (.A1(_0285_),
    .A2(_0985_),
    .ZN(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2742_ (.A1(_0285_),
    .A2(_0985_),
    .B(_0986_),
    .C(_0982_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2743_ (.A1(_0285_),
    .A2(_0985_),
    .B(\u1.timer[24] ),
    .ZN(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2744_ (.A1(\u1.timer[24] ),
    .A2(_1327_),
    .A3(_0286_),
    .A4(_0981_),
    .Z(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2745_ (.A1(_0983_),
    .A2(_0987_),
    .A3(_0988_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2746_ (.A1(_1411_),
    .A2(_0988_),
    .ZN(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2747_ (.A1(_1411_),
    .A2(_0988_),
    .Z(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2748_ (.A1(_0983_),
    .A2(_0989_),
    .A3(_0990_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2749_ (.A1(_1410_),
    .A2(_0990_),
    .ZN(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2750_ (.A1(_1410_),
    .A2(_0990_),
    .B(_0991_),
    .C(_0982_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2751_ (.A1(_1410_),
    .A2(_0990_),
    .B(_1394_),
    .ZN(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2752_ (.A1(_1394_),
    .A2(_1345_),
    .A3(_1411_),
    .A4(_0988_),
    .Z(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2753_ (.A1(_0983_),
    .A2(_0992_),
    .A3(_0993_),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2754_ (.A1(_1413_),
    .A2(_0993_),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2755_ (.A1(_1413_),
    .A2(_0993_),
    .Z(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2756_ (.A1(_0982_),
    .A2(_0994_),
    .A3(_0995_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2757_ (.I(\u1.timer[29] ),
    .Z(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2758_ (.A1(_0996_),
    .A2(_0995_),
    .ZN(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2759_ (.A1(_0996_),
    .A2(_0995_),
    .B(_0997_),
    .C(_0934_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2760_ (.A1(_0996_),
    .A2(_0995_),
    .ZN(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2761_ (.A1(\u1.timer[30] ),
    .A2(_0996_),
    .A3(_1413_),
    .A4(_0993_),
    .Z(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2762_ (.A1(_1167_),
    .A2(_0998_),
    .B(_0999_),
    .C(_0934_),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2763_ (.A1(_1351_),
    .A2(_0999_),
    .ZN(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2764_ (.A1(_1351_),
    .A2(_0999_),
    .B(_1000_),
    .C(_0934_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2765_ (.I(net12),
    .ZN(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2766_ (.A1(_1001_),
    .A2(net30),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2767_ (.I(net11),
    .ZN(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2768_ (.A1(_1002_),
    .A2(net29),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2769_ (.I(net10),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2770_ (.A1(_1003_),
    .A2(net28),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2771_ (.I(net9),
    .ZN(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2772_ (.A1(_1004_),
    .A2(net27),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2773_ (.I(net8),
    .ZN(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2774_ (.A1(_1005_),
    .A2(net26),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2775_ (.I(net7),
    .ZN(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2776_ (.A1(_1006_),
    .A2(net25),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2777_ (.I(net6),
    .ZN(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2778_ (.A1(_1007_),
    .A2(net24),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2779_ (.I(net5),
    .ZN(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2780_ (.A1(_1008_),
    .A2(net23),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2781_ (.I(net21),
    .ZN(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2782_ (.A1(_1009_),
    .A2(net39),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2783_ (.I(\u1.ccr0[0] ),
    .ZN(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2784_ (.A1(_0393_),
    .A2(_0394_),
    .A3(_0351_),
    .ZN(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2785_ (.I(_1011_),
    .Z(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2786_ (.I(_1012_),
    .Z(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2787_ (.I(_1013_),
    .Z(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2788_ (.I(_1012_),
    .Z(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2789_ (.A1(_0392_),
    .A2(_1015_),
    .ZN(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2790_ (.A1(_1010_),
    .A2(_1014_),
    .B(_1016_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2791_ (.I(_1011_),
    .Z(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2792_ (.I0(\u1.ccr0[1] ),
    .I1(_0400_),
    .S(_1017_),
    .Z(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2793_ (.I(_1018_),
    .Z(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2794_ (.I0(\u1.ccr0[2] ),
    .I1(_0361_),
    .S(_1017_),
    .Z(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2795_ (.I(_1019_),
    .Z(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2796_ (.I0(\u1.ccr0[3] ),
    .I1(_0364_),
    .S(_1013_),
    .Z(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2797_ (.I(_1020_),
    .Z(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2798_ (.I(_1012_),
    .Z(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2799_ (.A1(_0409_),
    .A2(_1021_),
    .ZN(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2800_ (.A1(_1286_),
    .A2(_1014_),
    .B(_1022_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2801_ (.A1(_0411_),
    .A2(_1021_),
    .ZN(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2802_ (.A1(_1282_),
    .A2(_1014_),
    .B(_1023_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2803_ (.A1(_0470_),
    .A2(_1021_),
    .ZN(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2804_ (.A1(_1281_),
    .A2(_1014_),
    .B(_1024_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2805_ (.I(_1012_),
    .Z(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2806_ (.A1(_0373_),
    .A2(_1021_),
    .ZN(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2807_ (.A1(_1290_),
    .A2(_1025_),
    .B(_1026_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2808_ (.I0(\u1.ccr0[8] ),
    .I1(_0375_),
    .S(_1013_),
    .Z(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2809_ (.I(_1027_),
    .Z(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2810_ (.I0(\u1.ccr0[9] ),
    .I1(_0377_),
    .S(_1013_),
    .Z(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2811_ (.I(_1028_),
    .Z(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2812_ (.I(_1011_),
    .Z(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2813_ (.A1(net224),
    .A2(_1029_),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2814_ (.A1(_1296_),
    .A2(_1025_),
    .B(_1030_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2815_ (.I(\u1.ccr0[11] ),
    .ZN(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2816_ (.A1(net223),
    .A2(_1029_),
    .ZN(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2817_ (.A1(_1031_),
    .A2(_1025_),
    .B(_1032_),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2818_ (.A1(\u0.cmd[12] ),
    .A2(_1029_),
    .ZN(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2819_ (.A1(_1310_),
    .A2(_1025_),
    .B(_1033_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2820_ (.A1(net221),
    .A2(_1029_),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2821_ (.A1(_1301_),
    .A2(_1015_),
    .B(_1034_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2822_ (.A1(net220),
    .A2(_1017_),
    .ZN(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2823_ (.A1(_1305_),
    .A2(_1015_),
    .B(_1035_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2824_ (.A1(net219),
    .A2(_1017_),
    .ZN(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2825_ (.A1(_1304_),
    .A2(_1015_),
    .B(_1036_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2826_ (.A1(net4),
    .A2(net22),
    .Z(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2827_ (.I(_1037_),
    .Z(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2828_ (.A1(net13),
    .A2(net31),
    .Z(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2829_ (.I(_1038_),
    .Z(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2830_ (.A1(net14),
    .A2(net32),
    .Z(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2831_ (.I(_1039_),
    .Z(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2832_ (.D(net292),
    .CLK(clknet_leaf_10_clock),
    .Q(net204));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2833_ (.D(net293),
    .CLK(clknet_leaf_10_clock),
    .Q(net205));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2834_ (.D(\u1.row_sel[2] ),
    .CLK(clknet_leaf_9_clock),
    .Q(net206));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2835_ (.D(\u1.row_sel[3] ),
    .CLK(clknet_leaf_10_clock),
    .Q(net207));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2836_ (.D(net271),
    .CLK(clknet_leaf_10_clock),
    .Q(net208));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2837_ (.D(net276),
    .CLK(clknet_leaf_10_clock),
    .Q(net209));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2838_ (.D(net268),
    .CLK(clknet_leaf_15_clock),
    .Q(net83));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2839_ (.D(net295),
    .CLK(clknet_leaf_10_clock),
    .Q(net84));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2840_ (.D(net225),
    .CLK(clknet_leaf_15_clock),
    .Q(net85));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2841_ (.D(\u1.col_sel[3] ),
    .CLK(clknet_leaf_15_clock),
    .Q(net86));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2842_ (.D(net294),
    .CLK(clknet_leaf_15_clock),
    .Q(net87));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2843_ (.D(\u1.col_sel[5] ),
    .CLK(clknet_leaf_15_clock),
    .Q(net88));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2844_ (.D(\u0.cmd[0] ),
    .CLK(clknet_leaf_15_clock),
    .Q(net95));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2845_ (.D(\u0.cmd[1] ),
    .CLK(clknet_leaf_15_clock),
    .Q(net102));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2846_ (.D(\u0.cmd[2] ),
    .CLK(clknet_leaf_15_clock),
    .Q(net103));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2847_ (.D(net288),
    .CLK(clknet_leaf_10_clock),
    .Q(net104));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2848_ (.D(net290),
    .CLK(clknet_leaf_16_clock),
    .Q(net105));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2849_ (.D(net289),
    .CLK(clknet_leaf_16_clock),
    .Q(net106));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2850_ (.D(\u0.cmd[6] ),
    .CLK(clknet_leaf_15_clock),
    .Q(net107));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2851_ (.D(\u0.cmd[7] ),
    .CLK(clknet_leaf_15_clock),
    .Q(net108));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2852_ (.D(\u0.cmd[8] ),
    .CLK(clknet_leaf_16_clock),
    .Q(net109));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2853_ (.D(\u0.cmd[9] ),
    .CLK(clknet_leaf_16_clock),
    .Q(net110));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2854_ (.D(net224),
    .CLK(clknet_leaf_16_clock),
    .Q(net96));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2855_ (.D(net223),
    .CLK(clknet_leaf_16_clock),
    .Q(net97));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2856_ (.D(net222),
    .CLK(clknet_leaf_16_clock),
    .Q(net98));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2857_ (.D(net221),
    .CLK(clknet_leaf_15_clock),
    .Q(net99));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2858_ (.D(net220),
    .CLK(clknet_leaf_16_clock),
    .Q(net100));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2859_ (.D(net219),
    .CLK(clknet_leaf_16_clock),
    .Q(net101));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2860_ (.D(net249),
    .CLK(clknet_leaf_9_clock),
    .Q(net192));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2861_ (.D(net243),
    .CLK(clknet_leaf_5_clock),
    .Q(\latch_data_sync[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2862_ (.D(net272),
    .CLK(clknet_leaf_5_clock),
    .Q(\latch_data_sync[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2863_ (.D(net250),
    .CLK(clknet_leaf_4_clock),
    .Q(\control_trigger_sync[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2864_ (.D(net291),
    .CLK(clknet_leaf_4_clock),
    .Q(\control_trigger_sync[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2865_ (.D(net270),
    .CLK(clknet_leaf_33_clock),
    .Q(\reset_n_sync[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2866_ (.D(net259),
    .CLK(clknet_leaf_34_clock),
    .Q(\reset_n_sync[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2867_ (.D(_0024_),
    .CLK(clknet_leaf_32_clock),
    .Q(net160));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2868_ (.D(_0025_),
    .CLK(clknet_leaf_11_clock),
    .Q(\u1.col_sel[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2869_ (.D(_0026_),
    .CLK(clknet_leaf_10_clock),
    .Q(\u1.col_sel[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2870_ (.D(_0027_),
    .CLK(clknet_leaf_14_clock),
    .Q(\u1.col_sel[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2871_ (.D(_0028_),
    .CLK(clknet_leaf_15_clock),
    .Q(\u1.col_sel[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2872_ (.D(_0029_),
    .CLK(clknet_leaf_14_clock),
    .Q(\u1.col_sel[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2873_ (.D(_0030_),
    .CLK(clknet_leaf_16_clock),
    .Q(\u1.col_sel[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2874_ (.D(_0031_),
    .CLK(clknet_leaf_16_clock),
    .Q(\u1.col_sel[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2875_ (.D(\u0.latch_cmd ),
    .CLK(clknet_leaf_4_clock),
    .Q(\u0.update_cmd ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2876_ (.D(_0022_),
    .CLK(clknet_leaf_6_clock),
    .Q(\u0.write_config_n ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2877_ (.D(_0011_),
    .CLK(clknet_leaf_12_clock),
    .Q(\u0.timer_enable ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2878_ (.D(_0012_),
    .CLK(clknet_leaf_7_clock),
    .Q(\u0.mem_write_n[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2879_ (.D(_0013_),
    .CLK(clknet_leaf_7_clock),
    .Q(\u0.mem_write_n[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2880_ (.D(_0014_),
    .CLK(clknet_leaf_8_clock),
    .Q(\u0.mem_write_n[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2881_ (.D(_0015_),
    .CLK(clknet_leaf_8_clock),
    .Q(\u0.mem_write_n[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2882_ (.D(_0016_),
    .CLK(clknet_leaf_8_clock),
    .Q(\u0.mem_write_n[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2883_ (.D(_0017_),
    .CLK(clknet_leaf_9_clock),
    .Q(\u0.mem_write_n[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2884_ (.D(_0018_),
    .CLK(clknet_leaf_8_clock),
    .Q(\u0.mem_write_n[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2885_ (.D(_0019_),
    .CLK(clknet_leaf_8_clock),
    .Q(\u0.mem_write_n[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2886_ (.D(_0020_),
    .CLK(clknet_leaf_8_clock),
    .Q(\u0.mem_write_n[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2887_ (.D(_0021_),
    .CLK(clknet_leaf_8_clock),
    .Q(\u0.mem_write_n[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2888_ (.D(\u1.ccr1_flag ),
    .CLK(clknet_leaf_3_clock),
    .Q(\u1.u1.impulse_gen[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2889_ (.D(net279),
    .CLK(clknet_leaf_3_clock),
    .Q(\u1.u1.impulse_gen[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2890_ (.D(_0032_),
    .CLK(clknet_leaf_3_clock),
    .Q(\u1.ccr0[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2891_ (.D(_0033_),
    .CLK(clknet_leaf_2_clock),
    .Q(\u1.ccr0[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2892_ (.D(_0034_),
    .CLK(clknet_leaf_2_clock),
    .Q(\u1.ccr0[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2893_ (.D(_0035_),
    .CLK(clknet_leaf_2_clock),
    .Q(\u1.ccr0[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2894_ (.D(_0036_),
    .CLK(clknet_leaf_2_clock),
    .Q(\u1.ccr0[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2895_ (.D(_0037_),
    .CLK(clknet_leaf_3_clock),
    .Q(\u1.ccr0[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2896_ (.D(_0038_),
    .CLK(clknet_leaf_2_clock),
    .Q(\u1.ccr0[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2897_ (.D(_0039_),
    .CLK(clknet_leaf_2_clock),
    .Q(\u1.ccr0[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2898_ (.D(_0040_),
    .CLK(clknet_leaf_0_clock),
    .Q(\u1.ccr0[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2899_ (.D(_0041_),
    .CLK(clknet_leaf_36_clock),
    .Q(\u1.ccr0[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2900_ (.D(_0042_),
    .CLK(clknet_leaf_34_clock),
    .Q(\u1.ccr0[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2901_ (.D(_0043_),
    .CLK(clknet_leaf_34_clock),
    .Q(\u1.ccr0[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2902_ (.D(_0044_),
    .CLK(clknet_leaf_36_clock),
    .Q(\u1.ccr0[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2903_ (.D(_0045_),
    .CLK(clknet_leaf_36_clock),
    .Q(\u1.ccr0[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2904_ (.D(_0046_),
    .CLK(clknet_leaf_36_clock),
    .Q(\u1.ccr0[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2905_ (.D(_0047_),
    .CLK(clknet_leaf_0_clock),
    .Q(\u1.ccr0[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2906_ (.D(_0048_),
    .CLK(clknet_leaf_30_clock),
    .Q(\u1.ccr1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2907_ (.D(_0049_),
    .CLK(clknet_leaf_30_clock),
    .Q(\u1.ccr1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2908_ (.D(_0050_),
    .CLK(clknet_leaf_22_clock),
    .Q(\u1.ccr1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2909_ (.D(_0051_),
    .CLK(clknet_leaf_22_clock),
    .Q(\u1.ccr1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2910_ (.D(_0052_),
    .CLK(clknet_leaf_24_clock),
    .Q(\u1.ccr1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2911_ (.D(_0053_),
    .CLK(clknet_leaf_24_clock),
    .Q(\u1.ccr1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2912_ (.D(_0054_),
    .CLK(clknet_leaf_24_clock),
    .Q(\u1.ccr1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2913_ (.D(_0055_),
    .CLK(clknet_leaf_25_clock),
    .Q(\u1.ccr1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2914_ (.D(_0056_),
    .CLK(clknet_leaf_25_clock),
    .Q(\u1.ccr1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2915_ (.D(_0057_),
    .CLK(clknet_leaf_26_clock),
    .Q(\u1.ccr1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2916_ (.D(_0058_),
    .CLK(clknet_leaf_26_clock),
    .Q(\u1.ccr1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2917_ (.D(_0059_),
    .CLK(clknet_leaf_26_clock),
    .Q(\u1.ccr1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2918_ (.D(_0060_),
    .CLK(clknet_leaf_27_clock),
    .Q(\u1.ccr1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2919_ (.D(_0061_),
    .CLK(clknet_leaf_27_clock),
    .Q(\u1.ccr1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2920_ (.D(_0062_),
    .CLK(clknet_leaf_28_clock),
    .Q(\u1.ccr1[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2921_ (.D(_0063_),
    .CLK(clknet_leaf_29_clock),
    .Q(\u1.ccr1[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2922_ (.D(_0064_),
    .CLK(clknet_leaf_2_clock),
    .Q(\u1.ccr1[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2923_ (.D(_0065_),
    .CLK(clknet_leaf_2_clock),
    .Q(\u1.ccr1[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2924_ (.D(_0066_),
    .CLK(clknet_leaf_3_clock),
    .Q(\u1.ccr1[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2925_ (.D(_0067_),
    .CLK(clknet_leaf_30_clock),
    .Q(\u1.ccr1[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2926_ (.D(_0068_),
    .CLK(clknet_leaf_3_clock),
    .Q(\u1.ccr1[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2927_ (.D(_0069_),
    .CLK(clknet_leaf_2_clock),
    .Q(\u1.ccr1[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2928_ (.D(_0070_),
    .CLK(clknet_leaf_31_clock),
    .Q(\u1.ccr1[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2929_ (.D(_0071_),
    .CLK(clknet_leaf_2_clock),
    .Q(\u1.ccr1[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2930_ (.D(_0072_),
    .CLK(clknet_leaf_2_clock),
    .Q(\u1.ccr1[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2931_ (.D(_0073_),
    .CLK(clknet_leaf_0_clock),
    .Q(\u1.ccr1[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2932_ (.D(_0074_),
    .CLK(clknet_2_0__leaf_clock),
    .Q(\u1.ccr1[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2933_ (.D(_0075_),
    .CLK(clknet_leaf_2_clock),
    .Q(\u1.ccr1[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2934_ (.D(_0076_),
    .CLK(clknet_leaf_0_clock),
    .Q(\u1.ccr1[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2935_ (.D(_0077_),
    .CLK(clknet_leaf_0_clock),
    .Q(\u1.ccr1[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2936_ (.D(_0078_),
    .CLK(clknet_leaf_0_clock),
    .Q(\u1.ccr1[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2937_ (.D(_0079_),
    .CLK(clknet_leaf_0_clock),
    .Q(\u1.ccr1[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2938_ (.D(_0080_),
    .CLK(clknet_leaf_12_clock),
    .Q(\u1.ordering_complete[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2939_ (.D(_0081_),
    .CLK(clknet_leaf_4_clock),
    .Q(\u1.ordering_complete[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2940_ (.D(_0082_),
    .CLK(clknet_leaf_13_clock),
    .Q(\u1.ordering_complete[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2941_ (.D(_0083_),
    .CLK(clknet_leaf_14_clock),
    .Q(\u1.ordering_complete[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2942_ (.D(_0084_),
    .CLK(clknet_leaf_14_clock),
    .Q(\u1.ordering_complete[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2943_ (.D(_0085_),
    .CLK(clknet_leaf_14_clock),
    .Q(\u1.ordering_complete[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2944_ (.D(_0086_),
    .CLK(clknet_leaf_19_clock),
    .Q(\u1.ordering_complete[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2945_ (.D(_0087_),
    .CLK(clknet_leaf_19_clock),
    .Q(\u1.ordering_complete[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2946_ (.D(_0088_),
    .CLK(clknet_leaf_19_clock),
    .Q(\u1.ordering_complete[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2947_ (.D(_0089_),
    .CLK(clknet_leaf_20_clock),
    .Q(\u1.ordering_complete[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2948_ (.D(_0090_),
    .CLK(clknet_leaf_12_clock),
    .Q(\u1.ordering_complete[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2949_ (.D(_0091_),
    .CLK(clknet_leaf_12_clock),
    .Q(\u1.ordering_complete[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2950_ (.D(_0092_),
    .CLK(clknet_leaf_4_clock),
    .Q(\u1.ordering_complete[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2951_ (.D(_0093_),
    .CLK(clknet_leaf_4_clock),
    .Q(\u1.ordering_complete[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2952_ (.D(_0094_),
    .CLK(clknet_leaf_3_clock),
    .Q(\u1.ordering_complete[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2953_ (.D(_0095_),
    .CLK(clknet_leaf_3_clock),
    .Q(\u1.ordering_complete[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2954_ (.D(_0096_),
    .CLK(clknet_leaf_3_clock),
    .Q(\u1.ordering_complete[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2955_ (.D(_0097_),
    .CLK(clknet_leaf_3_clock),
    .Q(\u1.ordering_complete[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2956_ (.D(_0098_),
    .CLK(clknet_leaf_3_clock),
    .Q(\u1.ordering_complete[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2957_ (.D(_0099_),
    .CLK(clknet_leaf_3_clock),
    .Q(\u1.ordering_complete[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2958_ (.D(_0100_),
    .CLK(clknet_leaf_20_clock),
    .Q(\u1.ordering_complete[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2959_ (.D(_0101_),
    .CLK(clknet_leaf_20_clock),
    .Q(\u1.ordering_complete[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2960_ (.D(_0102_),
    .CLK(clknet_leaf_20_clock),
    .Q(\u1.ordering_complete[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2961_ (.D(_0103_),
    .CLK(clknet_leaf_21_clock),
    .Q(\u1.ordering_complete[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2962_ (.D(_0104_),
    .CLK(clknet_leaf_20_clock),
    .Q(\u1.ordering_complete[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2963_ (.D(_0105_),
    .CLK(clknet_leaf_20_clock),
    .Q(\u1.ordering_complete[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2964_ (.D(_0106_),
    .CLK(clknet_leaf_24_clock),
    .Q(\u1.ordering_complete[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2965_ (.D(_0107_),
    .CLK(clknet_leaf_24_clock),
    .Q(\u1.ordering_complete[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2966_ (.D(_0108_),
    .CLK(clknet_leaf_3_clock),
    .Q(\u1.ordering_complete[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2967_ (.D(_0109_),
    .CLK(clknet_leaf_23_clock),
    .Q(\u1.ordering_complete[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2968_ (.D(_0110_),
    .CLK(clknet_leaf_22_clock),
    .Q(\u1.ordering_complete[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2969_ (.D(_0111_),
    .CLK(clknet_leaf_22_clock),
    .Q(\u1.ordering_complete[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2970_ (.D(_0112_),
    .CLK(clknet_leaf_12_clock),
    .Q(\u1.row_limit[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2971_ (.D(_0113_),
    .CLK(clknet_leaf_11_clock),
    .Q(\u1.row_limit[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2972_ (.D(_0114_),
    .CLK(clknet_leaf_9_clock),
    .Q(\u1.row_limit[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2973_ (.D(_0115_),
    .CLK(clknet_leaf_11_clock),
    .Q(\u1.row_limit[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2974_ (.D(_0116_),
    .CLK(clknet_leaf_11_clock),
    .Q(\u1.row_limit[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2975_ (.D(_0117_),
    .CLK(clknet_leaf_11_clock),
    .Q(\u1.row_limit[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2976_ (.D(_0118_),
    .CLK(clknet_leaf_11_clock),
    .Q(\u1.row_limit[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2977_ (.D(_0119_),
    .CLK(clknet_leaf_11_clock),
    .Q(\u1.col_limit[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2978_ (.D(_0120_),
    .CLK(clknet_leaf_11_clock),
    .Q(\u1.col_limit[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2979_ (.D(_0121_),
    .CLK(clknet_leaf_14_clock),
    .Q(\u1.col_limit[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2980_ (.D(_0122_),
    .CLK(clknet_leaf_14_clock),
    .Q(\u1.col_limit[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2981_ (.D(_0123_),
    .CLK(clknet_leaf_16_clock),
    .Q(\u1.col_limit[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2982_ (.D(_0124_),
    .CLK(clknet_leaf_16_clock),
    .Q(\u1.col_limit[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2983_ (.D(_0125_),
    .CLK(clknet_leaf_14_clock),
    .Q(\u1.col_limit[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2984_ (.D(_0126_),
    .CLK(clknet_leaf_18_clock),
    .Q(\u1.inverter_select[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2985_ (.D(_0127_),
    .CLK(clknet_leaf_16_clock),
    .Q(\u1.inverter_select[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2986_ (.D(_0128_),
    .CLK(clknet_leaf_16_clock),
    .Q(\u1.inverter_select[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2987_ (.D(_0129_),
    .CLK(clknet_leaf_18_clock),
    .Q(\u1.inverter_select[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2988_ (.D(_0130_),
    .CLK(clknet_leaf_18_clock),
    .Q(\u1.inverter_select[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2989_ (.D(_0131_),
    .CLK(clknet_leaf_18_clock),
    .Q(\u1.inverter_select[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2990_ (.D(_0132_),
    .CLK(clknet_leaf_17_clock),
    .Q(\u1.inverter_select[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2991_ (.D(_0133_),
    .CLK(clknet_leaf_17_clock),
    .Q(\u1.inverter_select[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2992_ (.D(_0134_),
    .CLK(clknet_leaf_18_clock),
    .Q(\u1.inverter_select[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2993_ (.D(_0135_),
    .CLK(clknet_leaf_18_clock),
    .Q(\u1.inverter_select[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2994_ (.D(_0136_),
    .CLK(clknet_leaf_16_clock),
    .Q(\u1.row_col_select[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2995_ (.D(_0137_),
    .CLK(clknet_leaf_16_clock),
    .Q(\u1.row_col_select[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2996_ (.D(_0138_),
    .CLK(clknet_leaf_16_clock),
    .Q(\u1.row_col_select[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2997_ (.D(_0139_),
    .CLK(clknet_leaf_16_clock),
    .Q(\u1.row_col_select[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2998_ (.D(_0140_),
    .CLK(clknet_leaf_18_clock),
    .Q(\u1.row_col_select[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2999_ (.D(_0141_),
    .CLK(clknet_leaf_18_clock),
    .Q(\u1.row_col_select[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3000_ (.D(_0142_),
    .CLK(clknet_leaf_18_clock),
    .Q(\u1.row_col_select[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3001_ (.D(_0143_),
    .CLK(clknet_leaf_17_clock),
    .Q(\u1.row_col_select[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3002_ (.D(_0144_),
    .CLK(clknet_leaf_18_clock),
    .Q(\u1.row_col_select[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3003_ (.D(_0145_),
    .CLK(clknet_leaf_18_clock),
    .Q(\u1.row_col_select[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3004_ (.D(_0146_),
    .CLK(clknet_leaf_13_clock),
    .Q(\u1.ordering_timer[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3005_ (.D(_0147_),
    .CLK(clknet_leaf_12_clock),
    .Q(\u1.ordering_timer[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3006_ (.D(_0148_),
    .CLK(clknet_leaf_12_clock),
    .Q(\u1.ordering_timer[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3007_ (.D(_0149_),
    .CLK(clknet_leaf_12_clock),
    .Q(\u1.ordering_timer[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3008_ (.D(_0150_),
    .CLK(clknet_leaf_14_clock),
    .Q(\u1.ordering_timer[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3009_ (.D(_0151_),
    .CLK(clknet_leaf_16_clock),
    .Q(\u1.ordering_timer[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3010_ (.D(_0152_),
    .CLK(clknet_leaf_19_clock),
    .Q(\u1.ordering_timer[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3011_ (.D(_0153_),
    .CLK(clknet_leaf_19_clock),
    .Q(\u1.ordering_timer[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3012_ (.D(_0154_),
    .CLK(clknet_leaf_19_clock),
    .Q(\u1.ordering_timer[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3013_ (.D(_0155_),
    .CLK(clknet_leaf_19_clock),
    .Q(\u1.ordering_timer[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3014_ (.D(_0156_),
    .CLK(clknet_leaf_21_clock),
    .Q(\u1.ordering_timer[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3015_ (.D(_0157_),
    .CLK(clknet_leaf_14_clock),
    .Q(\u1.ordering_timer[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3016_ (.D(_0158_),
    .CLK(clknet_leaf_14_clock),
    .Q(\u1.ordering_timer[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3017_ (.D(_0159_),
    .CLK(clknet_leaf_13_clock),
    .Q(\u1.ordering_timer[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3018_ (.D(_0160_),
    .CLK(clknet_leaf_13_clock),
    .Q(\u1.ordering_timer[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3019_ (.D(_0161_),
    .CLK(clknet_leaf_13_clock),
    .Q(\u1.ordering_timer[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3020_ (.D(_0162_),
    .CLK(clknet_leaf_13_clock),
    .Q(\u1.ordering_timer[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3021_ (.D(_0163_),
    .CLK(clknet_leaf_13_clock),
    .Q(\u1.ordering_timer[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3022_ (.D(_0164_),
    .CLK(clknet_leaf_30_clock),
    .Q(\u1.ordering_timer[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3023_ (.D(_0165_),
    .CLK(clknet_leaf_21_clock),
    .Q(\u1.ordering_timer[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3024_ (.D(_0166_),
    .CLK(clknet_leaf_21_clock),
    .Q(\u1.ordering_timer[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3025_ (.D(_0167_),
    .CLK(clknet_leaf_20_clock),
    .Q(\u1.ordering_timer[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3026_ (.D(_0168_),
    .CLK(clknet_leaf_20_clock),
    .Q(\u1.ordering_timer[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3027_ (.D(_0169_),
    .CLK(clknet_leaf_20_clock),
    .Q(\u1.ordering_timer[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3028_ (.D(_0170_),
    .CLK(clknet_leaf_24_clock),
    .Q(\u1.ordering_timer[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3029_ (.D(_0171_),
    .CLK(clknet_leaf_24_clock),
    .Q(\u1.ordering_timer[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3030_ (.D(_0172_),
    .CLK(clknet_leaf_24_clock),
    .Q(\u1.ordering_timer[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3031_ (.D(_0173_),
    .CLK(clknet_leaf_24_clock),
    .Q(\u1.ordering_timer[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3032_ (.D(_0174_),
    .CLK(clknet_leaf_21_clock),
    .Q(\u1.ordering_timer[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3033_ (.D(_0175_),
    .CLK(clknet_leaf_22_clock),
    .Q(\u1.ordering_timer[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3034_ (.D(_0176_),
    .CLK(clknet_leaf_22_clock),
    .Q(\u1.ordering_timer[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3035_ (.D(_0177_),
    .CLK(clknet_leaf_22_clock),
    .Q(\u1.ordering_timer[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3036_ (.D(_0178_),
    .CLK(clknet_leaf_3_clock),
    .Q(\u0.cmd[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3037_ (.D(_0179_),
    .CLK(clknet_leaf_3_clock),
    .Q(\u0.cmd[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3038_ (.D(_0180_),
    .CLK(clknet_leaf_3_clock),
    .Q(\u0.cmd[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3039_ (.D(_0181_),
    .CLK(clknet_leaf_4_clock),
    .Q(\u0.cmd[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3040_ (.D(_0182_),
    .CLK(clknet_leaf_4_clock),
    .Q(\u0.cmd[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3041_ (.D(_0183_),
    .CLK(clknet_leaf_4_clock),
    .Q(\u0.cmd[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3042_ (.D(_0184_),
    .CLK(clknet_leaf_3_clock),
    .Q(\u0.cmd[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3043_ (.D(_0185_),
    .CLK(clknet_leaf_3_clock),
    .Q(\u0.cmd[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3044_ (.D(_0186_),
    .CLK(clknet_leaf_1_clock),
    .Q(\u0.cmd[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3045_ (.D(_0187_),
    .CLK(clknet_leaf_1_clock),
    .Q(\u0.cmd[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3046_ (.D(_0188_),
    .CLK(clknet_leaf_1_clock),
    .Q(\u0.cmd[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3047_ (.D(_0189_),
    .CLK(clknet_leaf_1_clock),
    .Q(\u0.cmd[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3048_ (.D(_0190_),
    .CLK(clknet_leaf_5_clock),
    .Q(\u0.cmd[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3049_ (.D(_0191_),
    .CLK(clknet_leaf_4_clock),
    .Q(\u0.cmd[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3050_ (.D(_0192_),
    .CLK(clknet_leaf_1_clock),
    .Q(\u0.cmd[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3051_ (.D(_0193_),
    .CLK(clknet_leaf_1_clock),
    .Q(\u0.cmd[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3052_ (.D(_0194_),
    .CLK(clknet_leaf_5_clock),
    .Q(\u0.cmd[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3053_ (.D(_0195_),
    .CLK(clknet_leaf_5_clock),
    .Q(\u0.cmd[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3054_ (.D(_0196_),
    .CLK(clknet_leaf_5_clock),
    .Q(\u0.cmd[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3055_ (.D(_0197_),
    .CLK(clknet_leaf_5_clock),
    .Q(\u0.cmd[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _3056_ (.D(_0198_),
    .CLK(clknet_leaf_5_clock),
    .Q(\u0.cmd[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _3057_ (.D(_0199_),
    .CLK(clknet_leaf_5_clock),
    .Q(\u0.cmd[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3058_ (.D(_0200_),
    .CLK(clknet_leaf_6_clock),
    .Q(\u0.cmd[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3059_ (.D(_0201_),
    .CLK(clknet_leaf_6_clock),
    .Q(\u0.cmd[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3060_ (.D(_0202_),
    .CLK(clknet_leaf_7_clock),
    .Q(\u0.cmd[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3061_ (.D(_0203_),
    .CLK(clknet_leaf_7_clock),
    .Q(\u0.cmd[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3062_ (.D(_0204_),
    .CLK(clknet_leaf_8_clock),
    .Q(\u0.cmd[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3063_ (.D(_0205_),
    .CLK(clknet_leaf_6_clock),
    .Q(\u0.cmd[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3064_ (.D(_0206_),
    .CLK(clknet_leaf_6_clock),
    .Q(\u0.cmd[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3065_ (.D(_0207_),
    .CLK(clknet_leaf_6_clock),
    .Q(\u0.cmd[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3066_ (.D(_0208_),
    .CLK(clknet_leaf_6_clock),
    .Q(\u0.cmd[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3067_ (.D(_0209_),
    .CLK(clknet_leaf_6_clock),
    .Q(\u0.cmd[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3068_ (.D(_0023_),
    .CLK(clknet_leaf_4_clock),
    .Q(\u1.output_active ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3069_ (.D(_0210_),
    .CLK(clknet_leaf_9_clock),
    .Q(\u1.row_sel[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3070_ (.D(_0211_),
    .CLK(clknet_leaf_9_clock),
    .Q(\u1.row_sel[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3071_ (.D(_0212_),
    .CLK(clknet_leaf_9_clock),
    .Q(\u1.row_sel[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3072_ (.D(_0213_),
    .CLK(clknet_leaf_10_clock),
    .Q(\u1.row_sel[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3073_ (.D(_0214_),
    .CLK(clknet_leaf_10_clock),
    .Q(\u1.row_sel[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3074_ (.D(_0215_),
    .CLK(clknet_leaf_10_clock),
    .Q(\u1.row_sel[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3075_ (.D(_0216_),
    .CLK(clknet_leaf_11_clock),
    .Q(\u1.row_sel[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3076_ (.D(_0217_),
    .CLK(clknet_leaf_5_clock),
    .Q(\u0.u11.impulse_gen[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3077_ (.D(_0218_),
    .CLK(clknet_leaf_4_clock),
    .Q(\u0.u11.impulse_gen[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3078_ (.D(_0006_),
    .CLK(clknet_leaf_9_clock),
    .Q(\u0.run_state[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3079_ (.D(_0004_),
    .CLK(clknet_leaf_12_clock),
    .Q(\u0.run_state[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3080_ (.D(_0005_),
    .CLK(clknet_leaf_12_clock),
    .Q(\u0.run_state[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3081_ (.D(_0007_),
    .CLK(clknet_leaf_4_clock),
    .Q(\u0.run_state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3082_ (.D(_0008_),
    .CLK(clknet_leaf_4_clock),
    .Q(\u0.run_state[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3083_ (.D(_0009_),
    .CLK(clknet_leaf_4_clock),
    .Q(\u0.run_state[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3084_ (.D(_0010_),
    .CLK(clknet_leaf_4_clock),
    .Q(\u0.run_state[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3085_ (.D(_0219_),
    .CLK(clknet_leaf_35_clock),
    .Q(net149));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3086_ (.D(_0220_),
    .CLK(clknet_leaf_29_clock),
    .Q(\u1.timer[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3087_ (.D(_0221_),
    .CLK(clknet_leaf_29_clock),
    .Q(\u1.timer[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3088_ (.D(_0222_),
    .CLK(clknet_leaf_29_clock),
    .Q(\u1.timer[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3089_ (.D(_0223_),
    .CLK(clknet_leaf_29_clock),
    .Q(\u1.timer[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3090_ (.D(_0224_),
    .CLK(clknet_leaf_23_clock),
    .Q(\u1.timer[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3091_ (.D(_0225_),
    .CLK(clknet_leaf_25_clock),
    .Q(\u1.timer[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3092_ (.D(_0226_),
    .CLK(clknet_leaf_25_clock),
    .Q(\u1.timer[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3093_ (.D(_0227_),
    .CLK(clknet_leaf_26_clock),
    .Q(\u1.timer[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3094_ (.D(_0228_),
    .CLK(clknet_leaf_26_clock),
    .Q(\u1.timer[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3095_ (.D(_0229_),
    .CLK(clknet_leaf_26_clock),
    .Q(\u1.timer[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3096_ (.D(_0230_),
    .CLK(clknet_leaf_27_clock),
    .Q(\u1.timer[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3097_ (.D(_0231_),
    .CLK(clknet_leaf_26_clock),
    .Q(\u1.timer[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3098_ (.D(_0232_),
    .CLK(clknet_leaf_27_clock),
    .Q(\u1.timer[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3099_ (.D(_0233_),
    .CLK(clknet_leaf_29_clock),
    .Q(\u1.timer[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3100_ (.D(_0234_),
    .CLK(clknet_leaf_29_clock),
    .Q(\u1.timer[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3101_ (.D(_0235_),
    .CLK(clknet_leaf_28_clock),
    .Q(\u1.timer[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3102_ (.D(_0236_),
    .CLK(clknet_leaf_28_clock),
    .Q(\u1.timer[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3103_ (.D(_0237_),
    .CLK(clknet_leaf_32_clock),
    .Q(\u1.timer[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3104_ (.D(_0238_),
    .CLK(clknet_leaf_30_clock),
    .Q(\u1.timer[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3105_ (.D(_0239_),
    .CLK(clknet_leaf_31_clock),
    .Q(\u1.timer[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3106_ (.D(_0240_),
    .CLK(clknet_leaf_31_clock),
    .Q(\u1.timer[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3107_ (.D(_0241_),
    .CLK(clknet_leaf_31_clock),
    .Q(\u1.timer[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3108_ (.D(_0242_),
    .CLK(clknet_leaf_31_clock),
    .Q(\u1.timer[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3109_ (.D(_0243_),
    .CLK(clknet_leaf_31_clock),
    .Q(\u1.timer[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3110_ (.D(_0244_),
    .CLK(clknet_leaf_33_clock),
    .Q(\u1.timer[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3111_ (.D(_0245_),
    .CLK(clknet_leaf_34_clock),
    .Q(\u1.timer[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3112_ (.D(_0246_),
    .CLK(clknet_leaf_34_clock),
    .Q(\u1.timer[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3113_ (.D(_0247_),
    .CLK(clknet_leaf_34_clock),
    .Q(\u1.timer[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3114_ (.D(_0248_),
    .CLK(clknet_leaf_36_clock),
    .Q(\u1.timer[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3115_ (.D(_0249_),
    .CLK(clknet_leaf_36_clock),
    .Q(\u1.timer[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3116_ (.D(_0250_),
    .CLK(clknet_leaf_36_clock),
    .Q(\u1.timer[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3117_ (.D(_0251_),
    .CLK(clknet_leaf_36_clock),
    .Q(\u1.timer[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3118_ (.D(net40),
    .CLK(net227),
    .Q(\spi_data_crossing[0].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3119_ (.D(\spi_data_crossing[0].A ),
    .CLK(clknet_leaf_35_clock),
    .Q(\spi_data_crossing[0].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3120_ (.D(net51),
    .CLK(net229),
    .Q(\spi_data_crossing[1].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3121_ (.D(\spi_data_crossing[1].A ),
    .CLK(clknet_leaf_35_clock),
    .Q(\spi_data_crossing[1].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3122_ (.D(net62),
    .CLK(net229),
    .Q(\spi_data_crossing[2].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3123_ (.D(\spi_data_crossing[2].A ),
    .CLK(clknet_leaf_36_clock),
    .Q(\spi_data_crossing[2].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3124_ (.D(net65),
    .CLK(net227),
    .Q(\spi_data_crossing[3].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3125_ (.D(\spi_data_crossing[3].A ),
    .CLK(clknet_leaf_36_clock),
    .Q(\spi_data_crossing[3].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3126_ (.D(net66),
    .CLK(net227),
    .Q(\spi_data_crossing[4].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3127_ (.D(\spi_data_crossing[4].A ),
    .CLK(clknet_leaf_36_clock),
    .Q(\spi_data_crossing[4].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3128_ (.D(net67),
    .CLK(net227),
    .Q(\spi_data_crossing[5].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3129_ (.D(\spi_data_crossing[5].A ),
    .CLK(clknet_leaf_0_clock),
    .Q(\spi_data_crossing[5].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3130_ (.D(net68),
    .CLK(net228),
    .Q(\spi_data_crossing[6].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3131_ (.D(\spi_data_crossing[6].A ),
    .CLK(clknet_leaf_0_clock),
    .Q(\spi_data_crossing[6].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3132_ (.D(net69),
    .CLK(net228),
    .Q(\spi_data_crossing[7].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3133_ (.D(\spi_data_crossing[7].A ),
    .CLK(clknet_leaf_5_clock),
    .Q(\spi_data_crossing[7].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3134_ (.D(net70),
    .CLK(net230),
    .Q(\spi_data_crossing[8].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3135_ (.D(\spi_data_crossing[8].A ),
    .CLK(clknet_leaf_0_clock),
    .Q(\spi_data_crossing[8].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3136_ (.D(net71),
    .CLK(net230),
    .Q(\spi_data_crossing[9].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3137_ (.D(\spi_data_crossing[9].A ),
    .CLK(clknet_leaf_0_clock),
    .Q(\spi_data_crossing[9].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3138_ (.D(net41),
    .CLK(net230),
    .Q(\spi_data_crossing[10].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3139_ (.D(\spi_data_crossing[10].A ),
    .CLK(clknet_leaf_0_clock),
    .Q(\spi_data_crossing[10].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3140_ (.D(net42),
    .CLK(net230),
    .Q(\spi_data_crossing[11].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3141_ (.D(\spi_data_crossing[11].A ),
    .CLK(clknet_leaf_0_clock),
    .Q(\spi_data_crossing[11].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3142_ (.D(net43),
    .CLK(net231),
    .Q(\spi_data_crossing[12].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3143_ (.D(\spi_data_crossing[12].A ),
    .CLK(clknet_leaf_0_clock),
    .Q(\spi_data_crossing[12].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3144_ (.D(net44),
    .CLK(net231),
    .Q(\spi_data_crossing[13].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3145_ (.D(\spi_data_crossing[13].A ),
    .CLK(clknet_leaf_1_clock),
    .Q(\spi_data_crossing[13].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3146_ (.D(net45),
    .CLK(net234),
    .Q(\spi_data_crossing[14].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3147_ (.D(\spi_data_crossing[14].A ),
    .CLK(clknet_leaf_1_clock),
    .Q(\spi_data_crossing[14].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3148_ (.D(net46),
    .CLK(net234),
    .Q(\spi_data_crossing[15].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3149_ (.D(\spi_data_crossing[15].A ),
    .CLK(clknet_leaf_1_clock),
    .Q(\spi_data_crossing[15].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3150_ (.D(net47),
    .CLK(net234),
    .Q(\spi_data_crossing[16].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3151_ (.D(\spi_data_crossing[16].A ),
    .CLK(clknet_leaf_5_clock),
    .Q(\spi_data_crossing[16].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3152_ (.D(net48),
    .CLK(net234),
    .Q(\spi_data_crossing[17].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3153_ (.D(\spi_data_crossing[17].A ),
    .CLK(clknet_leaf_5_clock),
    .Q(\spi_data_crossing[17].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3154_ (.D(net49),
    .CLK(net235),
    .Q(\spi_data_crossing[18].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3155_ (.D(\spi_data_crossing[18].A ),
    .CLK(clknet_leaf_5_clock),
    .Q(\spi_data_crossing[18].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3156_ (.D(net50),
    .CLK(net235),
    .Q(\spi_data_crossing[19].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3157_ (.D(\spi_data_crossing[19].A ),
    .CLK(clknet_leaf_5_clock),
    .Q(\spi_data_crossing[19].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3158_ (.D(net52),
    .CLK(net235),
    .Q(\spi_data_crossing[20].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3159_ (.D(\spi_data_crossing[20].A ),
    .CLK(clknet_leaf_6_clock),
    .Q(\spi_data_crossing[20].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3160_ (.D(net53),
    .CLK(net239),
    .Q(\spi_data_crossing[21].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3161_ (.D(\spi_data_crossing[21].A ),
    .CLK(clknet_leaf_6_clock),
    .Q(\spi_data_crossing[21].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3162_ (.D(net54),
    .CLK(net239),
    .Q(\spi_data_crossing[22].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3163_ (.D(\spi_data_crossing[22].A ),
    .CLK(clknet_leaf_6_clock),
    .Q(\spi_data_crossing[22].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3164_ (.D(net55),
    .CLK(net239),
    .Q(\spi_data_crossing[23].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3165_ (.D(\spi_data_crossing[23].A ),
    .CLK(clknet_leaf_6_clock),
    .Q(\spi_data_crossing[23].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3166_ (.D(net56),
    .CLK(net237),
    .Q(\spi_data_crossing[24].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3167_ (.D(\spi_data_crossing[24].A ),
    .CLK(clknet_leaf_7_clock),
    .Q(\spi_data_crossing[24].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3168_ (.D(net57),
    .CLK(net237),
    .Q(\spi_data_crossing[25].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3169_ (.D(\spi_data_crossing[25].A ),
    .CLK(clknet_leaf_7_clock),
    .Q(\spi_data_crossing[25].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3170_ (.D(net58),
    .CLK(net237),
    .Q(\spi_data_crossing[26].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3171_ (.D(\spi_data_crossing[26].A ),
    .CLK(clknet_leaf_7_clock),
    .Q(\spi_data_crossing[26].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3172_ (.D(net59),
    .CLK(net240),
    .Q(\spi_data_crossing[27].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3173_ (.D(\spi_data_crossing[27].A ),
    .CLK(clknet_leaf_7_clock),
    .Q(\spi_data_crossing[27].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3174_ (.D(net60),
    .CLK(net240),
    .Q(\spi_data_crossing[28].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3175_ (.D(\spi_data_crossing[28].A ),
    .CLK(clknet_leaf_7_clock),
    .Q(\spi_data_crossing[28].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3176_ (.D(net61),
    .CLK(net238),
    .Q(\spi_data_crossing[29].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3177_ (.D(\spi_data_crossing[29].A ),
    .CLK(clknet_leaf_7_clock),
    .Q(\spi_data_crossing[29].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3178_ (.D(net63),
    .CLK(net237),
    .Q(\spi_data_crossing[30].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3179_ (.D(\spi_data_crossing[30].A ),
    .CLK(clknet_leaf_6_clock),
    .Q(\spi_data_crossing[30].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3180_ (.D(net64),
    .CLK(net240),
    .Q(\spi_data_crossing[31].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3181_ (.D(\spi_data_crossing[31].A ),
    .CLK(clknet_leaf_7_clock),
    .Q(\spi_data_crossing[31].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3182_ (.D(_0252_),
    .CLK(clknet_leaf_32_clock),
    .Q(net148));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3183_ (.D(_0253_),
    .CLK(clknet_leaf_28_clock),
    .Q(net146));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3184_ (.D(_0254_),
    .CLK(clknet_leaf_33_clock),
    .Q(net144));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3185_ (.D(_0255_),
    .CLK(clknet_leaf_33_clock),
    .Q(net142));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3186_ (.D(_0256_),
    .CLK(clknet_leaf_33_clock),
    .Q(net140));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3187_ (.D(_0257_),
    .CLK(clknet_leaf_33_clock),
    .Q(net157));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3188_ (.D(_0258_),
    .CLK(clknet_leaf_33_clock),
    .Q(net155));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3189_ (.D(_0259_),
    .CLK(clknet_leaf_35_clock),
    .Q(net153));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3190_ (.D(_0260_),
    .CLK(clknet_leaf_35_clock),
    .Q(net151));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3191_ (.D(_0261_),
    .CLK(clknet_leaf_23_clock),
    .Q(\u1.ccr0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3192_ (.D(_0262_),
    .CLK(clknet_leaf_30_clock),
    .Q(\u1.ccr0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3193_ (.D(_0263_),
    .CLK(clknet_leaf_30_clock),
    .Q(\u1.ccr0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3194_ (.D(_0264_),
    .CLK(clknet_leaf_30_clock),
    .Q(\u1.ccr0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3195_ (.D(_0265_),
    .CLK(clknet_leaf_23_clock),
    .Q(\u1.ccr0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3196_ (.D(_0266_),
    .CLK(clknet_leaf_24_clock),
    .Q(\u1.ccr0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3197_ (.D(_0267_),
    .CLK(clknet_leaf_23_clock),
    .Q(\u1.ccr0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3198_ (.D(_0268_),
    .CLK(clknet_leaf_23_clock),
    .Q(\u1.ccr0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3199_ (.D(_0269_),
    .CLK(clknet_leaf_31_clock),
    .Q(\u1.ccr0[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3200_ (.D(_0270_),
    .CLK(clknet_leaf_31_clock),
    .Q(\u1.ccr0[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3201_ (.D(_0271_),
    .CLK(clknet_leaf_23_clock),
    .Q(\u1.ccr0[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3202_ (.D(_0272_),
    .CLK(clknet_leaf_23_clock),
    .Q(\u1.ccr0[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3203_ (.D(_0273_),
    .CLK(clknet_leaf_23_clock),
    .Q(\u1.ccr0[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3204_ (.D(_0274_),
    .CLK(clknet_leaf_23_clock),
    .Q(\u1.ccr0[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3205_ (.D(_0275_),
    .CLK(clknet_leaf_23_clock),
    .Q(\u1.ccr0[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3206_ (.D(_0276_),
    .CLK(clknet_leaf_29_clock),
    .Q(\u1.ccr0[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3207_ (.D(_0277_),
    .CLK(clknet_leaf_35_clock),
    .Q(net159));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3208_ (.D(_0278_),
    .CLK(clknet_leaf_35_clock),
    .Q(net158));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3209_ (.D(_0001_),
    .CLK(clknet_leaf_28_clock),
    .Q(net161));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3210_ (.D(_0279_),
    .CLK(clknet_leaf_35_clock),
    .Q(net137));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3211_ (.D(_0003_),
    .CLK(clknet_leaf_33_clock),
    .Q(reset_n));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3212_ (.D(_0002_),
    .CLK(clknet_leaf_34_clock),
    .Q(latch_data));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3213_ (.D(_0000_),
    .CLK(clknet_leaf_32_clock),
    .Q(control_trigger));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3214_ (.D(net267),
    .CLK(clknet_leaf_17_clock),
    .Q(net127));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3215_ (.D(net277),
    .CLK(clknet_leaf_17_clock),
    .Q(net128));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3216_ (.D(net275),
    .CLK(clknet_leaf_17_clock),
    .Q(net129));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3217_ (.D(net253),
    .CLK(clknet_leaf_16_clock),
    .Q(net130));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3218_ (.D(net262),
    .CLK(clknet_leaf_17_clock),
    .Q(net131));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3219_ (.D(net261),
    .CLK(clknet_leaf_17_clock),
    .Q(net132));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3220_ (.D(net281),
    .CLK(clknet_leaf_17_clock),
    .Q(net133));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3221_ (.D(net282),
    .CLK(clknet_leaf_17_clock),
    .Q(net134));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3222_ (.D(net278),
    .CLK(clknet_leaf_18_clock),
    .Q(net135));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3223_ (.D(net265),
    .CLK(clknet_leaf_17_clock),
    .Q(net136));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3224_ (.D(net287),
    .CLK(clknet_leaf_16_clock),
    .Q(net194));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3225_ (.D(net273),
    .CLK(clknet_leaf_17_clock),
    .Q(net195));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3226_ (.D(net283),
    .CLK(clknet_leaf_16_clock),
    .Q(net196));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3227_ (.D(net274),
    .CLK(clknet_leaf_17_clock),
    .Q(net197));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3228_ (.D(net263),
    .CLK(clknet_leaf_17_clock),
    .Q(net198));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3229_ (.D(net280),
    .CLK(clknet_leaf_18_clock),
    .Q(net199));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3230_ (.D(net264),
    .CLK(clknet_leaf_17_clock),
    .Q(net200));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3231_ (.D(net284),
    .CLK(clknet_leaf_17_clock),
    .Q(net201));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3232_ (.D(net266),
    .CLK(clknet_leaf_17_clock),
    .Q(net202));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3233_ (.D(net260),
    .CLK(clknet_leaf_17_clock),
    .Q(net203));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3234_ (.D(\u0.cmd[16] ),
    .CLK(clknet_leaf_7_clock),
    .Q(net162));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3235_ (.D(net269),
    .CLK(clknet_leaf_7_clock),
    .Q(net163));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3236_ (.D(\u0.cmd[18] ),
    .CLK(clknet_leaf_7_clock),
    .Q(net164));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3237_ (.D(net218),
    .CLK(clknet_leaf_7_clock),
    .Q(net165));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3238_ (.D(\u0.cmd[20] ),
    .CLK(clknet_leaf_7_clock),
    .Q(net166));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3239_ (.D(\u0.cmd[21] ),
    .CLK(clknet_leaf_7_clock),
    .Q(net167));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3240_ (.D(net258),
    .CLK(clknet_leaf_7_clock),
    .Q(net168));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3241_ (.D(net254),
    .CLK(clknet_leaf_7_clock),
    .Q(net169));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3242_ (.D(net285),
    .CLK(clknet_leaf_7_clock),
    .Q(net170));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3243_ (.D(net286),
    .CLK(clknet_leaf_7_clock),
    .Q(net171));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3244_ (.D(net252),
    .CLK(clknet_leaf_8_clock),
    .Q(net182));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3245_ (.D(net251),
    .CLK(clknet_leaf_8_clock),
    .Q(net183));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3246_ (.D(net256),
    .CLK(clknet_leaf_8_clock),
    .Q(net184));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3247_ (.D(net255),
    .CLK(clknet_leaf_8_clock),
    .Q(net185));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3248_ (.D(net247),
    .CLK(clknet_leaf_9_clock),
    .Q(net186));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3249_ (.D(net248),
    .CLK(clknet_leaf_10_clock),
    .Q(net187));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3250_ (.D(net257),
    .CLK(clknet_leaf_8_clock),
    .Q(net188));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3251_ (.D(net245),
    .CLK(clknet_leaf_9_clock),
    .Q(net189));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3252_ (.D(net246),
    .CLK(clknet_leaf_9_clock),
    .Q(net190));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3253_ (.D(net244),
    .CLK(clknet_leaf_9_clock),
    .Q(net191));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3254_ (.I(clknet_leaf_9_clock),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3255_ (.I(clknet_leaf_9_clock),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3256_ (.I(clknet_leaf_9_clock),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3257_ (.I(clknet_leaf_9_clock),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3258_ (.I(clknet_leaf_9_clock),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3259_ (.I(clknet_leaf_10_clock),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3260_ (.I(clknet_leaf_10_clock),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3261_ (.I(clknet_leaf_10_clock),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3262_ (.I(clknet_leaf_10_clock),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3263_ (.I(clknet_leaf_10_clock),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3264_ (.I(net83),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3265_ (.I(net84),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3266_ (.I(net85),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3267_ (.I(net86),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3268_ (.I(net87),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3269_ (.I(net88),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3270_ (.I(net95),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3271_ (.I(net102),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3272_ (.I(net103),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3273_ (.I(net104),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3274_ (.I(net105),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3275_ (.I(net106),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3276_ (.I(net107),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3277_ (.I(net108),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3278_ (.I(net109),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3279_ (.I(net110),
    .Z(net126));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3280_ (.I(net96),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3281_ (.I(net97),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3282_ (.I(net98),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3283_ (.I(net99),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3284_ (.I(net100),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3285_ (.I(net101),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3286_ (.I(net149),
    .Z(net138));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3287_ (.I(net151),
    .Z(net150));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3288_ (.I(net153),
    .Z(net152));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3289_ (.I(net155),
    .Z(net154));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3290_ (.I(net157),
    .Z(net156));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3291_ (.I(net140),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3292_ (.I(net142),
    .Z(net141));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3293_ (.I(net144),
    .Z(net143));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3294_ (.I(net146),
    .Z(net145));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3295_ (.I(net148),
    .Z(net147));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3296_ (.I(net162),
    .Z(net172));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3297_ (.I(net163),
    .Z(net173));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3298_ (.I(net164),
    .Z(net174));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3299_ (.I(net165),
    .Z(net175));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3300_ (.I(net166),
    .Z(net176));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3301_ (.I(net167),
    .Z(net177));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3302_ (.I(net168),
    .Z(net178));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3303_ (.I(net169),
    .Z(net179));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3304_ (.I(net170),
    .Z(net180));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3305_ (.I(net171),
    .Z(net181));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3306_ (.I(net192),
    .Z(net193));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3307_ (.I(net204),
    .Z(net210));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3308_ (.I(net205),
    .Z(net211));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3309_ (.I(net206),
    .Z(net212));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3310_ (.I(net207),
    .Z(net213));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3311_ (.I(net208),
    .Z(net214));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3312_ (.I(net209),
    .Z(net215));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input1 (.I(io_control_trigger_in),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input2 (.I(io_latch_data_in),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input3 (.I(io_reset_n_in),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input4 (.I(la_data_in[0]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input5 (.I(la_data_in[10]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input6 (.I(la_data_in[11]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input7 (.I(la_data_in[12]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input8 (.I(la_data_in[13]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input9 (.I(la_data_in[14]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input10 (.I(la_data_in[15]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input11 (.I(la_data_in[16]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input12 (.I(la_data_in[17]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input13 (.I(la_data_in[1]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input14 (.I(la_data_in[2]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input15 (.I(la_data_in[3]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input16 (.I(la_data_in[4]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input17 (.I(la_data_in[5]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input18 (.I(la_data_in[6]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input19 (.I(la_data_in[7]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input20 (.I(la_data_in[8]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input21 (.I(la_data_in[9]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input22 (.I(la_oenb[0]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input23 (.I(la_oenb[10]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input24 (.I(la_oenb[11]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input25 (.I(la_oenb[12]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input26 (.I(la_oenb[13]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input27 (.I(la_oenb[14]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input28 (.I(la_oenb[15]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input29 (.I(la_oenb[16]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input30 (.I(la_oenb[17]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input31 (.I(la_oenb[1]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input32 (.I(la_oenb[2]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input33 (.I(la_oenb[3]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input34 (.I(la_oenb[4]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input35 (.I(la_oenb[5]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input36 (.I(la_oenb[6]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input37 (.I(la_oenb[7]),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input38 (.I(la_oenb[8]),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input39 (.I(la_oenb[9]),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input40 (.I(spi_data[0]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input41 (.I(spi_data[10]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input42 (.I(spi_data[11]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input43 (.I(spi_data[12]),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input44 (.I(spi_data[13]),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input45 (.I(spi_data[14]),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input46 (.I(spi_data[15]),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input47 (.I(spi_data[16]),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input48 (.I(spi_data[17]),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input49 (.I(spi_data[18]),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input50 (.I(spi_data[19]),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input51 (.I(spi_data[1]),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input52 (.I(spi_data[20]),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input53 (.I(spi_data[21]),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input54 (.I(spi_data[22]),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input55 (.I(spi_data[23]),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input56 (.I(spi_data[24]),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input57 (.I(spi_data[25]),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input58 (.I(spi_data[26]),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input59 (.I(spi_data[27]),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input60 (.I(spi_data[28]),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input61 (.I(spi_data[29]),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input62 (.I(spi_data[2]),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input63 (.I(spi_data[30]),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input64 (.I(spi_data[31]),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input65 (.I(spi_data[3]),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input66 (.I(spi_data[4]),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input67 (.I(spi_data[5]),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input68 (.I(spi_data[6]),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input69 (.I(spi_data[7]),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input70 (.I(spi_data[8]),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input71 (.I(spi_data[9]),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input72 (.I(spi_data_clock),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 output73 (.I(net73),
    .Z(clock_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 output74 (.I(net74),
    .Z(clock_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 output75 (.I(net75),
    .Z(clock_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 output76 (.I(net76),
    .Z(clock_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 output77 (.I(net77),
    .Z(clock_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 output78 (.I(net78),
    .Z(clock_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 output79 (.I(net79),
    .Z(clock_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 output80 (.I(net80),
    .Z(clock_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 output81 (.I(net81),
    .Z(clock_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 output82 (.I(net82),
    .Z(clock_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output83 (.I(net83),
    .Z(col_select_left[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output84 (.I(net84),
    .Z(col_select_left[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output85 (.I(net85),
    .Z(col_select_left[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output86 (.I(net86),
    .Z(col_select_left[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output87 (.I(net87),
    .Z(col_select_left[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output88 (.I(net88),
    .Z(col_select_left[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output89 (.I(net89),
    .Z(col_select_right[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output90 (.I(net90),
    .Z(col_select_right[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output91 (.I(net91),
    .Z(col_select_right[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output92 (.I(net92),
    .Z(col_select_right[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output93 (.I(net93),
    .Z(col_select_right[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output94 (.I(net94),
    .Z(col_select_right[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output95 (.I(net95),
    .Z(data_out_left[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output96 (.I(net96),
    .Z(data_out_left[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output97 (.I(net97),
    .Z(data_out_left[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output98 (.I(net98),
    .Z(data_out_left[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output99 (.I(net99),
    .Z(data_out_left[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output100 (.I(net100),
    .Z(data_out_left[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output101 (.I(net101),
    .Z(data_out_left[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output102 (.I(net102),
    .Z(data_out_left[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output103 (.I(net103),
    .Z(data_out_left[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output104 (.I(net104),
    .Z(data_out_left[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output105 (.I(net105),
    .Z(data_out_left[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output106 (.I(net106),
    .Z(data_out_left[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output107 (.I(net107),
    .Z(data_out_left[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output108 (.I(net108),
    .Z(data_out_left[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output109 (.I(net109),
    .Z(data_out_left[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output110 (.I(net110),
    .Z(data_out_left[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output111 (.I(net111),
    .Z(data_out_right[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output112 (.I(net112),
    .Z(data_out_right[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output113 (.I(net113),
    .Z(data_out_right[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output114 (.I(net114),
    .Z(data_out_right[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output115 (.I(net115),
    .Z(data_out_right[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output116 (.I(net116),
    .Z(data_out_right[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output117 (.I(net117),
    .Z(data_out_right[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output118 (.I(net118),
    .Z(data_out_right[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output119 (.I(net119),
    .Z(data_out_right[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output120 (.I(net120),
    .Z(data_out_right[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output121 (.I(net121),
    .Z(data_out_right[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output122 (.I(net122),
    .Z(data_out_right[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output123 (.I(net123),
    .Z(data_out_right[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output124 (.I(net124),
    .Z(data_out_right[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output125 (.I(net125),
    .Z(data_out_right[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output126 (.I(net126),
    .Z(data_out_right[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output127 (.I(net127),
    .Z(inverter_select[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output128 (.I(net128),
    .Z(inverter_select[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output129 (.I(net129),
    .Z(inverter_select[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output130 (.I(net130),
    .Z(inverter_select[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output131 (.I(net131),
    .Z(inverter_select[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output132 (.I(net132),
    .Z(inverter_select[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output133 (.I(net133),
    .Z(inverter_select[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output134 (.I(net134),
    .Z(inverter_select[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output135 (.I(net135),
    .Z(inverter_select[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output136 (.I(net136),
    .Z(inverter_select[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output137 (.I(net137),
    .Z(io_control_trigger_oeb));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output138 (.I(net138),
    .Z(io_driver_io_oeb[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output139 (.I(net139),
    .Z(io_driver_io_oeb[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output140 (.I(net140),
    .Z(io_driver_io_oeb[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output141 (.I(net141),
    .Z(io_driver_io_oeb[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output142 (.I(net142),
    .Z(io_driver_io_oeb[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output143 (.I(net143),
    .Z(io_driver_io_oeb[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output144 (.I(net144),
    .Z(io_driver_io_oeb[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output145 (.I(net145),
    .Z(io_driver_io_oeb[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output146 (.I(net146),
    .Z(io_driver_io_oeb[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output147 (.I(net147),
    .Z(io_driver_io_oeb[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output148 (.I(net148),
    .Z(io_driver_io_oeb[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output149 (.I(net149),
    .Z(io_driver_io_oeb[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output150 (.I(net150),
    .Z(io_driver_io_oeb[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output151 (.I(net151),
    .Z(io_driver_io_oeb[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output152 (.I(net152),
    .Z(io_driver_io_oeb[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output153 (.I(net153),
    .Z(io_driver_io_oeb[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output154 (.I(net154),
    .Z(io_driver_io_oeb[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output155 (.I(net155),
    .Z(io_driver_io_oeb[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output156 (.I(net156),
    .Z(io_driver_io_oeb[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output157 (.I(net157),
    .Z(io_driver_io_oeb[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output158 (.I(net158),
    .Z(io_latch_data_oeb));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output159 (.I(net159),
    .Z(io_reset_n_oeb));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output160 (.I(net160),
    .Z(io_update_cycle_complete_oeb));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output161 (.I(net161),
    .Z(io_update_cycle_complete_out));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output162 (.I(net162),
    .Z(mem_address_left[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output163 (.I(net163),
    .Z(mem_address_left[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output164 (.I(net164),
    .Z(mem_address_left[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output165 (.I(net165),
    .Z(mem_address_left[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output166 (.I(net166),
    .Z(mem_address_left[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output167 (.I(net167),
    .Z(mem_address_left[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output168 (.I(net168),
    .Z(mem_address_left[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output169 (.I(net169),
    .Z(mem_address_left[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output170 (.I(net170),
    .Z(mem_address_left[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output171 (.I(net171),
    .Z(mem_address_left[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output172 (.I(net172),
    .Z(mem_address_right[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output173 (.I(net173),
    .Z(mem_address_right[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output174 (.I(net174),
    .Z(mem_address_right[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output175 (.I(net175),
    .Z(mem_address_right[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output176 (.I(net176),
    .Z(mem_address_right[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output177 (.I(net177),
    .Z(mem_address_right[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output178 (.I(net178),
    .Z(mem_address_right[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output179 (.I(net179),
    .Z(mem_address_right[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output180 (.I(net180),
    .Z(mem_address_right[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output181 (.I(net181),
    .Z(mem_address_right[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output182 (.I(net182),
    .Z(mem_write_n[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output183 (.I(net183),
    .Z(mem_write_n[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output184 (.I(net184),
    .Z(mem_write_n[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output185 (.I(net185),
    .Z(mem_write_n[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output186 (.I(net186),
    .Z(mem_write_n[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output187 (.I(net187),
    .Z(mem_write_n[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output188 (.I(net188),
    .Z(mem_write_n[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output189 (.I(net189),
    .Z(mem_write_n[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output190 (.I(net190),
    .Z(mem_write_n[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output191 (.I(net191),
    .Z(mem_write_n[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output192 (.I(net192),
    .Z(output_active_left));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output193 (.I(net193),
    .Z(output_active_right));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output194 (.I(net194),
    .Z(row_col_select[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output195 (.I(net195),
    .Z(row_col_select[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output196 (.I(net196),
    .Z(row_col_select[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output197 (.I(net197),
    .Z(row_col_select[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output198 (.I(net198),
    .Z(row_col_select[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output199 (.I(net199),
    .Z(row_col_select[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output200 (.I(net200),
    .Z(row_col_select[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output201 (.I(net201),
    .Z(row_col_select[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output202 (.I(net202),
    .Z(row_col_select[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output203 (.I(net203),
    .Z(row_col_select[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output204 (.I(net204),
    .Z(row_select_left[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output205 (.I(net205),
    .Z(row_select_left[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output206 (.I(net206),
    .Z(row_select_left[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output207 (.I(net207),
    .Z(row_select_left[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output208 (.I(net208),
    .Z(row_select_left[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output209 (.I(net209),
    .Z(row_select_left[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output210 (.I(net210),
    .Z(row_select_right[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output211 (.I(net211),
    .Z(row_select_right[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output212 (.I(net212),
    .Z(row_select_right[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output213 (.I(net213),
    .Z(row_select_right[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output214 (.I(net214),
    .Z(row_select_right[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output215 (.I(net215),
    .Z(row_select_right[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout216 (.I(\u1.row_sel[5] ),
    .Z(net216));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout217 (.I(\u1.row_sel[4] ),
    .Z(net217));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout218 (.I(\u0.cmd[19] ),
    .Z(net218));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout219 (.I(\u0.cmd[15] ),
    .Z(net219));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout220 (.I(\u0.cmd[14] ),
    .Z(net220));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout221 (.I(\u0.cmd[13] ),
    .Z(net221));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout222 (.I(\u0.cmd[12] ),
    .Z(net222));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout223 (.I(\u0.cmd[11] ),
    .Z(net223));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout224 (.I(\u0.cmd[10] ),
    .Z(net224));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout225 (.I(\u1.col_sel[2] ),
    .Z(net225));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout226 (.I(\u1.col_sel[0] ),
    .Z(net226));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout227 (.I(net229),
    .Z(net227));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout228 (.I(net229),
    .Z(net228));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout229 (.I(net233),
    .Z(net229));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout230 (.I(net232),
    .Z(net230));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout231 (.I(net232),
    .Z(net231));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout232 (.I(net233),
    .Z(net232));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout233 (.I(net242),
    .Z(net233));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout234 (.I(net236),
    .Z(net234));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout235 (.I(net236),
    .Z(net235));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout236 (.I(net241),
    .Z(net236));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout237 (.I(net238),
    .Z(net237));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout238 (.I(net239),
    .Z(net238));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout239 (.I(net240),
    .Z(net239));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout240 (.I(net241),
    .Z(net240));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout241 (.I(net242),
    .Z(net241));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout242 (.I(net72),
    .Z(net242));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_0_clock (.I(clknet_2_0__leaf_clock),
    .Z(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_clock (.I(clknet_2_0__leaf_clock),
    .Z(clknet_leaf_1_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_clock (.I(clknet_2_0__leaf_clock),
    .Z(clknet_leaf_2_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_3_clock (.I(clknet_2_1__leaf_clock),
    .Z(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_4_clock (.I(clknet_2_1__leaf_clock),
    .Z(clknet_leaf_4_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_5_clock (.I(clknet_2_1__leaf_clock),
    .Z(clknet_leaf_5_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_6_clock (.I(clknet_2_1__leaf_clock),
    .Z(clknet_leaf_6_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_7_clock (.I(clknet_2_1__leaf_clock),
    .Z(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_8_clock (.I(clknet_2_1__leaf_clock),
    .Z(clknet_leaf_8_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_9_clock (.I(clknet_2_1__leaf_clock),
    .Z(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_10_clock (.I(clknet_2_1__leaf_clock),
    .Z(clknet_leaf_10_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_11_clock (.I(clknet_2_1__leaf_clock),
    .Z(clknet_leaf_11_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_12_clock (.I(clknet_2_1__leaf_clock),
    .Z(clknet_leaf_12_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_13_clock (.I(clknet_2_1__leaf_clock),
    .Z(clknet_leaf_13_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_14_clock (.I(clknet_2_3__leaf_clock),
    .Z(clknet_leaf_14_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_clock (.I(clknet_2_3__leaf_clock),
    .Z(clknet_leaf_15_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_16_clock (.I(clknet_2_3__leaf_clock),
    .Z(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_17_clock (.I(clknet_2_3__leaf_clock),
    .Z(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_18_clock (.I(clknet_2_3__leaf_clock),
    .Z(clknet_leaf_18_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_19_clock (.I(clknet_2_3__leaf_clock),
    .Z(clknet_leaf_19_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_20_clock (.I(clknet_2_3__leaf_clock),
    .Z(clknet_leaf_20_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_21_clock (.I(clknet_2_3__leaf_clock),
    .Z(clknet_leaf_21_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_22_clock (.I(clknet_2_2__leaf_clock),
    .Z(clknet_leaf_22_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_23_clock (.I(clknet_2_2__leaf_clock),
    .Z(clknet_leaf_23_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_24_clock (.I(clknet_2_2__leaf_clock),
    .Z(clknet_leaf_24_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_25_clock (.I(clknet_2_2__leaf_clock),
    .Z(clknet_leaf_25_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_26_clock (.I(clknet_2_2__leaf_clock),
    .Z(clknet_leaf_26_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_27_clock (.I(clknet_2_2__leaf_clock),
    .Z(clknet_leaf_27_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_28_clock (.I(clknet_2_2__leaf_clock),
    .Z(clknet_leaf_28_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_29_clock (.I(clknet_2_2__leaf_clock),
    .Z(clknet_leaf_29_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_30_clock (.I(clknet_2_0__leaf_clock),
    .Z(clknet_leaf_30_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_31_clock (.I(clknet_2_0__leaf_clock),
    .Z(clknet_leaf_31_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_32_clock (.I(clknet_2_0__leaf_clock),
    .Z(clknet_leaf_32_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_33_clock (.I(clknet_2_0__leaf_clock),
    .Z(clknet_leaf_33_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_34_clock (.I(clknet_2_0__leaf_clock),
    .Z(clknet_leaf_34_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_35_clock (.I(clknet_2_0__leaf_clock),
    .Z(clknet_leaf_35_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_36_clock (.I(clknet_2_0__leaf_clock),
    .Z(clknet_leaf_36_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_clock (.I(clock),
    .Z(clknet_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_0__f_clock (.I(clknet_0_clock),
    .Z(clknet_2_0__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_1__f_clock (.I(clknet_0_clock),
    .Z(clknet_2_1__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_2__f_clock (.I(clknet_0_clock),
    .Z(clknet_2_2__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_3__f_clock (.I(clknet_0_clock),
    .Z(clknet_2_3__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold1 (.I(latch_data),
    .Z(net243));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold2 (.I(\u0.mem_write_n[9] ),
    .Z(net244));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold3 (.I(\u0.mem_write_n[7] ),
    .Z(net245));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold4 (.I(\u0.mem_write_n[8] ),
    .Z(net246));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold5 (.I(\u0.mem_write_n[4] ),
    .Z(net247));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold6 (.I(\u0.mem_write_n[5] ),
    .Z(net248));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold7 (.I(\u1.output_active ),
    .Z(net249));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold8 (.I(control_trigger),
    .Z(net250));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold9 (.I(\u0.mem_write_n[1] ),
    .Z(net251));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold10 (.I(\u0.mem_write_n[0] ),
    .Z(net252));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold11 (.I(\u1.inverter_select[3] ),
    .Z(net253));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold12 (.I(\u0.cmd[23] ),
    .Z(net254));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold13 (.I(\u0.mem_write_n[3] ),
    .Z(net255));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold14 (.I(\u0.mem_write_n[2] ),
    .Z(net256));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold15 (.I(\u0.mem_write_n[6] ),
    .Z(net257));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold16 (.I(\u0.cmd[22] ),
    .Z(net258));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold17 (.I(\reset_n_sync[0] ),
    .Z(net259));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold18 (.I(\u1.row_col_select[9] ),
    .Z(net260));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold19 (.I(\u1.inverter_select[5] ),
    .Z(net261));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold20 (.I(\u1.inverter_select[4] ),
    .Z(net262));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold21 (.I(\u1.row_col_select[4] ),
    .Z(net263));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold22 (.I(\u1.row_col_select[6] ),
    .Z(net264));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold23 (.I(\u1.inverter_select[9] ),
    .Z(net265));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold24 (.I(\u1.row_col_select[8] ),
    .Z(net266));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold25 (.I(\u1.inverter_select[0] ),
    .Z(net267));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold26 (.I(\u1.col_sel[0] ),
    .Z(net268));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold27 (.I(\u0.cmd[17] ),
    .Z(net269));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold28 (.I(reset_n),
    .Z(net270));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold29 (.I(\u1.row_sel[4] ),
    .Z(net271));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold30 (.I(\latch_data_sync[0] ),
    .Z(net272));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold31 (.I(\u1.row_col_select[1] ),
    .Z(net273));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold32 (.I(\u1.row_col_select[3] ),
    .Z(net274));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold33 (.I(\u1.inverter_select[2] ),
    .Z(net275));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold34 (.I(\u1.row_sel[5] ),
    .Z(net276));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold35 (.I(\u1.inverter_select[1] ),
    .Z(net277));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold36 (.I(\u1.inverter_select[8] ),
    .Z(net278));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold37 (.I(\u1.u1.impulse_gen[0] ),
    .Z(net279));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold38 (.I(\u1.row_col_select[5] ),
    .Z(net280));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold39 (.I(\u1.inverter_select[6] ),
    .Z(net281));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold40 (.I(\u1.inverter_select[7] ),
    .Z(net282));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold41 (.I(\u1.row_col_select[2] ),
    .Z(net283));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold42 (.I(\u1.row_col_select[7] ),
    .Z(net284));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold43 (.I(\u0.cmd[24] ),
    .Z(net285));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold44 (.I(\u0.cmd[25] ),
    .Z(net286));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold45 (.I(\u1.row_col_select[0] ),
    .Z(net287));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold46 (.I(\u0.cmd[3] ),
    .Z(net288));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold47 (.I(\u0.cmd[5] ),
    .Z(net289));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold48 (.I(\u0.cmd[4] ),
    .Z(net290));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold49 (.I(\control_trigger_sync[0] ),
    .Z(net291));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold50 (.I(\u1.row_sel[0] ),
    .Z(net292));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold51 (.I(\u1.row_sel[1] ),
    .Z(net293));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold52 (.I(\u1.col_sel[4] ),
    .Z(net294));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold53 (.I(\u1.col_sel[1] ),
    .Z(net295));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3212__D (.I(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3211__D (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3068__D (.I(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3020__D (.I(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3022__D (.I(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3036__D (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3085__D (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3097__D (.I(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3100__D (.I(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3182__D (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3183__D (.I(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3184__D (.I(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3185__D (.I(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3186__D (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3187__D (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3188__D (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3189__D (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3190__D (.I(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3210__D (.I(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1807__A3 (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2743__A1 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2742__A1 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2741__A1 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1805__A1 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2744__A3 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2739__A1 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2738__A1 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1805__A2 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1806__A2 (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1839__A3 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1835__A1 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1824__A2 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1840__A3 (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1836__A1 (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1828__A2 (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1841__A1 (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1840__A1 (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1839__A1 (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1834__A1 (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1838__A4 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1837__A3 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1836__A2 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1835__A2 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1844__A1 (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2597__A1 (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1869__A2 (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1867__A1 (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1876__A1 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1875__A1 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1873__A1 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1857__A1 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2594__A1 (.I(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1860__C2 (.I(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2611__C (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2408__A1 (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2392__A1 (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1867__B (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1888__A1 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1885__A1 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1874__A1 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1872__A1 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1876__A2 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1875__A3 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1873__A2 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1872__A2 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1886__A2 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1884__A2 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1883__A2 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2163__A1 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2101__A1 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2051__A1 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1890__I (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2202__I0 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2179__I0 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2141__I0 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1899__I1 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2556__A1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2159__A2 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2139__A2 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1896__A2 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1905__I (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1897__I (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1940__I (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1921__I (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1908__I (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1898__I (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1918__S (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1915__S (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1903__S (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1899__S (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2165__A1 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2103__A1 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2053__A1 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1902__I (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2204__I0 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2181__I0 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2143__I0 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1903__I1 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1933__I (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1931__S (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1928__S (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1906__I (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1926__A2 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1923__A2 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1913__A2 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1910__A2 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2794__I1 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2516__A1 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2011__I1 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1909__A1 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1951__A2 (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1948__A2 (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1912__A2 (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1909__A2 (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2796__I1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__A1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2208__I0 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1912__A1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2522__A1 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2211__I0 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2018__I1 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1915__I1 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2524__A1 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2213__I0 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2020__I1 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1918__I1 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2526__A1 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2022__A1 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1981__A1 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1922__A1 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2806__A1 (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2024__A1 (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1983__A1 (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1925__A1 (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2808__I1 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2532__A1 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2026__I1 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1928__I1 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2810__I1 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2534__A1 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2029__I1 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1931__I1 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1945__A2 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1942__A2 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1939__A2 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1936__A2 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2536__A1 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2031__A1 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1990__I1 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1935__A1 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2538__A1 (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2033__A1 (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1993__A1 (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1938__A1 (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2544__A1 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2089__I0 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2038__I1 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1944__A1 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2546__A1 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2040__I1 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1999__A1 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1947__A1 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2548__A1 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2042__I1 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2001__A1 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1950__A1 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2789__A1 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2512__A1 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2005__I1 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1959__I1 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2784__A1 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2554__A1 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2159__A1 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1956__A1 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1967__I (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1957__I (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1987__I (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1977__I (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1964__I (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1958__I (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2792__I1 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2514__A1 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2007__I1 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1962__I1 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1992__I (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1990__S (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1980__I (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1965__I (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1979__A2 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1975__A2 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1972__A2 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1969__A2 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2167__A1 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2106__A1 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2055__I (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1968__A1 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2002__A2 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1974__A2 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1971__A2 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1968__A2 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2108__A1 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2059__I (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2016__A1 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1971__A1 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2799__A1 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2151__A1 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2062__I (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1974__A1 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1975__B (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2801__A1 (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2154__A1 (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2065__I (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1978__A1 (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1997__A2 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1995__A2 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1993__A2 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1988__A2 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2000__A2 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1998__A2 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1996__A2 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1994__A2 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2000__B (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2002__B (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2015__I (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2009__I (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2004__I (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2033__A2 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2031__A2 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2007__S (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2005__S (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2042__S (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2028__I (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2014__I (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2010__I (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2026__S (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2020__S (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2018__S (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2011__S (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2032__A2 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2025__A2 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2023__A2 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2017__A2 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2034__A2 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2024__A2 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2022__A2 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2016__A2 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2040__S (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2038__S (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2036__S (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2029__S (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2542__A1 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2131__I0 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2087__I0 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2036__I1 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2082__I (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2070__I (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2056__I (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2048__I (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2089__S (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2087__S (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2050__I (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2049__I (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2086__A2 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2084__A2 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2054__A2 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2052__A2 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2094__A2 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2092__A2 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2053__A2 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2051__A2 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2206__I0 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2183__I0 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2145__I0 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2057__I0 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2066__S (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2063__S (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2060__S (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2057__S (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2185__I0 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2169__I0 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2147__I0 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2060__I0 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2188__I0 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2171__I0 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2111__I0 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2063__I0 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2190__I0 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2173__I0 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2113__I0 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2066__I0 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2803__A1 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2175__A1 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2157__A1 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2069__I (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2215__I0 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2192__I0 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2115__I0 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2071__I0 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2080__S (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2077__S (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2074__S (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2071__S (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2528__A1 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2217__I0 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2194__I0 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2074__I0 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2219__I0 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2196__I0 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2120__I0 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2077__I0 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2221__I0 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2198__I0 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2122__I0 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2080__I0 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2099__I (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2097__I (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2131__S (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2122__S (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2117__I (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2098__I (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2109__A2 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2107__A2 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2104__A2 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2102__A2 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2128__I (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2110__I (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2105__I (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2100__I (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2138__A2 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2136__A2 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2103__A2 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2101__A2 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2125__A2 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2118__A2 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2108__A2 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2106__A2 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2120__S (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2115__S (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2113__S (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2111__S (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2134__A2 (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2130__A2 (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2126__A2 (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2119__A2 (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2119__B (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2126__B (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2137__A2 (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2135__A2 (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2133__A2 (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2129__A2 (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2130__B (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2150__I (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2147__S (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2145__S (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2140__I (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2157__A2 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2154__A2 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2143__S (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2141__S (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2162__I (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2160__I (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2173__S (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2171__S (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2169__S (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2161__I (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2176__A2 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2168__A2 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2166__A2 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2164__A2 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2175__A2 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2167__A2 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2165__A2 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2163__A2 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2198__S (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2196__S (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2187__I (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2178__I (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2185__S (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2183__S (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2181__S (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2179__S (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2221__S (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2219__S (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2210__I (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2201__I (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2208__S (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2206__S (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2204__S (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2202__S (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2217__S (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2215__S (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2213__S (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2211__S (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2498__A1 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2491__B2 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2262__A1 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2257__A1 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2235__C (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2240__A3 (.I(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2246__A2 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2246__A3 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2246__B1 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2248__A2 (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2253__A4 (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2266__I (.I(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2259__A2 (.I(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2254__I (.I(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2436__I (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2357__I (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2324__I (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2255__I (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2484__A1 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2283__A2 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2278__A2 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2256__A2 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2288__I (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2262__A2 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2260__I (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2434__I (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2390__I (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2383__I (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2261__I (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2498__A2 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2285__A2 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2280__A2 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2270__A2 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2442__I (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2297__I (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2263__I (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2503__A1 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2485__B (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2480__B (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2264__I (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2295__B1 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2285__B1 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2280__B1 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2270__B1 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2430__S (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2379__S (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2367__S (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2269__S (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2395__I (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2338__I (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2307__I (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2273__I (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2304__A1 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2294__A1 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2284__A1 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2279__A1 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2318__A2 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2311__A2 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2305__A2 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2295__A2 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2314__A4 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2300__A2 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2299__A3 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2291__A2 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2316__A2 (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2309__A2 (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2303__A2 (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2293__A2 (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2327__B1 (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2318__B1 (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2311__B1 (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2305__B1 (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2335__A1 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2326__A1 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2317__A1 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2310__A1 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2457__A4 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2332__A4 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2322__A2 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2315__A2 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2457__A3 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2332__A3 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2330__A1 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2327__A1 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2350__A2 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2342__A2 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2336__A2 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2327__A2 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2348__A2 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2340__A2 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2334__A2 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2325__A2 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2360__B1 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2350__B1 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2342__B1 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2336__B1 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2364__A3 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2346__A2 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2339__A2 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2333__A2 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2337__I (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2373__A1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2359__A1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2349__A1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2341__A1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2355__A2 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2353__A1 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2350__A1 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2345__I (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2351__I (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2380__A2 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2374__A2 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2368__A2 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2360__A2 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2366__A2 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2356__A2 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2420__A2 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2415__A2 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2372__A2 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2358__A2 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2402__B1 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2380__B1 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2374__B1 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2368__B1 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2386__A3 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2377__A2 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2371__A2 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2366__B (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2459__A2 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2386__A2 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2377__A1 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2374__A1 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2375__I (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2459__A1 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2386__A1 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2380__A1 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2378__A1 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2381__I (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2486__A2 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2481__A2 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2409__A2 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2393__A2 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2479__A2 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2472__A1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2407__A1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2391__A1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2489__B (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2406__A2 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2400__C (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2389__A2 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2497__A2 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2473__A2 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2407__C (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2391__C (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2431__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2422__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2417__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2402__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2490__A2 (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2485__A2 (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2447__A2 (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2401__A2 (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2427__A3 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2412__A2 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2405__A2 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2399__I (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2403__I (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2460__A2 (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2413__A2 (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2409__A1 (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2405__A1 (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2439__B1 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2431__B1 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2422__B1 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2417__B1 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2453__A1 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2438__A1 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2421__A1 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2416__A1 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2424__A2 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2419__A2 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2414__A2 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2429__A2 (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2460__A4 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2426__I (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2468__A4 (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2428__I (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2465__A2 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2454__A2 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2448__A2 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2439__A2 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2471__A2 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2452__A2 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2446__A1 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2437__A2 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2473__B1 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2465__B1 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2454__B1 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2448__B1 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2451__A2 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2446__A3 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2449__I (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2475__A2 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2468__A1 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2465__A1 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2462__A1 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2458__A3 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2461__A4 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2475__A3 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2462__A2 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2502__S (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2495__C (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2477__I (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2464__S (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2488__A4 (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2478__A2 (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2494__A2 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2487__A2 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2483__A2 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2478__B (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2492__A2 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2478__C (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2501__A1 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2488__A2 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2486__A1 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2483__A1 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2495__A2 (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2489__A2 (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2496__A2 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2501__A2 (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2550__I (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2507__I (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2540__I (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2530__I (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2520__I (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2508__I (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2541__I (.I(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2531__I (.I(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2521__I (.I(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2511__I (.I(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2513__I (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2515__I (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__I (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2549__I (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2582__I (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2572__I (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2562__I (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2551__I (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2583__I (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2573__I (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2563__I (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2553__I (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2580__A2 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2578__A2 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2576__A2 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2574__A2 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2580__B1 (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2578__B1 (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2576__B1 (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2574__B1 (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2593__A3 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2597__A2 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2615__A2 (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2614__A2 (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2612__A1 (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2617__A1 (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2604__B2 (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2602__A2 (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2627__A1 (.I(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2624__A1 (.I(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2621__A1 (.I(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2613__I (.I(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2632__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2630__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2618__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2616__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2623__A2 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2622__A2 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2621__A2 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2621__A3 (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2637__A1 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2650__A2 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2650__B (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2648__B (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2650__C (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2658__A2 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2658__B (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2664__A3 (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2737__I (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2683__I (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2671__I (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2666__I (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2764__C (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2762__C (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2759__C (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2667__I (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2711__A1 (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2682__A1 (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2670__A1 (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2668__A2 (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2732__A1 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2680__A1 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2677__A1 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2674__A1 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2689__A3 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2679__A2 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2678__A2 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2677__A3 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2687__A2 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2686__A1 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2681__A2 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2680__A2 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2735__I (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2715__I (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2700__I (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2684__I (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2699__A1 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2695__A1 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2692__A1 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2688__A1 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2689__A4 (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2686__A2 (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2714__A1 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2709__A1 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2706__A1 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2703__A1 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2712__A4 (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2708__A2 (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2707__A2 (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2706__A2 (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2713__A2 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2710__A2 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2709__A2 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2717__A2 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2716__A2 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2714__A2 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2730__A1 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2727__A1 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2724__A1 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2719__A1 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2726__A4 (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2723__A3 (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2718__I (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2722__A2 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2721__B1 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2720__A2 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2719__A3 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2744__A4 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2739__A2 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2738__A2 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2736__B (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2756__A1 (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2750__C (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2742__C (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2736__C (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2753__A1 (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2748__A1 (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2745__A1 (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2740__A1 (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2752__A4 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2747__A2 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2746__A2 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2745__A3 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2761__A4 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2755__A2 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2754__A2 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2753__A3 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2770__A1 (.I(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2772__A1 (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2774__A1 (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2776__A1 (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2778__A1 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2780__A1 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2782__A1 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2812__I (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2791__I (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2785__I (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2805__I (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2798__I (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2788__I (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2786__I (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2810__S (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2808__S (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2796__S (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2787__I (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2804__A2 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2802__A2 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2800__A2 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2790__A2 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2824__A2 (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2822__A2 (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2794__S (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2792__S (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2806__A2 (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2803__A2 (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2801__A2 (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2799__A2 (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2827__I (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2829__I (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2831__I (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2590__A1 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1820__A1 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1533__A1 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1418__A1 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2505__I (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1417__I (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2633__A4 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2509__A1 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1533__A3 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1418__A3 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1544__A1 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1530__A1 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1525__A1 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1522__A1 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1527__A2 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1420__A2 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2419__A1 (.I(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1431__A1 (.I(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1426__B1 (.I(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2246__B2 (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1431__B (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2246__A1 (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1445__A1 (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2242__A2 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2109__A1 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1438__A2 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2397__A2 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2387__A1 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2382__I (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1438__B1 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2102__A1 (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1438__B2 (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1437__B2 (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2401__A1 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2104__A1 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1444__B2 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1437__A2 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2460__A1 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2413__A1 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1441__A1 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2402__A1 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2400__A1 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2397__A1 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1444__B1 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2138__A1 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1458__A2 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1449__A2 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2251__B (.I(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1450__C (.I(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2491__A1 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2488__A1 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1452__A1 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2136__A1 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1458__B2 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1455__A2 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2497__A1 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2495__A1 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2493__A1 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1458__B1 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2251__A1 (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1459__A3 (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2248__A1 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1470__A1 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2476__A3 (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2461__A1 (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2450__I (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1465__A1 (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2470__A1 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1469__B1 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1464__A1 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2247__C1 (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1465__B (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1470__A2 (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2247__C2 (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1470__A3 (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2488__A3 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2481__A1 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2478__A1 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1469__A1 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2252__A1 (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2224__A2 (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1519__A2 (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2398__A1 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2376__I (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2229__I (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1474__A1 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2094__A1 (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1480__A2 (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1474__A2 (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2092__A1 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1474__B2 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2371__A1 (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1477__A1 (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2354__A1 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1482__A1 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1481__B1 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2086__A1 (.I(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1489__A2 (.I(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1480__B2 (.I(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2234__B (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1495__A1 (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2334__A1 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2232__A2 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2080__I1 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1490__A2 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2325__A1 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2077__I1 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1493__A2 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1490__B2 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2084__A1 (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1489__B2 (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2234__A1 (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1490__C (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2458__A2 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2364__A2 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2346__A1 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1492__A1 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2235__A1 (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1519__A3 (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2301__A1 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1506__B1 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1498__A1 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2291__A1 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1505__B1 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1498__B1 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2315__A1 (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1504__A1 (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1501__A1 (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1512__A1 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1505__A1 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2228__B2 (.I(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1505__C (.I(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2052__A1 (.I(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1510__A2 (.I(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2054__A1 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1515__A2 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1510__B2 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2225__A1 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1518__A2 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2276__A1 (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1516__A1 (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1512__B1 (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2225__A2 (.I(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1517__B (.I(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1816__A2 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1786__A2 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1543__A2 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1520__I (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1542__B1 (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1528__A2 (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1841__A3 (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1817__A3 (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1534__B (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1539__I (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2580__A1 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1838__A2 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1832__A2 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1542__B2 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2663__A1 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1552__C (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1782__A1 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1738__A1 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1567__A2 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1554__A2 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2663__A2 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1557__A1 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2662__A2 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1733__A1 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1566__A2 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1556__B2 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2663__B1 (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1569__A2 (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2662__C1 (.I(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1564__B (.I(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2661__A2 (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1564__C (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2663__C (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1568__A3 (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2659__A1 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2237__A1 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1661__A1 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2644__A2 (.I(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1663__I (.I(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1583__B2 (.I(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1571__I (.I(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2643__A2 (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1668__A1 (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1577__A2 (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1668__B2 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1577__B2 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2644__B1 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1979__A1 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1580__A1 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1984__A1 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1583__A1 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2644__A1 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1982__A1 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1583__B1 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2647__C (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2240__A1 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1604__A1 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2673__B (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1790__A4 (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1598__B2 (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1586__I (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2672__A3 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1753__A1 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1751__B2 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1587__A2 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2646__A1 (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2239__A1 (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1593__A2 (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2597__B (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2253__A1 (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1785__I (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1603__A1 (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2675__A1 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1790__A3 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1750__I (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1598__A2 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2646__A2 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1602__A1 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1661__A2 (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2731__A1 (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1721__A1 (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1718__B2 (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1617__A2 (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2656__B (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2651__A1 (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1614__A1 (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2736__A1 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1720__A1 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1718__A1 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1616__A2 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2657__B1 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2237__A2 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1628__A1 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1719__A1 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1717__A1 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1624__A2 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1620__A2 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1722__A1 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1717__B2 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1625__A2 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1620__B2 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2698__A1 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1791__A3 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1657__A2 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1633__A2 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2694__A1 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2693__A1 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1791__A4 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1633__B2 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2000__A1 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1637__B1 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2713__B (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2712__A1 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1689__B2 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1637__B2 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1788__A1 (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1768__A1 (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1690__A1 (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1641__A2 (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1788__A2 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1690__B2 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1641__B2 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2642__B1 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1648__A1 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2650__A1 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1659__A2 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2696__A2 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1697__A1 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1692__B2 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1658__A2 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2638__B2 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1677__B2 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1656__A2 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1655__B2 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2638__A2 (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1680__A1 (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1677__A1 (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1652__A2 (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2705__A1 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2704__A1 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1791__A1 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1655__A2 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2649__A1 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2240__A2 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1660__A2 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2721__A1 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2665__A1 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1662__I (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2802__A1 (.I(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1671__A2 (.I(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1667__B1 (.I(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2687__A1 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1789__A3 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1671__A1 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1667__B2 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2807__A1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1763__A2 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1674__A2 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1784__A1 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1761__A1 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2696__A1 (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1692__A1 (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1682__A1 (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1765__B1 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1758__A1 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1700__A1 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2717__A1 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2716__A1 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2641__A2 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1689__A1 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2819__A1 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1696__A2 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1695__B1 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2708__A1 (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2707__A1 (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1787__I (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1695__B2 (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1757__A1 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2652__A2 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1799__I (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1708__A1 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1706__A1 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1913__A1 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1708__A2 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1706__A2 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1910__A1 (.I(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1707__A2 (.I(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1706__B1 (.I(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2726__A1 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2652__B (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1707__A1 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1705__I (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2729__A2 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2725__A1 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1802__A2 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1706__B2 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1926__A1 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1714__A2 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1713__A2 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1923__A1 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1713__B1 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1776__B1 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1757__A2 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1939__A1 (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1778__A2 (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1729__A2 (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1936__A1 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1778__B1 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1729__B1 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2764__A1 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2763__A1 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1797__A1 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1737__A1 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1782__B1 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1739__A3 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1781__A1 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1744__A2 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1783__A1 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1756__A1 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1761__A2 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1754__B (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1764__A1 (.I(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1764__B (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1776__B2 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1783__B (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1784__B (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2664__A1 (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2223__I (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1866__I (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1786__A1 (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2259__A1 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1808__A2 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1807__A1 (.I(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1792__A1 (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1792__A3 (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1807__A2 (.I(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1798__A2 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_clock_I (.I(clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold8_I (.I(control_trigger));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1523__A2 (.I(control_trigger));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1419__A2 (.I(control_trigger));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_control_trigger_in));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_latch_data_in));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_reset_n_in));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(la_data_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(la_data_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(la_data_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(la_data_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(la_data_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(la_data_in[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(la_data_in[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(la_data_in[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(la_data_in[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(la_data_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(la_data_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(la_data_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(la_data_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(la_data_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(la_data_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(la_data_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(la_data_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(la_data_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(la_oenb[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(la_oenb[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(la_oenb[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(la_oenb[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(la_oenb[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(la_oenb[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(la_oenb[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(la_oenb[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(la_oenb[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(la_oenb[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(la_oenb[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(la_oenb[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(la_oenb[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(la_oenb[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(la_oenb[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(la_oenb[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_I (.I(la_oenb[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_I (.I(la_oenb[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold1_I (.I(latch_data));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2633__A2 (.I(latch_data));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_I (.I(spi_data[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_I (.I(spi_data[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input42_I (.I(spi_data[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input43_I (.I(spi_data[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input44_I (.I(spi_data[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input45_I (.I(spi_data[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input46_I (.I(spi_data[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input47_I (.I(spi_data[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input48_I (.I(spi_data[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input49_I (.I(spi_data[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input50_I (.I(spi_data[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input51_I (.I(spi_data[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input52_I (.I(spi_data[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input53_I (.I(spi_data[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input54_I (.I(spi_data[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input55_I (.I(spi_data[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input56_I (.I(spi_data[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input57_I (.I(spi_data[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input58_I (.I(spi_data[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input59_I (.I(spi_data[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input60_I (.I(spi_data[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input61_I (.I(spi_data[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input62_I (.I(spi_data[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input63_I (.I(spi_data[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input64_I (.I(spi_data[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input65_I (.I(spi_data[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input66_I (.I(spi_data[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input67_I (.I(spi_data[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input68_I (.I(spi_data[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input69_I (.I(spi_data[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input70_I (.I(spi_data[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input71_I (.I(spi_data[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input72_I (.I(spi_data_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3119__D (.I(\spi_data_crossing[0].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2512__B2 (.I(\spi_data_crossing[0].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2536__B2 (.I(\spi_data_crossing[10].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2538__B2 (.I(\spi_data_crossing[11].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3143__D (.I(\spi_data_crossing[12].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3145__D (.I(\spi_data_crossing[13].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2546__B2 (.I(\spi_data_crossing[14].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2548__B2 (.I(\spi_data_crossing[15].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2560__B2 (.I(\spi_data_crossing[19].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3121__D (.I(\spi_data_crossing[1].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2514__B2 (.I(\spi_data_crossing[1].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2574__B2 (.I(\spi_data_crossing[24].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3169__D (.I(\spi_data_crossing[25].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3171__D (.I(\spi_data_crossing[26].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3173__D (.I(\spi_data_crossing[27].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3177__D (.I(\spi_data_crossing[29].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2586__B2 (.I(\spi_data_crossing[29].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2516__B2 (.I(\spi_data_crossing[2].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3179__D (.I(\spi_data_crossing[30].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__B2 (.I(\spi_data_crossing[3].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2522__B2 (.I(\spi_data_crossing[4].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3129__D (.I(\spi_data_crossing[5].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2524__B2 (.I(\spi_data_crossing[5].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3131__D (.I(\spi_data_crossing[6].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2526__B2 (.I(\spi_data_crossing[6].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3133__D (.I(\spi_data_crossing[7].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2528__B2 (.I(\spi_data_crossing[7].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2532__B2 (.I(\spi_data_crossing[8].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2534__B2 (.I(\spi_data_crossing[9].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2844__D (.I(\u0.cmd[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1952__I (.I(\u0.cmd[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1889__I (.I(\u0.cmd[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout224_I (.I(\u0.cmd[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2125__A1 (.I(\u0.cmd[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout223_I (.I(\u0.cmd[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2129__A1 (.I(\u0.cmd[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout222_I (.I(\u0.cmd[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2818__A1 (.I(\u0.cmd[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout221_I (.I(\u0.cmd[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2133__A1 (.I(\u0.cmd[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout220_I (.I(\u0.cmd[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2135__A1 (.I(\u0.cmd[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout219_I (.I(\u0.cmd[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2137__A1 (.I(\u0.cmd[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3234__D (.I(\u0.cmd[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2044__A1 (.I(\u0.cmd[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1953__I (.I(\u0.cmd[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1891__I (.I(\u0.cmd[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold27_I (.I(\u0.cmd[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1954__I (.I(\u0.cmd[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1892__I (.I(\u0.cmd[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3236__D (.I(\u0.cmd[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2558__A1 (.I(\u0.cmd[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2045__A1 (.I(\u0.cmd[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1894__A2 (.I(\u0.cmd[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout218_I (.I(\u0.cmd[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2200__A1 (.I(\u0.cmd[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2845__D (.I(\u0.cmd[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1961__I (.I(\u0.cmd[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1901__I (.I(\u0.cmd[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3238__D (.I(\u0.cmd[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2564__A1 (.I(\u0.cmd[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2046__A3 (.I(\u0.cmd[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1894__A4 (.I(\u0.cmd[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3239__D (.I(\u0.cmd[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2566__A1 (.I(\u0.cmd[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2046__A2 (.I(\u0.cmd[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1894__A3 (.I(\u0.cmd[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold16_I (.I(\u0.cmd[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2568__A1 (.I(\u0.cmd[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1830__A1 (.I(\u0.cmd[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1825__I (.I(\u0.cmd[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1823__A2 (.I(\u0.cmd[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1420__A1 (.I(\u0.cmd[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2584__A1 (.I(\u0.cmd[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1833__I (.I(\u0.cmd[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1821__A1 (.I(\u0.cmd[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1524__A1 (.I(\u0.cmd[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2586__A1 (.I(\u0.cmd[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1834__A2 (.I(\u0.cmd[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1821__A2 (.I(\u0.cmd[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1531__I (.I(\u0.cmd[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2846__D (.I(\u0.cmd[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1966__I (.I(\u0.cmd[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1907__I (.I(\u0.cmd[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2588__A1 (.I(\u0.cmd[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1819__I (.I(\u0.cmd[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1533__A2 (.I(\u0.cmd[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1418__A2 (.I(\u0.cmd[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold46_I (.I(\u0.cmd[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1970__I (.I(\u0.cmd[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1911__I (.I(\u0.cmd[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold48_I (.I(\u0.cmd[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1973__I (.I(\u0.cmd[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1914__I (.I(\u0.cmd[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold47_I (.I(\u0.cmd[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1976__I (.I(\u0.cmd[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1917__I (.I(\u0.cmd[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2850__D (.I(\u0.cmd[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2068__I (.I(\u0.cmd[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1920__I (.I(\u0.cmd[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2851__D (.I(\u0.cmd[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2118__A1 (.I(\u0.cmd[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2073__I (.I(\u0.cmd[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1924__I (.I(\u0.cmd[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2852__D (.I(\u0.cmd[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2076__I (.I(\u0.cmd[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1985__A1 (.I(\u0.cmd[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1927__I (.I(\u0.cmd[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2853__D (.I(\u0.cmd[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2079__I (.I(\u0.cmd[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1988__A1 (.I(\u0.cmd[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1930__I (.I(\u0.cmd[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1869__A1 (.I(\u0.timer_enable ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1594__I (.I(\u0.timer_enable ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2783__I (.I(\u1.ccr0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1754__A2 (.I(\u1.ccr0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1748__B1 (.I(\u1.ccr0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1915__I0 (.I(\u1.ccr0[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1721__A2 (.I(\u1.ccr0[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1718__B1 (.I(\u1.ccr0[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1715__A2 (.I(\u1.ccr0[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1712__I (.I(\u1.ccr0[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1931__I0 (.I(\u1.ccr0[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1731__B1 (.I(\u1.ccr0[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1730__A2 (.I(\u1.ccr0[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1731__A2 (.I(\u1.ccr0[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1727__I (.I(\u1.ccr0[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1733__B1 (.I(\u1.ccr0[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1726__I (.I(\u1.ccr0[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1741__I (.I(\u1.ccr0[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1733__A2 (.I(\u1.ccr0[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1782__A2 (.I(\u1.ccr0[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1738__A2 (.I(\u1.ccr0[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1735__I (.I(\u1.ccr0[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2796__I0 (.I(\u1.ccr0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1752__A2 (.I(\u1.ccr0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1751__A2 (.I(\u1.ccr0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2808__I0 (.I(\u1.ccr0[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1697__A2 (.I(\u1.ccr0[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1692__B1 (.I(\u1.ccr0[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2810__I0 (.I(\u1.ccr0[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1692__A2 (.I(\u1.ccr0[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1682__A2 (.I(\u1.ccr0[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1959__I0 (.I(\u1.ccr1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1599__A2 (.I(\u1.ccr1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1592__A2 (.I(\u1.ccr1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2638__B1 (.I(\u1.ccr1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1990__I0 (.I(\u1.ccr1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1656__A1 (.I(\u1.ccr1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1655__B1 (.I(\u1.ccr1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1645__I (.I(\u1.ccr1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1641__C1 (.I(\u1.ccr1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2005__I0 (.I(\u1.ccr1[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1625__A1 (.I(\u1.ccr1[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1620__B1 (.I(\u1.ccr1[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2007__I0 (.I(\u1.ccr1[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1624__A1 (.I(\u1.ccr1[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1620__A1 (.I(\u1.ccr1[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2655__A1 (.I(\u1.ccr1[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2011__I0 (.I(\u1.ccr1[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1622__A1 (.I(\u1.ccr1[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1962__I0 (.I(\u1.ccr1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1600__A1 (.I(\u1.ccr1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1592__B1 (.I(\u1.ccr1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2020__I0 (.I(\u1.ccr1[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1616__A1 (.I(\u1.ccr1[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1613__C1 (.I(\u1.ccr1[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2656__A1 (.I(\u1.ccr1[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1613__A1 (.I(\u1.ccr1[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1607__I (.I(\u1.ccr1[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2660__A1 (.I(\u1.ccr1[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2029__I0 (.I(\u1.ccr1[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1565__A1 (.I(\u1.ccr1[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1552__A1 (.I(\u1.ccr1[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2662__A1 (.I(\u1.ccr1[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2036__I0 (.I(\u1.ccr1[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1566__A1 (.I(\u1.ccr1[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1556__B1 (.I(\u1.ccr1[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1578__I (.I(\u1.ccr1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1574__B1 (.I(\u1.ccr1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1582__I (.I(\u1.ccr1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1574__A1 (.I(\u1.ccr1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2643__A1 (.I(\u1.ccr1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1581__I (.I(\u1.ccr1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1577__A1 (.I(\u1.ccr1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1658__A1 (.I(\u1.ccr1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1631__I (.I(\u1.ccr1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2888__D (.I(\u1.ccr1_flag ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2595__A2 (.I(\u1.col_limit[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2169__I1 (.I(\u1.col_limit[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1860__A2 (.I(\u1.col_limit[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1852__A2 (.I(\u1.col_limit[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2171__I1 (.I(\u1.col_limit[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1861__B2 (.I(\u1.col_limit[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1852__B2 (.I(\u1.col_limit[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2173__I1 (.I(\u1.col_limit[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1861__A2 (.I(\u1.col_limit[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1849__A2 (.I(\u1.col_limit[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2841__D (.I(\u1.col_sel[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1879__A1 (.I(\u1.col_sel[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1878__A1 (.I(\u1.col_sel[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1850__I (.I(\u1.col_sel[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold35_I (.I(\u1.inverter_select[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2181__I1 (.I(\u1.inverter_select[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1517__A2 (.I(\u1.ordering_complete[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1508__I (.I(\u1.ordering_complete[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2340__A1 (.I(\u1.ordering_complete[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1492__A2 (.I(\u1.ordering_complete[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1488__I (.I(\u1.ordering_complete[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2348__A1 (.I(\u1.ordering_complete[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1479__I (.I(\u1.ordering_complete[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2358__A1 (.I(\u1.ordering_complete[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2087__I1 (.I(\u1.ordering_complete[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1482__A2 (.I(\u1.ordering_complete[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1481__B2 (.I(\u1.ordering_complete[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2367__I0 (.I(\u1.ordering_complete[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2089__I1 (.I(\u1.ordering_complete[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1481__A2 (.I(\u1.ordering_complete[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1477__B2 (.I(\u1.ordering_complete[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2372__A1 (.I(\u1.ordering_complete[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1477__A2 (.I(\u1.ordering_complete[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1473__I (.I(\u1.ordering_complete[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2379__I0 (.I(\u1.ordering_complete[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2231__A2 (.I(\u1.ordering_complete[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1472__I (.I(\u1.ordering_complete[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2389__A1 (.I(\u1.ordering_complete[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1435__I (.I(\u1.ordering_complete[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2406__A1 (.I(\u1.ordering_complete[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1442__I (.I(\u1.ordering_complete[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1441__B2 (.I(\u1.ordering_complete[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2415__A1 (.I(\u1.ordering_complete[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1441__A2 (.I(\u1.ordering_complete[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1433__I (.I(\u1.ordering_complete[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2269__I0 (.I(\u1.ordering_complete[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1509__I (.I(\u1.ordering_complete[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2420__A1 (.I(\u1.ordering_complete[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2111__I1 (.I(\u1.ordering_complete[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1431__A2 (.I(\u1.ordering_complete[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1426__B2 (.I(\u1.ordering_complete[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2430__I0 (.I(\u1.ordering_complete[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2113__I1 (.I(\u1.ordering_complete[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1428__B2 (.I(\u1.ordering_complete[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1426__A2 (.I(\u1.ordering_complete[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2437__A1 (.I(\u1.ordering_complete[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2115__I1 (.I(\u1.ordering_complete[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1428__A2 (.I(\u1.ordering_complete[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1423__B2 (.I(\u1.ordering_complete[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2452__A1 (.I(\u1.ordering_complete[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2120__I1 (.I(\u1.ordering_complete[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1461__I (.I(\u1.ordering_complete[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2471__A1 (.I(\u1.ordering_complete[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2124__I (.I(\u1.ordering_complete[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1469__B2 (.I(\u1.ordering_complete[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1464__A2 (.I(\u1.ordering_complete[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2127__I (.I(\u1.ordering_complete[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1469__A2 (.I(\u1.ordering_complete[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1450__B2 (.I(\u1.ordering_complete[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2485__A1 (.I(\u1.ordering_complete[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2131__I1 (.I(\u1.ordering_complete[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1452__B2 (.I(\u1.ordering_complete[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1450__A2 (.I(\u1.ordering_complete[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2490__A1 (.I(\u1.ordering_complete[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1454__I (.I(\u1.ordering_complete[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1452__A2 (.I(\u1.ordering_complete[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2502__I0 (.I(\u1.ordering_complete[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1448__I (.I(\u1.ordering_complete[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2283__A1 (.I(\u1.ordering_complete[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2060__I1 (.I(\u1.ordering_complete[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1512__A2 (.I(\u1.ordering_complete[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1505__A2 (.I(\u1.ordering_complete[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2293__A1 (.I(\u1.ordering_complete[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2063__I1 (.I(\u1.ordering_complete[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1505__B2 (.I(\u1.ordering_complete[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1498__B2 (.I(\u1.ordering_complete[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2303__A1 (.I(\u1.ordering_complete[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2066__I1 (.I(\u1.ordering_complete[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1506__B2 (.I(\u1.ordering_complete[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1498__A2 (.I(\u1.ordering_complete[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2309__A1 (.I(\u1.ordering_complete[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2071__I1 (.I(\u1.ordering_complete[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1506__A2 (.I(\u1.ordering_complete[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1501__B2 (.I(\u1.ordering_complete[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2316__A1 (.I(\u1.ordering_complete[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2074__I1 (.I(\u1.ordering_complete[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1504__A2 (.I(\u1.ordering_complete[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1501__A2 (.I(\u1.ordering_complete[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2232__B2 (.I(\u1.ordering_complete[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1487__I (.I(\u1.ordering_complete[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1492__B2 (.I(\u1.ordering_complete[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1485__I (.I(\u1.ordering_complete[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2342__A1 (.I(\u1.ordering_timer[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2339__A1 (.I(\u1.ordering_timer[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1491__I (.I(\u1.ordering_timer[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1489__B1 (.I(\u1.ordering_timer[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2344__I (.I(\u1.ordering_timer[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1489__A1 (.I(\u1.ordering_timer[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1480__B1 (.I(\u1.ordering_timer[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2368__A1 (.I(\u1.ordering_timer[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2363__A1 (.I(\u1.ordering_timer[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1476__I (.I(\u1.ordering_timer[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2398__A2 (.I(\u1.ordering_timer[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2370__I (.I(\u1.ordering_timer[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1475__I (.I(\u1.ordering_timer[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1474__B1 (.I(\u1.ordering_timer[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2427__A2 (.I(\u1.ordering_timer[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2412__A1 (.I(\u1.ordering_timer[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1444__A1 (.I(\u1.ordering_timer[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1440__I (.I(\u1.ordering_timer[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2241__I (.I(\u1.ordering_timer[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1439__I (.I(\u1.ordering_timer[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1438__A1 (.I(\u1.ordering_timer[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2431__A1 (.I(\u1.ordering_timer[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2425__A1 (.I(\u1.ordering_timer[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1424__I (.I(\u1.ordering_timer[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2468__A3 (.I(\u1.ordering_timer[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2433__I (.I(\u1.ordering_timer[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1422__I (.I(\u1.ordering_timer[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2441__I (.I(\u1.ordering_timer[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1430__A1 (.I(\u1.ordering_timer[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1421__I (.I(\u1.ordering_timer[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2467__I (.I(\u1.ordering_timer[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2247__B1 (.I(\u1.ordering_timer[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1462__I (.I(\u1.ordering_timer[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2500__A1 (.I(\u1.ordering_timer[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2476__A1 (.I(\u1.ordering_timer[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2247__A1 (.I(\u1.ordering_timer[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1447__I (.I(\u1.ordering_timer[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2494__A1 (.I(\u1.ordering_timer[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2487__A1 (.I(\u1.ordering_timer[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1446__I (.I(\u1.ordering_timer[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2290__A4 (.I(\u1.ordering_timer[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2280__A1 (.I(\u1.ordering_timer[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2274__A3 (.I(\u1.ordering_timer[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1511__I (.I(\u1.ordering_timer[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1457__I (.I(\u1.ordering_timer[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1455__A1 (.I(\u1.ordering_timer[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2314__A1 (.I(\u1.ordering_timer[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2311__A1 (.I(\u1.ordering_timer[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2308__A1 (.I(\u1.ordering_timer[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1500__I (.I(\u1.ordering_timer[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2457__A2 (.I(\u1.ordering_timer[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2336__A1 (.I(\u1.ordering_timer[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2332__A2 (.I(\u1.ordering_timer[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1484__I (.I(\u1.ordering_timer[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold45_I (.I(\u1.row_col_select[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2202__I1 (.I(\u1.row_col_select[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold42_I (.I(\u1.row_col_select[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2217__I1 (.I(\u1.row_col_select[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold24_I (.I(\u1.row_col_select[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2219__I1 (.I(\u1.row_col_select[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2605__B1 (.I(\u1.row_limit[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2604__A1 (.I(\u1.row_limit[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2145__I1 (.I(\u1.row_limit[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold50_I (.I(\u1.row_sel[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2615__A1 (.I(\u1.row_sel[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2614__A1 (.I(\u1.row_sel[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2601__I (.I(\u1.row_sel[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold51_I (.I(\u1.row_sel[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2620__A1 (.I(\u1.row_sel[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2619__A2 (.I(\u1.row_sel[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2600__I (.I(\u1.row_sel[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2834__D (.I(\u1.row_sel[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2620__B (.I(\u1.row_sel[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2619__A1 (.I(\u1.row_sel[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2603__I (.I(\u1.row_sel[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1683__I (.I(\u1.timer[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1646__A2 (.I(\u1.timer[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1640__I (.I(\u1.timer[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1686__I (.I(\u1.timer[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1638__I (.I(\u1.timer[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1637__A2 (.I(\u1.timer[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2726__A3 (.I(\u1.timer[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2723__A2 (.I(\u1.timer[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1801__I (.I(\u1.timer[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1619__I (.I(\u1.timer[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2676__A2 (.I(\u1.timer[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1590__I (.I(\u1.timer[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2734__A1 (.I(\u1.timer[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1805__A3 (.I(\u1.timer[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1612__I (.I(\u1.timer[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2744__A1 (.I(\u1.timer[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2743__B (.I(\u1.timer[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1795__A4 (.I(\u1.timer[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1547__I (.I(\u1.timer[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2761__A1 (.I(\u1.timer[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1797__A2 (.I(\u1.timer[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1737__B2 (.I(\u1.timer[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1549__I (.I(\u1.timer[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2689__A2 (.I(\u1.timer[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1670__I (.I(\u1.timer[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1580__B2 (.I(\u1.timer[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1576__I (.I(\u1.timer[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2689__A1 (.I(\u1.timer[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1672__I (.I(\u1.timer[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1583__A2 (.I(\u1.timer[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1575__I (.I(\u1.timer[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1813__I1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1811__I1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1809__I1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2826__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2767__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2765__I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2828__A1 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2830__A1 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1809__I0 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1811__I0 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1813__I0 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1815__A1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1811__S (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3172__D (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3174__D (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3122__D (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3180__D (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output85_I (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3266__I (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output86_I (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3267__I (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output88_I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3269__I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output95_I (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3270__I (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output96_I (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3280__I (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output97_I (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3281__I (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output98_I (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3282__I (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output99_I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3283__I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output100_I (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3284__I (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output101_I (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3285__I (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output102_I (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3271__I (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output103_I (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3272__I (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output104_I (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3273__I (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output105_I (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3274__I (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output106_I (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3275__I (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output107_I (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3276__I (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output108_I (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3277__I (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output109_I (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3278__I (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output110_I (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3279__I (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output119_I (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output126_I (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output129_I (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output130_I (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output131_I (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output146_I (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3294__I (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output159_I (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output160_I (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output161_I (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output162_I (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3296__I (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output163_I (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3297__I (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output164_I (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3298__I (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output165_I (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3299__I (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output166_I (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3300__I (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output167_I (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3301__I (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output168_I (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3302__I (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output169_I (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3303__I (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output170_I (.I(net170));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3304__I (.I(net170));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output181_I (.I(net181));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output187_I (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output192_I (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3306__I (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output196_I (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output197_I (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output201_I (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output203_I (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output204_I (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3307__I (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output205_I (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3308__I (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output206_I (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3309__I (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output207_I (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3310__I (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output209_I (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3312__I (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2608__A2 (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2609__B2 (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2631__A1 (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2628__I (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2625__A1 (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2626__A1 (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2598__I (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2608__B2 (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2177__A1 (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1893__I (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3237__D (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2560__A1 (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2859__D (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2824__A1 (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2093__A1 (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1949__I (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2858__D (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2822__A1 (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1946__I (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2091__A1 (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1997__A1 (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2857__D (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2820__A1 (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1943__I (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1995__A1 (.I(net222));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2856__D (.I(net222));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2035__I (.I(net222));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1941__A1 (.I(net222));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2855__D (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2816__A1 (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2085__A1 (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1937__I (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2854__D (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2813__A1 (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2083__A1 (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1934__I (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3122__CLK (.I(net229));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3120__CLK (.I(net229));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout227_I (.I(net229));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout228_I (.I(net229));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout232_I (.I(net233));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout229_I (.I(net233));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3176__CLK (.I(net238));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout237_I (.I(net238));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout238_I (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3164__CLK (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3162__CLK (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3160__CLK (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3180__CLK (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3174__CLK (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3172__CLK (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout239_I (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout240_I (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout236_I (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout241_I (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout233_I (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3129__CLK (.I(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3143__CLK (.I(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3141__CLK (.I(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3131__CLK (.I(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2934__CLK (.I(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2935__CLK (.I(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3139__CLK (.I(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2936__CLK (.I(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2937__CLK (.I(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3137__CLK (.I(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3135__CLK (.I(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2905__CLK (.I(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2931__CLK (.I(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2898__CLK (.I(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3047__CLK (.I(clknet_leaf_1_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3051__CLK (.I(clknet_leaf_1_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3050__CLK (.I(clknet_leaf_1_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3044__CLK (.I(clknet_leaf_1_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3045__CLK (.I(clknet_leaf_1_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3046__CLK (.I(clknet_leaf_1_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3145__CLK (.I(clknet_leaf_1_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3149__CLK (.I(clknet_leaf_1_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3147__CLK (.I(clknet_leaf_1_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2891__CLK (.I(clknet_leaf_2_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2894__CLK (.I(clknet_leaf_2_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2893__CLK (.I(clknet_leaf_2_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2922__CLK (.I(clknet_leaf_2_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2927__CLK (.I(clknet_leaf_2_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2929__CLK (.I(clknet_leaf_2_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2897__CLK (.I(clknet_leaf_2_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2933__CLK (.I(clknet_leaf_2_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2896__CLK (.I(clknet_leaf_2_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2892__CLK (.I(clknet_leaf_2_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2930__CLK (.I(clknet_leaf_2_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2923__CLK (.I(clknet_leaf_2_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3042__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3043__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2888__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2954__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2955__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2889__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2952__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2953__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2957__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3038__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2956__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2966__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3037__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2924__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2926__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2895__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3036__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2890__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3049__CLK (.I(clknet_leaf_4_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3068__CLK (.I(clknet_leaf_4_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3039__CLK (.I(clknet_leaf_4_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3084__CLK (.I(clknet_leaf_4_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3040__CLK (.I(clknet_leaf_4_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2875__CLK (.I(clknet_leaf_4_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3077__CLK (.I(clknet_leaf_4_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3081__CLK (.I(clknet_leaf_4_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3082__CLK (.I(clknet_leaf_4_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2864__CLK (.I(clknet_leaf_4_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3083__CLK (.I(clknet_leaf_4_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2939__CLK (.I(clknet_leaf_4_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3041__CLK (.I(clknet_leaf_4_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2863__CLK (.I(clknet_leaf_4_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2951__CLK (.I(clknet_leaf_4_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2950__CLK (.I(clknet_leaf_4_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3157__CLK (.I(clknet_leaf_5_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3057__CLK (.I(clknet_leaf_5_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3056__CLK (.I(clknet_leaf_5_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3055__CLK (.I(clknet_leaf_5_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3053__CLK (.I(clknet_leaf_5_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3155__CLK (.I(clknet_leaf_5_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3153__CLK (.I(clknet_leaf_5_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3133__CLK (.I(clknet_leaf_5_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3151__CLK (.I(clknet_leaf_5_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3048__CLK (.I(clknet_leaf_5_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2861__CLK (.I(clknet_leaf_5_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3052__CLK (.I(clknet_leaf_5_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3054__CLK (.I(clknet_leaf_5_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3076__CLK (.I(clknet_leaf_5_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2862__CLK (.I(clknet_leaf_5_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3063__CLK (.I(clknet_leaf_6_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3065__CLK (.I(clknet_leaf_6_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3067__CLK (.I(clknet_leaf_6_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2876__CLK (.I(clknet_leaf_6_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3066__CLK (.I(clknet_leaf_6_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3064__CLK (.I(clknet_leaf_6_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3179__CLK (.I(clknet_leaf_6_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3058__CLK (.I(clknet_leaf_6_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3059__CLK (.I(clknet_leaf_6_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3165__CLK (.I(clknet_leaf_6_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3163__CLK (.I(clknet_leaf_6_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3161__CLK (.I(clknet_leaf_6_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3159__CLK (.I(clknet_leaf_6_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2879__CLK (.I(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2878__CLK (.I(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3243__CLK (.I(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3238__CLK (.I(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3237__CLK (.I(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3236__CLK (.I(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3235__CLK (.I(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3239__CLK (.I(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3240__CLK (.I(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3241__CLK (.I(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3061__CLK (.I(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3242__CLK (.I(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3169__CLK (.I(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3177__CLK (.I(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3167__CLK (.I(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3234__CLK (.I(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3181__CLK (.I(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3175__CLK (.I(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3060__CLK (.I(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3171__CLK (.I(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3173__CLK (.I(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3062__CLK (.I(clknet_leaf_8_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2887__CLK (.I(clknet_leaf_8_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2886__CLK (.I(clknet_leaf_8_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2885__CLK (.I(clknet_leaf_8_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2880__CLK (.I(clknet_leaf_8_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2881__CLK (.I(clknet_leaf_8_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2884__CLK (.I(clknet_leaf_8_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2882__CLK (.I(clknet_leaf_8_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3250__CLK (.I(clknet_leaf_8_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3246__CLK (.I(clknet_leaf_8_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3244__CLK (.I(clknet_leaf_8_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3245__CLK (.I(clknet_leaf_8_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3247__CLK (.I(clknet_leaf_8_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3258__I (.I(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3257__I (.I(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3248__CLK (.I(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3255__I (.I(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3256__I (.I(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3251__CLK (.I(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2860__CLK (.I(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3252__CLK (.I(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3254__I (.I(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2834__CLK (.I(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3069__CLK (.I(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3070__CLK (.I(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3071__CLK (.I(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3253__CLK (.I(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2883__CLK (.I(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2972__CLK (.I(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3078__CLK (.I(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3074__CLK (.I(clknet_leaf_10_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3072__CLK (.I(clknet_leaf_10_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3073__CLK (.I(clknet_leaf_10_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2869__CLK (.I(clknet_leaf_10_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2839__CLK (.I(clknet_leaf_10_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2837__CLK (.I(clknet_leaf_10_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2836__CLK (.I(clknet_leaf_10_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2847__CLK (.I(clknet_leaf_10_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2835__CLK (.I(clknet_leaf_10_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2833__CLK (.I(clknet_leaf_10_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2832__CLK (.I(clknet_leaf_10_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3263__I (.I(clknet_leaf_10_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3261__I (.I(clknet_leaf_10_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3262__I (.I(clknet_leaf_10_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3260__I (.I(clknet_leaf_10_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3259__I (.I(clknet_leaf_10_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3249__CLK (.I(clknet_leaf_10_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2971__CLK (.I(clknet_leaf_11_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2973__CLK (.I(clknet_leaf_11_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2974__CLK (.I(clknet_leaf_11_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2975__CLK (.I(clknet_leaf_11_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2976__CLK (.I(clknet_leaf_11_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2978__CLK (.I(clknet_leaf_11_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2977__CLK (.I(clknet_leaf_11_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2868__CLK (.I(clknet_leaf_11_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3075__CLK (.I(clknet_leaf_11_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3005__CLK (.I(clknet_leaf_12_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3007__CLK (.I(clknet_leaf_12_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3006__CLK (.I(clknet_leaf_12_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2949__CLK (.I(clknet_leaf_12_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2948__CLK (.I(clknet_leaf_12_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2938__CLK (.I(clknet_leaf_12_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2877__CLK (.I(clknet_leaf_12_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2970__CLK (.I(clknet_leaf_12_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3079__CLK (.I(clknet_leaf_12_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3080__CLK (.I(clknet_leaf_12_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2940__CLK (.I(clknet_leaf_13_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3017__CLK (.I(clknet_leaf_13_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3020__CLK (.I(clknet_leaf_13_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3021__CLK (.I(clknet_leaf_13_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3018__CLK (.I(clknet_leaf_13_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3019__CLK (.I(clknet_leaf_13_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3004__CLK (.I(clknet_leaf_13_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2872__CLK (.I(clknet_leaf_14_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2870__CLK (.I(clknet_leaf_14_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2979__CLK (.I(clknet_leaf_14_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2983__CLK (.I(clknet_leaf_14_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2980__CLK (.I(clknet_leaf_14_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2943__CLK (.I(clknet_leaf_14_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3008__CLK (.I(clknet_leaf_14_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3016__CLK (.I(clknet_leaf_14_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3015__CLK (.I(clknet_leaf_14_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2942__CLK (.I(clknet_leaf_14_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2941__CLK (.I(clknet_leaf_14_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2850__CLK (.I(clknet_leaf_15_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2846__CLK (.I(clknet_leaf_15_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2857__CLK (.I(clknet_leaf_15_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2843__CLK (.I(clknet_leaf_15_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2842__CLK (.I(clknet_leaf_15_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2845__CLK (.I(clknet_leaf_15_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2851__CLK (.I(clknet_leaf_15_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2841__CLK (.I(clknet_leaf_15_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2844__CLK (.I(clknet_leaf_15_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2840__CLK (.I(clknet_leaf_15_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2838__CLK (.I(clknet_leaf_15_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2871__CLK (.I(clknet_leaf_15_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3224__CLK (.I(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3226__CLK (.I(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3217__CLK (.I(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2995__CLK (.I(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2994__CLK (.I(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2996__CLK (.I(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2985__CLK (.I(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2986__CLK (.I(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2997__CLK (.I(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2981__CLK (.I(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3009__CLK (.I(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2854__CLK (.I(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2982__CLK (.I(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2848__CLK (.I(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2852__CLK (.I(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2859__CLK (.I(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2874__CLK (.I(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2873__CLK (.I(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2858__CLK (.I(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2853__CLK (.I(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2849__CLK (.I(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2855__CLK (.I(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2856__CLK (.I(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3233__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2990__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2991__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3223__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3219__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3218__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3221__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3215__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3220__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3214__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3231__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3230__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3232__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3001__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3228__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3216__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3225__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3227__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2987__CLK (.I(clknet_leaf_18_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2998__CLK (.I(clknet_leaf_18_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2999__CLK (.I(clknet_leaf_18_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3000__CLK (.I(clknet_leaf_18_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3229__CLK (.I(clknet_leaf_18_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2984__CLK (.I(clknet_leaf_18_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3003__CLK (.I(clknet_leaf_18_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3002__CLK (.I(clknet_leaf_18_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2992__CLK (.I(clknet_leaf_18_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3222__CLK (.I(clknet_leaf_18_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2993__CLK (.I(clknet_leaf_18_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2989__CLK (.I(clknet_leaf_18_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2988__CLK (.I(clknet_leaf_18_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2944__CLK (.I(clknet_leaf_19_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2946__CLK (.I(clknet_leaf_19_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3013__CLK (.I(clknet_leaf_19_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3012__CLK (.I(clknet_leaf_19_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2945__CLK (.I(clknet_leaf_19_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3011__CLK (.I(clknet_leaf_19_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3010__CLK (.I(clknet_leaf_19_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3025__CLK (.I(clknet_leaf_20_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3027__CLK (.I(clknet_leaf_20_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2963__CLK (.I(clknet_leaf_20_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3026__CLK (.I(clknet_leaf_20_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2960__CLK (.I(clknet_leaf_20_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2959__CLK (.I(clknet_leaf_20_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2958__CLK (.I(clknet_leaf_20_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2947__CLK (.I(clknet_leaf_20_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2962__CLK (.I(clknet_leaf_20_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3023__CLK (.I(clknet_leaf_21_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3014__CLK (.I(clknet_leaf_21_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3024__CLK (.I(clknet_leaf_21_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3032__CLK (.I(clknet_leaf_21_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2961__CLK (.I(clknet_leaf_21_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3035__CLK (.I(clknet_leaf_22_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3033__CLK (.I(clknet_leaf_22_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3034__CLK (.I(clknet_leaf_22_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2909__CLK (.I(clknet_leaf_22_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2908__CLK (.I(clknet_leaf_22_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2968__CLK (.I(clknet_leaf_22_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2969__CLK (.I(clknet_leaf_22_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2967__CLK (.I(clknet_leaf_23_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3195__CLK (.I(clknet_leaf_23_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3197__CLK (.I(clknet_leaf_23_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3198__CLK (.I(clknet_leaf_23_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3090__CLK (.I(clknet_leaf_23_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3202__CLK (.I(clknet_leaf_23_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3201__CLK (.I(clknet_leaf_23_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3203__CLK (.I(clknet_leaf_23_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3205__CLK (.I(clknet_leaf_23_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3204__CLK (.I(clknet_leaf_23_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3191__CLK (.I(clknet_leaf_23_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2912__CLK (.I(clknet_leaf_24_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2910__CLK (.I(clknet_leaf_24_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2911__CLK (.I(clknet_leaf_24_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3029__CLK (.I(clknet_leaf_24_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3030__CLK (.I(clknet_leaf_24_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3028__CLK (.I(clknet_leaf_24_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2964__CLK (.I(clknet_leaf_24_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2965__CLK (.I(clknet_leaf_24_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3196__CLK (.I(clknet_leaf_24_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3031__CLK (.I(clknet_leaf_24_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3092__CLK (.I(clknet_leaf_25_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3091__CLK (.I(clknet_leaf_25_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2914__CLK (.I(clknet_leaf_25_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2913__CLK (.I(clknet_leaf_25_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2916__CLK (.I(clknet_leaf_26_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2915__CLK (.I(clknet_leaf_26_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2917__CLK (.I(clknet_leaf_26_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3097__CLK (.I(clknet_leaf_26_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3094__CLK (.I(clknet_leaf_26_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3093__CLK (.I(clknet_leaf_26_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3095__CLK (.I(clknet_leaf_26_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3098__CLK (.I(clknet_leaf_27_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2918__CLK (.I(clknet_leaf_27_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2919__CLK (.I(clknet_leaf_27_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3096__CLK (.I(clknet_leaf_27_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2920__CLK (.I(clknet_leaf_28_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3102__CLK (.I(clknet_leaf_28_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3101__CLK (.I(clknet_leaf_28_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3183__CLK (.I(clknet_leaf_28_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3209__CLK (.I(clknet_leaf_28_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3087__CLK (.I(clknet_leaf_29_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3088__CLK (.I(clknet_leaf_29_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3089__CLK (.I(clknet_leaf_29_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3206__CLK (.I(clknet_leaf_29_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3099__CLK (.I(clknet_leaf_29_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3100__CLK (.I(clknet_leaf_29_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2921__CLK (.I(clknet_leaf_29_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3086__CLK (.I(clknet_leaf_29_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3104__CLK (.I(clknet_leaf_30_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3194__CLK (.I(clknet_leaf_30_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2925__CLK (.I(clknet_leaf_30_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2906__CLK (.I(clknet_leaf_30_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2907__CLK (.I(clknet_leaf_30_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3022__CLK (.I(clknet_leaf_30_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3193__CLK (.I(clknet_leaf_30_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3192__CLK (.I(clknet_leaf_30_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3107__CLK (.I(clknet_leaf_31_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3109__CLK (.I(clknet_leaf_31_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3108__CLK (.I(clknet_leaf_31_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3106__CLK (.I(clknet_leaf_31_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3199__CLK (.I(clknet_leaf_31_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3200__CLK (.I(clknet_leaf_31_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2928__CLK (.I(clknet_leaf_31_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3105__CLK (.I(clknet_leaf_31_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3182__CLK (.I(clknet_leaf_32_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2867__CLK (.I(clknet_leaf_32_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3213__CLK (.I(clknet_leaf_32_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3103__CLK (.I(clknet_leaf_32_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3110__CLK (.I(clknet_leaf_33_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2865__CLK (.I(clknet_leaf_33_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3211__CLK (.I(clknet_leaf_33_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3188__CLK (.I(clknet_leaf_33_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3187__CLK (.I(clknet_leaf_33_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3186__CLK (.I(clknet_leaf_33_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3185__CLK (.I(clknet_leaf_33_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3184__CLK (.I(clknet_leaf_33_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2866__CLK (.I(clknet_leaf_34_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3212__CLK (.I(clknet_leaf_34_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3111__CLK (.I(clknet_leaf_34_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3112__CLK (.I(clknet_leaf_34_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3113__CLK (.I(clknet_leaf_34_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2901__CLK (.I(clknet_leaf_34_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2900__CLK (.I(clknet_leaf_34_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3210__CLK (.I(clknet_leaf_35_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3208__CLK (.I(clknet_leaf_35_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3085__CLK (.I(clknet_leaf_35_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3119__CLK (.I(clknet_leaf_35_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3121__CLK (.I(clknet_leaf_35_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3190__CLK (.I(clknet_leaf_35_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3207__CLK (.I(clknet_leaf_35_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3189__CLK (.I(clknet_leaf_35_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3114__CLK (.I(clknet_leaf_36_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2902__CLK (.I(clknet_leaf_36_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2904__CLK (.I(clknet_leaf_36_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2903__CLK (.I(clknet_leaf_36_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3117__CLK (.I(clknet_leaf_36_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3116__CLK (.I(clknet_leaf_36_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2899__CLK (.I(clknet_leaf_36_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3127__CLK (.I(clknet_leaf_36_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3115__CLK (.I(clknet_leaf_36_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3123__CLK (.I(clknet_leaf_36_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3125__CLK (.I(clknet_leaf_36_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_3__f_clock_I (.I(clknet_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_2__f_clock_I (.I(clknet_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_1__f_clock_I (.I(clknet_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_0__f_clock_I (.I(clknet_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2932__CLK (.I(clknet_2_0__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_36_clock_I (.I(clknet_2_0__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_35_clock_I (.I(clknet_2_0__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_34_clock_I (.I(clknet_2_0__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_33_clock_I (.I(clknet_2_0__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_32_clock_I (.I(clknet_2_0__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_31_clock_I (.I(clknet_2_0__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_30_clock_I (.I(clknet_2_0__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_2_clock_I (.I(clknet_2_0__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_1_clock_I (.I(clknet_2_0__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_0_clock_I (.I(clknet_2_0__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_13_clock_I (.I(clknet_2_1__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_12_clock_I (.I(clknet_2_1__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_11_clock_I (.I(clknet_2_1__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_10_clock_I (.I(clknet_2_1__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_9_clock_I (.I(clknet_2_1__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_8_clock_I (.I(clknet_2_1__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_7_clock_I (.I(clknet_2_1__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_6_clock_I (.I(clknet_2_1__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_5_clock_I (.I(clknet_2_1__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_4_clock_I (.I(clknet_2_1__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_3_clock_I (.I(clknet_2_1__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_29_clock_I (.I(clknet_2_2__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_28_clock_I (.I(clknet_2_2__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_27_clock_I (.I(clknet_2_2__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_26_clock_I (.I(clknet_2_2__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_25_clock_I (.I(clknet_2_2__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_24_clock_I (.I(clknet_2_2__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_23_clock_I (.I(clknet_2_2__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_22_clock_I (.I(clknet_2_2__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_21_clock_I (.I(clknet_2_3__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_20_clock_I (.I(clknet_2_3__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_19_clock_I (.I(clknet_2_3__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_18_clock_I (.I(clknet_2_3__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_17_clock_I (.I(clknet_2_3__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_16_clock_I (.I(clknet_2_3__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_15_clock_I (.I(clknet_2_3__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_14_clock_I (.I(clknet_2_3__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2861__D (.I(net243));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3248__D (.I(net247));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2860__D (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2863__D (.I(net250));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3232__D (.I(net266));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3220__D (.I(net281));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3221__D (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2847__D (.I(net288));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2849__D (.I(net289));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2848__D (.I(net290));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1399 ();
endmodule


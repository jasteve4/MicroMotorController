// This is the unpowered netlist.
module spi_core (clock,
    clock_out,
    miso,
    miso_oeb,
    mosi,
    mosi_oeb,
    sclk,
    sclk_oeb,
    ss_n,
    ss_n_oeb,
    data_out,
    la_data_in,
    la_oenb);
 input clock;
 output clock_out;
 output miso;
 output miso_oeb;
 input mosi;
 output mosi_oeb;
 input sclk;
 output sclk_oeb;
 input ss_n;
 output ss_n_oeb;
 output [31:0] data_out;
 input [3:0] la_data_in;
 output [3:0] la_oenb;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire clknet_0_clock;
 wire net43;
 wire \mosi_reg[0] ;
 wire \mosi_reg[1] ;
 wire \mosi_reg[2] ;
 wire net44;
 wire \sclk_reg[0] ;
 wire \sclk_reg[1] ;
 wire \sclk_reg[2] ;
 wire net45;
 wire \ss_n_reg[0] ;
 wire \ss_n_reg[1] ;
 wire \ss_n_reg[2] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire clknet_2_0__leaf_clock;
 wire clknet_2_1__leaf_clock;
 wire clknet_2_2__leaf_clock;
 wire clknet_2_3__leaf_clock;

 gf180mcu_fd_sc_mcu7t5v0__and2_1 _078_ (.A1(\mosi_reg[2] ),
    .A2(\mosi_reg[1] ),
    .Z(_059_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _079_ (.I(\sclk_reg[2] ),
    .ZN(_060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _080_ (.A1(\ss_n_reg[2] ),
    .A2(\ss_n_reg[1] ),
    .ZN(_061_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _081_ (.A1(_060_),
    .A2(\sclk_reg[1] ),
    .A3(_061_),
    .ZN(_062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _082_ (.I(_062_),
    .Z(_063_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _083_ (.I(_063_),
    .Z(_064_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _084_ (.I0(_059_),
    .I1(net5),
    .S(_064_),
    .Z(_065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _085_ (.I(_065_),
    .Z(_000_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _086_ (.I0(net5),
    .I1(net16),
    .S(_064_),
    .Z(_066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _087_ (.I(_066_),
    .Z(_001_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _088_ (.I0(net16),
    .I1(net27),
    .S(_064_),
    .Z(_067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _089_ (.I(_067_),
    .Z(_002_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _090_ (.I0(net27),
    .I1(net30),
    .S(_064_),
    .Z(_068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _091_ (.I(_068_),
    .Z(_003_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _092_ (.I(_063_),
    .Z(_069_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _093_ (.I0(net30),
    .I1(net31),
    .S(_069_),
    .Z(_070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _094_ (.I(_070_),
    .Z(_004_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _095_ (.I0(net31),
    .I1(net32),
    .S(_069_),
    .Z(_071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _096_ (.I(_071_),
    .Z(_005_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _097_ (.I0(net32),
    .I1(net33),
    .S(_069_),
    .Z(_072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _098_ (.I(_072_),
    .Z(_006_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _099_ (.I0(net33),
    .I1(net34),
    .S(_069_),
    .Z(_073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _100_ (.I(_073_),
    .Z(_007_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _101_ (.I(_063_),
    .Z(_074_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _102_ (.I0(net34),
    .I1(net35),
    .S(_074_),
    .Z(_075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _103_ (.I(_075_),
    .Z(_008_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _104_ (.I0(net35),
    .I1(net36),
    .S(_074_),
    .Z(_076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _105_ (.I(_076_),
    .Z(_009_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _106_ (.I0(net36),
    .I1(net6),
    .S(_074_),
    .Z(_077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _107_ (.I(_077_),
    .Z(_010_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _108_ (.I0(net6),
    .I1(net7),
    .S(_074_),
    .Z(_032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _109_ (.I(_032_),
    .Z(_011_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _110_ (.I(_063_),
    .Z(_033_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _111_ (.I0(net7),
    .I1(net8),
    .S(_033_),
    .Z(_034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _112_ (.I(_034_),
    .Z(_012_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _113_ (.I0(net8),
    .I1(net9),
    .S(_033_),
    .Z(_035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _114_ (.I(_035_),
    .Z(_013_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _115_ (.I0(net9),
    .I1(net10),
    .S(_033_),
    .Z(_036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _116_ (.I(_036_),
    .Z(_014_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _117_ (.I0(net10),
    .I1(net11),
    .S(_033_),
    .Z(_037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _118_ (.I(_037_),
    .Z(_015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _119_ (.I(_062_),
    .Z(_038_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _120_ (.I(_038_),
    .Z(_039_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _121_ (.I0(net11),
    .I1(net12),
    .S(_039_),
    .Z(_040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _122_ (.I(_040_),
    .Z(_016_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _123_ (.I0(net12),
    .I1(net13),
    .S(_039_),
    .Z(_041_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _124_ (.I(_041_),
    .Z(_017_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _125_ (.I0(net13),
    .I1(net14),
    .S(_039_),
    .Z(_042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _126_ (.I(_042_),
    .Z(_018_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _127_ (.I0(net14),
    .I1(net15),
    .S(_039_),
    .Z(_043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _128_ (.I(_043_),
    .Z(_019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _129_ (.I(_038_),
    .Z(_044_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _130_ (.I0(net15),
    .I1(net17),
    .S(_044_),
    .Z(_045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _131_ (.I(_045_),
    .Z(_020_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _132_ (.I0(net17),
    .I1(net18),
    .S(_044_),
    .Z(_046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _133_ (.I(_046_),
    .Z(_021_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _134_ (.I0(net18),
    .I1(net19),
    .S(_044_),
    .Z(_047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _135_ (.I(_047_),
    .Z(_022_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _136_ (.I0(net19),
    .I1(net20),
    .S(_044_),
    .Z(_048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _137_ (.I(_048_),
    .Z(_023_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _138_ (.I(_038_),
    .Z(_049_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _139_ (.I0(net20),
    .I1(net21),
    .S(_049_),
    .Z(_050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _140_ (.I(_050_),
    .Z(_024_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _141_ (.I0(net21),
    .I1(net22),
    .S(_049_),
    .Z(_051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _142_ (.I(_051_),
    .Z(_025_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _143_ (.I0(net22),
    .I1(net23),
    .S(_049_),
    .Z(_052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _144_ (.I(_052_),
    .Z(_026_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _145_ (.I0(net23),
    .I1(net24),
    .S(_049_),
    .Z(_053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _146_ (.I(_053_),
    .Z(_027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _147_ (.I(_038_),
    .Z(_054_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _148_ (.I0(net24),
    .I1(net25),
    .S(_054_),
    .Z(_055_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _149_ (.I(_055_),
    .Z(_028_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _150_ (.I0(net25),
    .I1(net26),
    .S(_054_),
    .Z(_056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _151_ (.I(_056_),
    .Z(_029_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _152_ (.I0(net26),
    .I1(net28),
    .S(_054_),
    .Z(_057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _153_ (.I(_057_),
    .Z(_030_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _154_ (.I0(net28),
    .I1(net29),
    .S(_054_),
    .Z(_058_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _155_ (.I(_058_),
    .Z(_031_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _156_ (.D(net1),
    .CLK(clknet_2_1__leaf_clock),
    .Q(\mosi_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _157_ (.D(\mosi_reg[0] ),
    .CLK(clknet_2_0__leaf_clock),
    .Q(\mosi_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _158_ (.D(\mosi_reg[1] ),
    .CLK(clknet_2_0__leaf_clock),
    .Q(\mosi_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _159_ (.D(net3),
    .CLK(clknet_2_1__leaf_clock),
    .Q(\ss_n_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _160_ (.D(\ss_n_reg[0] ),
    .CLK(clknet_2_0__leaf_clock),
    .Q(\ss_n_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _161_ (.D(\ss_n_reg[1] ),
    .CLK(clknet_2_1__leaf_clock),
    .Q(\ss_n_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _162_ (.D(net2),
    .CLK(clknet_2_1__leaf_clock),
    .Q(\sclk_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _163_ (.D(\sclk_reg[0] ),
    .CLK(clknet_2_0__leaf_clock),
    .Q(\sclk_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _164_ (.D(\sclk_reg[1] ),
    .CLK(clknet_2_0__leaf_clock),
    .Q(\sclk_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _165_ (.D(_000_),
    .CLK(clknet_2_2__leaf_clock),
    .Q(net5));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _166_ (.D(_001_),
    .CLK(clknet_2_2__leaf_clock),
    .Q(net16));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _167_ (.D(_002_),
    .CLK(clknet_2_2__leaf_clock),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _168_ (.D(_003_),
    .CLK(clknet_2_2__leaf_clock),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _169_ (.D(_004_),
    .CLK(clknet_2_2__leaf_clock),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _170_ (.D(_005_),
    .CLK(clknet_2_2__leaf_clock),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _171_ (.D(_006_),
    .CLK(clknet_2_3__leaf_clock),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _172_ (.D(_007_),
    .CLK(clknet_2_3__leaf_clock),
    .Q(net34));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _173_ (.D(_008_),
    .CLK(clknet_2_3__leaf_clock),
    .Q(net35));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _174_ (.D(_009_),
    .CLK(clknet_2_3__leaf_clock),
    .Q(net36));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _175_ (.D(_010_),
    .CLK(clknet_2_3__leaf_clock),
    .Q(net6));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _176_ (.D(_011_),
    .CLK(clknet_2_3__leaf_clock),
    .Q(net7));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _177_ (.D(_012_),
    .CLK(clknet_2_2__leaf_clock),
    .Q(net8));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _178_ (.D(_013_),
    .CLK(clknet_2_2__leaf_clock),
    .Q(net9));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _179_ (.D(_014_),
    .CLK(clknet_2_2__leaf_clock),
    .Q(net10));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _180_ (.D(_015_),
    .CLK(clknet_2_2__leaf_clock),
    .Q(net11));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _181_ (.D(_016_),
    .CLK(clknet_2_2__leaf_clock),
    .Q(net12));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _182_ (.D(_017_),
    .CLK(clknet_2_0__leaf_clock),
    .Q(net13));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _183_ (.D(_018_),
    .CLK(clknet_2_0__leaf_clock),
    .Q(net14));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _184_ (.D(_019_),
    .CLK(clknet_2_1__leaf_clock),
    .Q(net15));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _185_ (.D(_020_),
    .CLK(clknet_2_1__leaf_clock),
    .Q(net17));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _186_ (.D(_021_),
    .CLK(clknet_2_1__leaf_clock),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _187_ (.D(_022_),
    .CLK(clknet_2_1__leaf_clock),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _188_ (.D(_023_),
    .CLK(clknet_2_1__leaf_clock),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _189_ (.D(_024_),
    .CLK(clknet_2_3__leaf_clock),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _190_ (.D(_025_),
    .CLK(clknet_2_3__leaf_clock),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _191_ (.D(_026_),
    .CLK(clknet_2_3__leaf_clock),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _192_ (.D(_027_),
    .CLK(clknet_2_3__leaf_clock),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _193_ (.D(_028_),
    .CLK(clknet_2_3__leaf_clock),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _194_ (.D(_029_),
    .CLK(clknet_2_3__leaf_clock),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _195_ (.D(_030_),
    .CLK(clknet_2_3__leaf_clock),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _196_ (.D(_031_),
    .CLK(clknet_2_1__leaf_clock),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_clock (.I(clock),
    .Z(clknet_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__tiel spi_core_39 (.ZN(net39));
 gf180mcu_fd_sc_mcu7t5v0__tiel spi_core_40 (.ZN(net40));
 gf180mcu_fd_sc_mcu7t5v0__tiel spi_core_41 (.ZN(net41));
 gf180mcu_fd_sc_mcu7t5v0__tiel spi_core_42 (.ZN(net42));
 gf180mcu_fd_sc_mcu7t5v0__tiel spi_core_43 (.ZN(net43));
 gf180mcu_fd_sc_mcu7t5v0__tiel spi_core_44 (.ZN(net44));
 gf180mcu_fd_sc_mcu7t5v0__tieh spi_core_45 (.Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _205_ (.I(clknet_2_2__leaf_clock),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _206_ (.I(net29),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(mosi),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(sclk),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(ss_n),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output4 (.I(net4),
    .Z(clock_out));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output5 (.I(net5),
    .Z(data_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output6 (.I(net6),
    .Z(data_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output7 (.I(net7),
    .Z(data_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output8 (.I(net8),
    .Z(data_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output9 (.I(net9),
    .Z(data_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output10 (.I(net10),
    .Z(data_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output11 (.I(net11),
    .Z(data_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output12 (.I(net12),
    .Z(data_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output13 (.I(net13),
    .Z(data_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output14 (.I(net14),
    .Z(data_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output15 (.I(net15),
    .Z(data_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output16 (.I(net16),
    .Z(data_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output17 (.I(net17),
    .Z(data_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output18 (.I(net18),
    .Z(data_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output19 (.I(net19),
    .Z(data_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output20 (.I(net20),
    .Z(data_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output21 (.I(net21),
    .Z(data_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output22 (.I(net22),
    .Z(data_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output23 (.I(net23),
    .Z(data_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output24 (.I(net24),
    .Z(data_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output25 (.I(net25),
    .Z(data_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output26 (.I(net26),
    .Z(data_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output27 (.I(net27),
    .Z(data_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output28 (.I(net28),
    .Z(data_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output29 (.I(net29),
    .Z(data_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output30 (.I(net30),
    .Z(data_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output31 (.I(net31),
    .Z(data_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output32 (.I(net32),
    .Z(data_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output33 (.I(net33),
    .Z(data_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output34 (.I(net34),
    .Z(data_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output35 (.I(net35),
    .Z(data_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output36 (.I(net36),
    .Z(data_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output37 (.I(net37),
    .Z(miso));
 gf180mcu_fd_sc_mcu7t5v0__tiel spi_core_38 (.ZN(net38));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_0__f_clock (.I(clknet_0_clock),
    .Z(clknet_2_0__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_1__f_clock (.I(clknet_0_clock),
    .Z(clknet_2_1__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_2__f_clock (.I(clknet_0_clock),
    .Z(clknet_2_2__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_3__f_clock (.I(clknet_0_clock),
    .Z(clknet_2_3__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__165__D (.I(_000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__167__D (.I(_002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__169__D (.I(_004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__170__D (.I(_005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__174__D (.I(_009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__175__D (.I(_010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__176__D (.I(_011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__177__D (.I(_012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__178__D (.I(_013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__179__D (.I(_014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__180__D (.I(_015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__181__D (.I(_016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__182__D (.I(_017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__183__D (.I(_018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__184__D (.I(_019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__185__D (.I(_020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__186__D (.I(_021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__187__D (.I(_022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__188__D (.I(_023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__189__D (.I(_024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__196__D (.I(_031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__127__S (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__125__S (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__123__S (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__121__S (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__137__I (.I(_048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__140__I (.I(_050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__142__I (.I(_051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__144__I (.I(_052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__146__I (.I(_053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__154__S (.I(_054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__152__S (.I(_054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__150__S (.I(_054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__148__S (.I(_054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__149__I (.I(_055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__151__I (.I(_056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__153__I (.I(_057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__090__S (.I(_064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__088__S (.I(_064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__086__S (.I(_064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__084__S (.I(_064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_clock_I (.I(clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_3__f_clock_I (.I(clknet_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_2__f_clock_I (.I(clknet_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_1__f_clock_I (.I(clknet_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_0__f_clock_I (.I(clknet_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(mosi));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__158__D (.I(\mosi_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__078__A2 (.I(\mosi_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__078__A1 (.I(\mosi_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(sclk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__164__D (.I(\sclk_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__081__A2 (.I(\sclk_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__079__I (.I(\sclk_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(ss_n));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__161__D (.I(\ss_n_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__080__A2 (.I(\ss_n_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__080__A1 (.I(\ss_n_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__156__D (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__159__D (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output4_I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output5_I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__086__I0 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__084__I1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output6_I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__108__I0 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__106__I1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output7_I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__111__I0 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__108__I1 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output8_I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__113__I0 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__111__I1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output9_I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__115__I0 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__113__I1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output10_I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__117__I0 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__115__I1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output11_I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__121__I0 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__117__I1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output12_I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__123__I0 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__121__I1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output13_I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__125__I0 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__123__I1 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output14_I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__127__I0 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__125__I1 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output15_I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__130__I0 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__127__I1 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output16_I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__088__I0 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__086__I1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output17_I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__132__I0 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__130__I1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output18_I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__134__I0 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__132__I1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output19_I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__136__I0 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__134__I1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output20_I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__139__I0 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__136__I1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output21_I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__141__I0 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__139__I1 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output22_I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__143__I0 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__141__I1 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output23_I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__145__I0 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__143__I1 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output24_I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__148__I0 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__145__I1 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output25_I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__150__I0 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__148__I1 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output26_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__152__I0 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__150__I1 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output27_I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__090__I0 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__088__I1 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output28_I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__154__I0 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__152__I1 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output29_I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__206__I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__154__I1 (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output30_I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__093__I0 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__090__I1 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output31_I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__095__I0 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__093__I1 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output32_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__097__I0 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__095__I1 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output33_I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__099__I0 (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__097__I1 (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output34_I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__102__I0 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__099__I1 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output35_I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__104__I0 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__102__I1 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output36_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__106__I0 (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__104__I1 (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output37_I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__157__CLK (.I(clknet_2_0__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__158__CLK (.I(clknet_2_0__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__160__CLK (.I(clknet_2_0__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__163__CLK (.I(clknet_2_0__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__164__CLK (.I(clknet_2_0__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__182__CLK (.I(clknet_2_0__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__183__CLK (.I(clknet_2_0__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__156__CLK (.I(clknet_2_1__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__159__CLK (.I(clknet_2_1__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__161__CLK (.I(clknet_2_1__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__162__CLK (.I(clknet_2_1__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__184__CLK (.I(clknet_2_1__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__185__CLK (.I(clknet_2_1__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__186__CLK (.I(clknet_2_1__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__187__CLK (.I(clknet_2_1__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__188__CLK (.I(clknet_2_1__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__196__CLK (.I(clknet_2_1__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__165__CLK (.I(clknet_2_2__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__166__CLK (.I(clknet_2_2__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__167__CLK (.I(clknet_2_2__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__168__CLK (.I(clknet_2_2__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__169__CLK (.I(clknet_2_2__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__170__CLK (.I(clknet_2_2__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__177__CLK (.I(clknet_2_2__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__178__CLK (.I(clknet_2_2__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__179__CLK (.I(clknet_2_2__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__180__CLK (.I(clknet_2_2__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__181__CLK (.I(clknet_2_2__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__205__I (.I(clknet_2_2__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__171__CLK (.I(clknet_2_3__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__172__CLK (.I(clknet_2_3__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__173__CLK (.I(clknet_2_3__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__174__CLK (.I(clknet_2_3__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__175__CLK (.I(clknet_2_3__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__176__CLK (.I(clknet_2_3__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__189__CLK (.I(clknet_2_3__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__190__CLK (.I(clknet_2_3__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__191__CLK (.I(clknet_2_3__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__192__CLK (.I(clknet_2_3__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__193__CLK (.I(clknet_2_3__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__194__CLK (.I(clknet_2_3__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__195__CLK (.I(clknet_2_3__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_419 ();
 assign la_oenb[0] = net38;
 assign la_oenb[1] = net39;
 assign la_oenb[2] = net40;
 assign la_oenb[3] = net41;
 assign miso_oeb = net45;
 assign mosi_oeb = net42;
 assign sclk_oeb = net43;
 assign ss_n_oeb = net44;
endmodule


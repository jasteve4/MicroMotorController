magic
tech gf180mcuC
magscale 1 10
timestamp 1670301642
<< metal1 >>
rect 398626 158398 398638 158450
rect 398690 158447 398702 158450
rect 399074 158447 399086 158450
rect 398690 158401 399086 158447
rect 398690 158398 398702 158401
rect 399074 158398 399086 158401
rect 399138 158398 399150 158450
rect 399522 158111 399534 158114
rect 399313 158065 399534 158111
rect 399313 158002 399359 158065
rect 399522 158062 399534 158065
rect 399586 158062 399598 158114
rect 399298 157950 399310 158002
rect 399362 157950 399374 158002
rect 399746 157999 399758 158002
rect 399537 157953 399758 157999
rect 399537 157890 399583 157953
rect 399746 157950 399758 157953
rect 399810 157950 399822 158002
rect 399522 157838 399534 157890
rect 399586 157838 399598 157890
rect 60722 29374 60734 29426
rect 60786 29423 60798 29426
rect 61058 29423 61070 29426
rect 60786 29377 61070 29423
rect 60786 29374 60798 29377
rect 61058 29374 61070 29377
rect 61122 29374 61134 29426
rect 60722 27134 60734 27186
rect 60786 27183 60798 27186
rect 61954 27183 61966 27186
rect 60786 27137 61966 27183
rect 60786 27134 60798 27137
rect 61954 27134 61966 27137
rect 62018 27134 62030 27186
rect 60722 23662 60734 23714
rect 60786 23711 60798 23714
rect 61058 23711 61070 23714
rect 60786 23665 61070 23711
rect 60786 23662 60798 23665
rect 61058 23662 61070 23665
rect 61122 23662 61134 23714
<< via1 >>
rect 398638 158398 398690 158450
rect 399086 158398 399138 158450
rect 399534 158062 399586 158114
rect 399310 157950 399362 158002
rect 399758 157950 399810 158002
rect 399534 157838 399586 157890
rect 60734 29374 60786 29426
rect 61070 29374 61122 29426
rect 60734 27134 60786 27186
rect 61966 27134 62018 27186
rect 60734 23662 60786 23714
rect 61070 23662 61122 23714
<< metal2 >>
rect 9688 591640 9912 593000
rect 26040 591640 26264 593000
rect 9688 591560 9940 591640
rect 9884 587972 9940 591560
rect 9884 587906 9940 587916
rect 26012 591560 26264 591640
rect 42392 591560 42616 593000
rect 58744 591560 58968 593000
rect 75096 591640 75320 593000
rect 91448 591640 91672 593000
rect 75068 591560 75320 591640
rect 91420 591560 91672 591640
rect 107800 591560 108024 593000
rect 124152 591560 124376 593000
rect 140504 591640 140728 593000
rect 156856 591640 157080 593000
rect 140504 591560 140756 591640
rect 156856 591560 157108 591640
rect 173208 591560 173432 593000
rect 189560 591560 189784 593000
rect 205912 591640 206136 593000
rect 222264 591640 222488 593000
rect 205884 591560 206136 591640
rect 222236 591560 222488 591640
rect 238616 591560 238840 593000
rect 254968 591560 255192 593000
rect 271320 591560 271544 593000
rect 287672 591560 287896 593000
rect 304024 591560 304248 593000
rect 320376 591560 320600 593000
rect 336728 591560 336952 593000
rect 353080 591560 353304 593000
rect 369432 591560 369656 593000
rect 385784 591560 386008 593000
rect 402136 591640 402360 593000
rect 402108 591560 402360 591640
rect 418488 591560 418712 593000
rect 434840 591560 435064 593000
rect 451192 591560 451416 593000
rect 467544 591640 467768 593000
rect 467516 591560 467768 591640
rect 483896 591560 484120 593000
rect 500248 591560 500472 593000
rect 516600 591560 516824 593000
rect 532588 591612 532868 591668
rect 532952 591640 533176 593000
rect 3276 587412 3332 587422
rect 3164 320964 3220 320974
rect 2492 268884 2548 268894
rect 28 225204 84 225214
rect 28 47124 84 225148
rect 28 47058 84 47068
rect 2492 21924 2548 268828
rect 2604 181860 2660 181870
rect 2604 35364 2660 181804
rect 3164 157332 3220 320908
rect 3276 319284 3332 587356
rect 26012 587412 26068 591560
rect 26012 587346 26068 587356
rect 8316 587300 8372 587310
rect 7532 507780 7588 507790
rect 5852 475188 5908 475198
rect 3388 431844 3444 431854
rect 3388 321076 3444 431788
rect 3388 321010 3444 321020
rect 4172 420868 4228 420878
rect 3276 319218 3332 319228
rect 3164 157266 3220 157276
rect 2604 35298 2660 35308
rect 3276 75684 3332 75694
rect 2492 21858 2548 21868
rect 3276 19460 3332 75628
rect 3276 19394 3332 19404
rect 4172 12852 4228 420812
rect 4172 12786 4228 12796
rect 4284 388276 4340 388286
rect 4284 8260 4340 388220
rect 4396 377412 4452 377422
rect 4396 70868 4452 377356
rect 4396 70802 4452 70812
rect 4508 344820 4564 344830
rect 4508 8372 4564 344764
rect 4732 333956 4788 333966
rect 4620 290500 4676 290510
rect 4620 18004 4676 290444
rect 4732 68964 4788 333900
rect 4844 301364 4900 301374
rect 4844 70756 4900 301308
rect 5852 159684 5908 475132
rect 6636 316708 6692 316718
rect 6524 310100 6580 310110
rect 6412 303268 6468 303278
rect 6300 301588 6356 301598
rect 5852 159618 5908 159628
rect 6076 160132 6132 160142
rect 4844 70690 4900 70700
rect 4956 79044 5012 79054
rect 4732 68898 4788 68908
rect 4956 21476 5012 78988
rect 6076 40516 6132 160076
rect 6300 157668 6356 301532
rect 6300 157602 6356 157612
rect 6412 155428 6468 303212
rect 6524 159572 6580 310044
rect 6524 159506 6580 159516
rect 6412 155362 6468 155372
rect 6636 148708 6692 316652
rect 7420 301812 7476 301822
rect 7420 157780 7476 301756
rect 7420 157714 7476 157724
rect 6636 148642 6692 148652
rect 6076 40450 6132 40460
rect 6524 74004 6580 74014
rect 4956 21410 5012 21420
rect 6524 21364 6580 73948
rect 6524 21298 6580 21308
rect 6636 72436 6692 72446
rect 6636 20020 6692 72380
rect 6636 19954 6692 19964
rect 7532 19796 7588 507724
rect 7868 464324 7924 464334
rect 7644 313572 7700 313582
rect 7644 159460 7700 313516
rect 7644 159394 7700 159404
rect 7756 310212 7812 310222
rect 7756 152852 7812 310156
rect 7756 152786 7812 152796
rect 7532 19730 7588 19740
rect 4620 17938 4676 17948
rect 7868 16548 7924 464268
rect 8204 317156 8260 317166
rect 8092 317044 8148 317054
rect 7980 316932 8036 316942
rect 7980 157444 8036 316876
rect 7980 157378 8036 157388
rect 8092 156996 8148 316988
rect 8092 156930 8148 156940
rect 8204 154196 8260 317100
rect 8204 154130 8260 154140
rect 8316 21140 8372 587244
rect 75068 587300 75124 591560
rect 75068 587234 75124 587244
rect 9996 587188 10052 587198
rect 9996 319172 10052 587132
rect 91420 587188 91476 591560
rect 91420 587122 91476 587132
rect 140700 587188 140756 591560
rect 157052 587300 157108 591560
rect 205884 587524 205940 591560
rect 205884 587458 205940 587468
rect 196476 587412 196532 587422
rect 157052 587234 157108 587244
rect 188972 587300 189028 587310
rect 140700 587122 140756 587132
rect 13244 319284 13300 320040
rect 13244 319218 13300 319228
rect 9996 319106 10052 319116
rect 17052 319172 17108 320040
rect 17052 319106 17108 319116
rect 20188 320012 20888 320068
rect 23548 320012 24696 320068
rect 26908 320012 28504 320068
rect 9660 317380 9716 317390
rect 9548 309988 9604 309998
rect 9436 303492 9492 303502
rect 9100 301700 9156 301710
rect 9100 157892 9156 301644
rect 9100 157826 9156 157836
rect 9212 247044 9268 247054
rect 9212 30212 9268 246988
rect 9324 203588 9380 203598
rect 9324 54852 9380 203532
rect 9436 157556 9492 303436
rect 9548 158788 9604 309932
rect 9660 159236 9716 317324
rect 9772 317268 9828 317278
rect 9772 159348 9828 317212
rect 9996 313796 10052 313806
rect 9772 159282 9828 159292
rect 9884 313684 9940 313694
rect 9660 159170 9716 159180
rect 9548 158722 9604 158732
rect 9436 157490 9492 157500
rect 9884 154420 9940 313628
rect 9884 154354 9940 154364
rect 9996 154308 10052 313740
rect 10444 313348 10500 313358
rect 10444 156212 10500 313292
rect 20188 301812 20244 320012
rect 20188 301746 20244 301756
rect 23548 301700 23604 320012
rect 26908 303492 26964 320012
rect 32284 317380 32340 320040
rect 32284 317314 32340 317324
rect 35308 320012 36120 320068
rect 26908 303426 26964 303436
rect 23548 301634 23604 301644
rect 35308 301588 35364 320012
rect 39900 317268 39956 320040
rect 39900 317202 39956 317212
rect 43708 317156 43764 320040
rect 43708 317090 43764 317100
rect 47068 320012 47544 320068
rect 50428 320012 51352 320068
rect 53788 320012 55160 320068
rect 47068 313796 47124 320012
rect 47068 313730 47124 313740
rect 50428 313684 50484 320012
rect 50428 313618 50484 313628
rect 53788 313572 53844 320012
rect 58940 317044 58996 320040
rect 58940 316978 58996 316988
rect 62748 316932 62804 320040
rect 62748 316866 62804 316876
rect 65548 320012 66584 320068
rect 68908 320012 70392 320068
rect 73948 320012 74200 320068
rect 77308 320012 78008 320068
rect 80668 320012 81816 320068
rect 53788 313506 53844 313516
rect 65548 313460 65604 320012
rect 65548 313394 65604 313404
rect 68908 313348 68964 320012
rect 68908 313282 68964 313292
rect 73948 310212 74004 320012
rect 73948 310146 74004 310156
rect 77308 310100 77364 320012
rect 77308 310034 77364 310044
rect 80668 303380 80724 320012
rect 85596 316820 85652 320040
rect 85596 316754 85652 316764
rect 89404 316708 89460 320040
rect 89404 316642 89460 316652
rect 92428 320012 93240 320068
rect 80668 303314 80724 303324
rect 92428 303268 92484 320012
rect 97020 316708 97076 320040
rect 97020 316642 97076 316652
rect 100828 306740 100884 320040
rect 104188 320012 104664 320068
rect 107548 320012 108472 320068
rect 104188 306852 104244 320012
rect 107548 306964 107604 320012
rect 112252 316820 112308 320040
rect 112252 316754 112308 316764
rect 115948 320012 116088 320068
rect 119308 320012 119896 320068
rect 122668 320012 123704 320068
rect 126028 320012 127512 320068
rect 115948 313348 116004 320012
rect 115948 313282 116004 313292
rect 119308 309988 119364 320012
rect 119308 309922 119364 309932
rect 122668 307076 122724 320012
rect 122668 307010 122724 307020
rect 107548 306898 107604 306908
rect 104188 306786 104244 306796
rect 100828 306674 100884 306684
rect 92428 303202 92484 303212
rect 126028 303268 126084 320012
rect 131292 316932 131348 320040
rect 131292 316866 131348 316876
rect 134428 320012 135128 320068
rect 137788 320012 138936 320068
rect 141148 320012 142744 320068
rect 134428 303380 134484 320012
rect 137788 303492 137844 320012
rect 141148 303604 141204 320012
rect 146524 317044 146580 320040
rect 150332 317156 150388 320040
rect 150332 317090 150388 317100
rect 152908 320012 154168 320068
rect 146524 316978 146580 316988
rect 152908 313460 152964 320012
rect 157948 313572 158004 320040
rect 161308 320012 161784 320068
rect 164668 320012 165592 320068
rect 168028 320012 169400 320068
rect 173068 320012 173208 320068
rect 161308 313684 161364 320012
rect 161308 313618 161364 313628
rect 157948 313506 158004 313516
rect 152908 313394 152964 313404
rect 164668 309988 164724 320012
rect 164668 309922 164724 309932
rect 168028 308308 168084 320012
rect 173068 311780 173124 320012
rect 176988 317268 177044 320040
rect 176988 317202 177044 317212
rect 179788 320012 180824 320068
rect 173068 311714 173124 311724
rect 168028 308242 168084 308252
rect 141148 303538 141204 303548
rect 137788 303426 137844 303436
rect 134428 303314 134484 303324
rect 126028 303202 126084 303212
rect 179788 302036 179844 320012
rect 184604 317380 184660 320040
rect 188972 319284 189028 587244
rect 188972 319218 189028 319228
rect 189868 587188 189924 587198
rect 184604 317314 184660 317324
rect 188300 317268 188356 317278
rect 188188 317156 188244 317166
rect 179788 301970 179844 301980
rect 188076 316820 188132 316830
rect 35308 301522 35364 301532
rect 188076 160244 188132 316764
rect 13244 157332 13300 160104
rect 17052 159684 17108 160104
rect 17052 159618 17108 159628
rect 20860 157780 20916 160104
rect 24668 157892 24724 160104
rect 20860 157714 20916 157724
rect 22652 157780 22708 157790
rect 13244 157266 13300 157276
rect 10444 156146 10500 156156
rect 9996 154242 10052 154252
rect 21868 145348 21924 145358
rect 21868 137788 21924 145292
rect 21868 137732 22148 137788
rect 11788 126084 11844 126094
rect 10892 116676 10948 116686
rect 9324 54786 9380 54796
rect 9996 74452 10052 74462
rect 9212 30146 9268 30156
rect 9996 21252 10052 74396
rect 10108 69076 10164 69086
rect 10108 62580 10164 69020
rect 10892 66948 10948 116620
rect 11676 77364 11732 77374
rect 10892 66882 10948 66892
rect 11564 70644 11620 70654
rect 10108 62514 10164 62524
rect 9996 21186 10052 21196
rect 10892 40628 10948 40638
rect 8316 21074 8372 21084
rect 7868 16482 7924 16492
rect 10892 16212 10948 40572
rect 11004 29764 11060 29774
rect 11004 20132 11060 29708
rect 11564 20244 11620 70588
rect 11564 20178 11620 20188
rect 11004 20066 11060 20076
rect 11676 19908 11732 77308
rect 11788 60564 11844 126028
rect 22092 115892 22148 137732
rect 22652 120148 22708 157724
rect 24668 156324 24724 157836
rect 28476 157556 28532 160104
rect 32284 159236 32340 160104
rect 32284 159170 32340 159180
rect 33292 159236 33348 159246
rect 28476 157220 28532 157500
rect 28476 157154 28532 157164
rect 31948 158900 32004 158910
rect 24668 156258 24724 156268
rect 27692 156324 27748 156334
rect 22652 120082 22708 120092
rect 26908 138628 26964 138638
rect 25564 119364 25620 119374
rect 24220 119252 24276 119262
rect 22092 115836 22904 115892
rect 24220 115864 24276 119196
rect 25564 115864 25620 119308
rect 26908 115864 26964 138572
rect 27692 135268 27748 156268
rect 27692 135202 27748 135212
rect 29372 143668 29428 143678
rect 27468 129444 27524 129454
rect 27468 115892 27524 129388
rect 28812 127764 28868 127774
rect 28812 115892 28868 127708
rect 29372 119252 29428 143612
rect 29372 119186 29428 119196
rect 30940 121044 30996 121054
rect 27468 115836 28280 115892
rect 28812 115836 29624 115892
rect 30940 115864 30996 120988
rect 31948 115892 32004 158844
rect 33292 156436 33348 159180
rect 33292 156370 33348 156380
rect 36092 157668 36148 160104
rect 36092 156324 36148 157612
rect 39900 159348 39956 160104
rect 39900 157108 39956 159292
rect 39900 157042 39956 157052
rect 41132 156436 41188 156446
rect 36092 156258 36148 156268
rect 37772 156324 37828 156334
rect 36988 133588 37044 133598
rect 34188 126084 34244 126094
rect 33628 121156 33684 121166
rect 31948 115836 32312 115892
rect 33628 115864 33684 121100
rect 34188 115892 34244 126028
rect 36876 116004 36932 116014
rect 36876 115892 36932 115948
rect 34188 115836 35000 115892
rect 36344 115836 36932 115892
rect 36988 115892 37044 133532
rect 37772 132692 37828 156268
rect 37772 132626 37828 132636
rect 41132 122612 41188 156380
rect 43708 154196 43764 160104
rect 46172 157220 46228 157230
rect 43708 154130 43764 154140
rect 44492 154196 44548 154206
rect 41132 122546 41188 122556
rect 43820 150388 43876 150398
rect 41692 119252 41748 119262
rect 40348 118468 40404 118478
rect 39004 118132 39060 118142
rect 36988 115836 37688 115892
rect 39004 115864 39060 118076
rect 40348 115864 40404 118412
rect 41692 115864 41748 119196
rect 43036 118692 43092 118702
rect 43036 115864 43092 118636
rect 43820 118132 43876 150332
rect 44492 129332 44548 154140
rect 44492 129266 44548 129276
rect 45388 148820 45444 148830
rect 43820 118066 43876 118076
rect 44380 123620 44436 123630
rect 44380 115864 44436 123564
rect 45388 119252 45444 148764
rect 46172 127652 46228 157164
rect 47516 154308 47572 160104
rect 51212 160076 51352 160132
rect 48748 155652 48804 155662
rect 47516 154242 47572 154252
rect 47852 154308 47908 154318
rect 46172 127586 46228 127596
rect 47068 137844 47124 137854
rect 47068 120708 47124 137788
rect 47852 136948 47908 154252
rect 47852 136882 47908 136892
rect 47068 120642 47124 120652
rect 47180 126980 47236 126990
rect 47180 120484 47236 126924
rect 45388 119186 45444 119196
rect 47068 120428 47236 120484
rect 47740 120708 47796 120718
rect 45724 118580 45780 118590
rect 45724 115864 45780 118524
rect 47068 115864 47124 120428
rect 47740 115892 47796 120652
rect 48748 118692 48804 155596
rect 51212 154420 51268 160076
rect 55132 159460 55188 160104
rect 58968 160076 59780 160132
rect 62776 160076 63140 160132
rect 55132 159394 55188 159404
rect 56364 159460 56420 159470
rect 55468 158788 55524 158798
rect 50428 140308 50484 140318
rect 48748 118626 48804 118636
rect 49756 119028 49812 119038
rect 47740 115836 48440 115892
rect 49756 115864 49812 118972
rect 50428 115892 50484 140252
rect 51212 124292 51268 154364
rect 51212 124226 51268 124236
rect 52892 155540 52948 155550
rect 52892 119028 52948 155484
rect 53788 150612 53844 150622
rect 53788 137788 53844 150556
rect 55468 137788 55524 158732
rect 56364 157220 56420 159404
rect 56364 157154 56420 157164
rect 59724 156996 59780 160076
rect 59612 143892 59668 143902
rect 53788 137732 54404 137788
rect 55468 137732 55748 137788
rect 52892 118962 52948 118972
rect 53788 118692 53844 118702
rect 52444 117684 52500 117694
rect 50428 115836 51128 115892
rect 52444 115864 52500 117628
rect 53788 115864 53844 118636
rect 54348 115892 54404 137732
rect 55692 115892 55748 137732
rect 57820 121828 57876 121838
rect 54348 115836 55160 115892
rect 55692 115836 56504 115892
rect 57820 115864 57876 121772
rect 59612 118692 59668 143836
rect 59724 131908 59780 156940
rect 62300 159012 62356 159022
rect 62300 137788 62356 158956
rect 63084 157444 63140 160076
rect 62972 152068 63028 152078
rect 62300 137732 62468 137788
rect 59724 131842 59780 131852
rect 59612 118626 59668 118636
rect 62412 115892 62468 137732
rect 62972 118580 63028 152012
rect 63084 128548 63140 157388
rect 66332 160076 66584 160132
rect 66332 154532 66388 160076
rect 63084 128482 63140 128492
rect 63868 148708 63924 148718
rect 62972 118514 63028 118524
rect 63868 115892 63924 148652
rect 65548 147028 65604 147038
rect 65548 118468 65604 146972
rect 66332 133700 66388 154476
rect 69692 156212 69748 156222
rect 68908 145460 68964 145470
rect 67228 141988 67284 141998
rect 67228 137788 67284 141932
rect 68908 137788 68964 145404
rect 67228 137732 67844 137788
rect 68908 137732 69188 137788
rect 66332 133634 66388 133644
rect 65548 118402 65604 118412
rect 67228 119252 67284 119262
rect 66556 116116 66612 116126
rect 66556 115892 66612 116060
rect 62412 115836 63224 115892
rect 63868 115836 64568 115892
rect 65912 115836 66612 115892
rect 67228 115864 67284 119196
rect 67788 115892 67844 137732
rect 69132 115892 69188 137732
rect 69692 131012 69748 156156
rect 70364 156212 70420 160104
rect 70364 156146 70420 156156
rect 71372 157108 71428 157118
rect 69692 130946 69748 130956
rect 70588 142100 70644 142110
rect 70588 115892 70644 142044
rect 71372 136052 71428 157052
rect 74172 156436 74228 160104
rect 77980 159572 78036 160104
rect 77980 159506 78036 159516
rect 78876 159572 78932 159582
rect 78876 157108 78932 159516
rect 78876 157042 78932 157052
rect 81788 159124 81844 160104
rect 74172 152852 74228 156380
rect 74172 152786 74228 152796
rect 78988 150500 79044 150510
rect 71372 135986 71428 135996
rect 73052 147028 73108 147038
rect 73052 119252 73108 146972
rect 75628 145572 75684 145582
rect 75628 137788 75684 145516
rect 77308 138740 77364 138750
rect 75628 137732 75908 137788
rect 73052 119186 73108 119196
rect 75852 115892 75908 137732
rect 77308 115892 77364 138684
rect 78988 115892 79044 150444
rect 81788 150388 81844 159068
rect 84812 160076 85624 160132
rect 89068 160076 89432 160132
rect 84812 156100 84868 160076
rect 81788 150322 81844 150332
rect 82348 155428 82404 155438
rect 82348 137788 82404 155372
rect 84028 153300 84084 153310
rect 82348 137732 82628 137788
rect 80668 118468 80724 118478
rect 67788 115836 68600 115892
rect 69132 115836 69944 115892
rect 70588 115836 71288 115892
rect 75852 115836 76664 115892
rect 77308 115836 78008 115892
rect 78988 115836 79352 115892
rect 80668 115864 80724 118412
rect 82012 116228 82068 116238
rect 82012 115864 82068 116172
rect 82572 115892 82628 137732
rect 84028 115892 84084 153244
rect 84812 147140 84868 156044
rect 84812 147074 84868 147084
rect 86492 157220 86548 157230
rect 85708 126196 85764 126206
rect 85708 115892 85764 126140
rect 86492 120372 86548 157164
rect 86716 157108 86772 157118
rect 86716 130228 86772 157052
rect 89068 149604 89124 160076
rect 93212 159236 93268 160104
rect 89068 148820 89124 149548
rect 89068 148754 89124 148764
rect 90636 157108 90692 157118
rect 87388 143780 87444 143790
rect 87388 137788 87444 143724
rect 87388 137732 88004 137788
rect 86716 130162 86772 130172
rect 86492 120306 86548 120316
rect 87388 118356 87444 118366
rect 82572 115836 83384 115892
rect 84028 115836 84728 115892
rect 85708 115836 86072 115892
rect 87388 115864 87444 118300
rect 87948 115892 88004 137732
rect 89068 125972 89124 125982
rect 89068 123620 89124 125916
rect 90636 125972 90692 157052
rect 90636 125906 90692 125916
rect 91532 156324 91588 156334
rect 89068 123554 89124 123564
rect 90076 125300 90132 125310
rect 89180 123508 89236 123518
rect 89180 118356 89236 123452
rect 89180 118290 89236 118300
rect 87948 115836 88760 115892
rect 90076 115864 90132 125244
rect 91420 125188 91476 125198
rect 91420 115864 91476 125132
rect 91532 123620 91588 156268
rect 93212 155652 93268 159180
rect 97020 157108 97076 160104
rect 100856 160076 100996 160132
rect 97020 157042 97076 157052
rect 97468 160020 97524 160030
rect 93212 155586 93268 155596
rect 96012 131124 96068 131134
rect 91532 123554 91588 123564
rect 94108 126868 94164 126878
rect 92764 120260 92820 120270
rect 92764 115864 92820 120204
rect 94108 115864 94164 126812
rect 95452 117908 95508 117918
rect 95452 115864 95508 117852
rect 96012 115892 96068 131068
rect 97468 115892 97524 159964
rect 100940 154532 100996 160076
rect 99148 153748 99204 153758
rect 99148 115892 99204 153692
rect 100828 152292 100884 152302
rect 100828 120708 100884 152236
rect 100940 152068 100996 154476
rect 100940 152002 100996 152012
rect 104188 160076 104664 160132
rect 107660 160076 108472 160132
rect 100828 120642 100884 120652
rect 101052 131236 101108 131246
rect 96012 115836 96824 115892
rect 97468 115836 98168 115892
rect 99148 115836 99512 115892
rect 101052 115780 101108 131180
rect 104188 129220 104244 160076
rect 107436 153860 107492 153870
rect 107324 139412 107380 139422
rect 104188 129154 104244 129164
rect 104972 139076 105028 139086
rect 104860 122724 104916 122734
rect 101500 120708 101556 120718
rect 101500 115892 101556 120652
rect 103516 119252 103572 119262
rect 101500 115836 102200 115892
rect 103516 115864 103572 119196
rect 104860 115864 104916 122668
rect 104972 119252 105028 139020
rect 107324 137844 107380 139356
rect 105532 129220 105588 129230
rect 105532 126980 105588 129164
rect 105532 126914 105588 126924
rect 107324 121940 107380 137788
rect 107436 124180 107492 153804
rect 107436 122724 107492 124124
rect 107436 122658 107492 122668
rect 107548 147140 107604 147150
rect 107324 121874 107380 121884
rect 104972 119186 105028 119196
rect 106204 119140 106260 119150
rect 106204 115864 106260 119084
rect 107548 115864 107604 147084
rect 107660 139412 107716 160076
rect 112252 159572 112308 160104
rect 116088 160076 116788 160132
rect 112252 155540 112308 159516
rect 116732 156996 116788 160076
rect 112252 155474 112308 155484
rect 114268 155540 114324 155550
rect 110012 153972 110068 153982
rect 107660 139346 107716 139356
rect 109228 148148 109284 148158
rect 107660 138964 107716 138974
rect 107660 137788 107716 138908
rect 109228 137788 109284 148092
rect 107660 137732 108164 137788
rect 109228 137732 109508 137788
rect 108108 115892 108164 137732
rect 109452 115892 109508 137732
rect 110012 119140 110068 153916
rect 110012 119074 110068 119084
rect 110908 152068 110964 152078
rect 110908 115892 110964 152012
rect 112588 142212 112644 142222
rect 112588 115892 112644 142156
rect 108108 115836 108920 115892
rect 109452 115836 110264 115892
rect 110908 115836 111608 115892
rect 112588 115836 112952 115892
rect 114268 115864 114324 155484
rect 116732 140308 116788 156940
rect 119420 160076 119896 160132
rect 122892 160104 123704 160132
rect 122892 160076 123732 160104
rect 116732 140242 116788 140252
rect 117628 155652 117684 155662
rect 116956 119476 117012 119486
rect 115612 117796 115668 117806
rect 115612 115864 115668 117740
rect 116956 115864 117012 119420
rect 117628 115892 117684 155596
rect 119308 152180 119364 152190
rect 119308 115892 119364 152124
rect 119420 143892 119476 160076
rect 122892 149548 122948 160076
rect 123676 159796 123732 160076
rect 123676 159730 123732 159740
rect 127484 153860 127540 160104
rect 131292 154420 131348 160104
rect 131292 153972 131348 154364
rect 131292 153906 131348 153916
rect 134428 160076 135128 160132
rect 137788 160076 138936 160132
rect 141148 160076 142744 160132
rect 146188 160076 146552 160132
rect 149548 160076 150360 160132
rect 153692 160076 154168 160132
rect 157976 160076 158788 160132
rect 161784 160076 162148 160132
rect 127484 153794 127540 153804
rect 127708 153860 127764 153870
rect 119420 143826 119476 143836
rect 122668 149492 122948 149548
rect 126028 152404 126084 152414
rect 122668 139076 122724 149492
rect 122668 139010 122724 139020
rect 122668 138852 122724 138862
rect 122668 137788 122724 138796
rect 122668 137732 122948 137788
rect 120988 126308 121044 126318
rect 117628 115836 118328 115892
rect 119308 115836 119672 115892
rect 120988 115864 121044 126252
rect 122332 124404 122388 124414
rect 122332 115864 122388 124348
rect 122892 115892 122948 137732
rect 125020 122724 125076 122734
rect 122892 115836 123704 115892
rect 125020 115864 125076 122668
rect 126028 115892 126084 152348
rect 127708 137788 127764 153804
rect 134428 149492 134484 160076
rect 134428 147140 134484 149436
rect 136892 148036 136948 148046
rect 134428 147074 134484 147084
rect 135212 147924 135268 147934
rect 127708 137732 128324 137788
rect 127708 118020 127764 118030
rect 126028 115836 126392 115892
rect 127708 115864 127764 117964
rect 128268 115892 128324 137732
rect 131068 137060 131124 137070
rect 130396 116340 130452 116350
rect 128268 115836 129080 115892
rect 130396 115864 130452 116284
rect 131068 115892 131124 137004
rect 135212 127652 135268 147868
rect 135212 126028 135268 127596
rect 134988 125972 135268 126028
rect 135324 135268 135380 135278
rect 133084 120148 133140 120158
rect 133084 119140 133140 120092
rect 131068 115836 131768 115892
rect 133084 115864 133140 119084
rect 134428 119252 134484 119262
rect 134428 115864 134484 119196
rect 134988 115892 135044 125972
rect 135324 119252 135380 135212
rect 135324 119186 135380 119196
rect 136892 119140 136948 147980
rect 137004 146244 137060 146254
rect 137004 137788 137060 146188
rect 137788 139412 137844 160076
rect 140252 149716 140308 149726
rect 137788 139346 137844 139356
rect 138572 142884 138628 142894
rect 137004 137732 137172 137788
rect 136892 119074 136948 119084
rect 137116 122612 137172 137732
rect 134988 115836 135800 115892
rect 137116 115864 137172 122556
rect 137788 132692 137844 132702
rect 137788 115892 137844 132636
rect 138572 132692 138628 142828
rect 138572 132626 138628 132636
rect 139468 136052 139524 136062
rect 139468 115892 139524 135996
rect 140252 136052 140308 149660
rect 141148 149548 141204 160076
rect 141036 149492 141204 149548
rect 141036 148148 141092 149492
rect 141036 137732 141092 148092
rect 146188 147812 146244 160076
rect 146188 147746 146244 147756
rect 149548 147028 149604 160076
rect 149548 146962 149604 146972
rect 153692 157668 153748 160076
rect 148652 146468 148708 146478
rect 141036 137666 141092 137676
rect 142044 146356 142100 146366
rect 140252 135986 140308 135996
rect 141932 136948 141988 136958
rect 141932 136500 141988 136892
rect 141148 129332 141204 129342
rect 137788 115836 138488 115892
rect 139468 115836 139832 115892
rect 141148 115864 141204 129276
rect 141932 115892 141988 136444
rect 142044 129332 142100 146300
rect 143724 144564 143780 144574
rect 143612 142996 143668 143006
rect 143612 136500 143668 142940
rect 143724 137788 143780 144508
rect 143724 137732 143892 137788
rect 143612 136434 143668 136444
rect 142044 129266 142100 129276
rect 143836 124292 143892 137732
rect 141932 115836 142520 115892
rect 143836 115864 143892 124236
rect 145292 131908 145348 131918
rect 145292 122836 145348 131852
rect 147868 128548 147924 128558
rect 145292 122770 145348 122780
rect 146524 122836 146580 122846
rect 145180 120372 145236 120382
rect 145180 119588 145236 120316
rect 145180 115864 145236 119532
rect 146524 115864 146580 122780
rect 147868 121268 147924 128492
rect 147868 115864 147924 121212
rect 148652 119252 148708 146412
rect 150332 144676 150388 144686
rect 148652 119186 148708 119196
rect 148876 133700 148932 133710
rect 148876 119252 148932 133644
rect 148876 115892 148932 119196
rect 149772 131012 149828 131022
rect 149772 115892 149828 130956
rect 150332 131012 150388 144620
rect 150332 130946 150388 130956
rect 151900 123620 151956 123630
rect 151900 119700 151956 123564
rect 153692 123508 153748 157612
rect 158732 156884 158788 160076
rect 156268 150388 156324 150398
rect 156268 137788 156324 150332
rect 157948 148820 158004 148830
rect 156268 137732 156548 137788
rect 153692 123442 153748 123452
rect 153804 130228 153860 130238
rect 153804 124516 153860 130172
rect 148876 115836 149240 115892
rect 149772 115836 150584 115892
rect 151900 115864 151956 119644
rect 153804 115892 153860 124460
rect 155932 123508 155988 123518
rect 153272 115836 153860 115892
rect 154588 118132 154644 118142
rect 154588 115864 154644 118076
rect 155932 115864 155988 123452
rect 156492 115892 156548 137732
rect 157948 115892 158004 148764
rect 158732 143780 158788 156828
rect 162092 157556 162148 160076
rect 158732 143714 158788 143724
rect 160412 152516 160468 152526
rect 159628 140308 159684 140318
rect 159628 115892 159684 140252
rect 160412 119252 160468 152460
rect 162092 125300 162148 157500
rect 165564 157444 165620 160104
rect 162092 125234 162148 125244
rect 163772 156324 163828 156334
rect 163772 125188 163828 156268
rect 165564 156324 165620 157388
rect 165564 156258 165620 156268
rect 166348 158788 166404 158798
rect 163772 125122 163828 125132
rect 160412 119186 160468 119196
rect 165340 118580 165396 118590
rect 156492 115836 157304 115892
rect 157948 115836 158648 115892
rect 159628 115836 159992 115892
rect 165340 115864 165396 118524
rect 166348 115892 166404 158732
rect 169372 157892 169428 160104
rect 173208 160076 173908 160132
rect 167132 156324 167188 156334
rect 167132 120260 167188 156268
rect 169372 156324 169428 157836
rect 169372 156258 169428 156268
rect 173852 157332 173908 160076
rect 168028 153972 168084 153982
rect 168028 137788 168084 153916
rect 169708 148932 169764 148942
rect 169708 137788 169764 148876
rect 168028 137732 168644 137788
rect 169708 137732 169988 137788
rect 167132 120194 167188 120204
rect 168028 116452 168084 116462
rect 166348 115836 166712 115892
rect 168028 115864 168084 116396
rect 168588 115892 168644 137732
rect 169932 115892 169988 137732
rect 171388 128548 171444 128558
rect 171388 115892 171444 128492
rect 173852 126868 173908 157276
rect 173852 126802 173908 126812
rect 175532 156324 175588 156334
rect 175532 123508 175588 156268
rect 176988 156324 177044 160104
rect 176988 156258 177044 156268
rect 180572 160076 180824 160132
rect 180572 157220 180628 160076
rect 180572 143668 180628 157164
rect 184604 153972 184660 160104
rect 188076 159572 188132 160188
rect 188076 159506 188132 159516
rect 184604 153906 184660 153916
rect 188188 145460 188244 317100
rect 188300 148820 188356 317212
rect 188972 317044 189028 317054
rect 188748 311780 188804 311790
rect 188300 148754 188356 148764
rect 188412 303604 188468 303614
rect 188412 302596 188468 303548
rect 188188 145394 188244 145404
rect 180572 143602 180628 143612
rect 188412 137732 188468 302540
rect 188524 303492 188580 303502
rect 188524 302484 188580 303436
rect 188524 139412 188580 302428
rect 188636 303380 188692 303390
rect 188636 149492 188692 303324
rect 188748 157332 188804 311724
rect 188860 308420 188916 308430
rect 188860 157892 188916 308364
rect 188860 157826 188916 157836
rect 188748 157266 188804 157276
rect 188972 157780 189028 316988
rect 188636 149426 188692 149436
rect 188972 147812 189028 157724
rect 189644 316932 189700 316942
rect 189644 161364 189700 316876
rect 189644 154420 189700 161308
rect 189644 154354 189700 154364
rect 188972 147746 189028 147756
rect 188524 139346 188580 139356
rect 188412 137666 188468 137676
rect 175532 123442 175588 123452
rect 188972 129444 189028 129454
rect 178780 118804 178836 118814
rect 173404 118692 173460 118702
rect 168588 115836 169400 115892
rect 169932 115836 170744 115892
rect 171388 115836 172088 115892
rect 173404 115864 173460 118636
rect 176876 117908 176932 117918
rect 176876 116788 176932 117852
rect 176876 116722 176932 116732
rect 178780 115864 178836 118748
rect 100856 115724 101108 115780
rect 180152 115388 180516 115444
rect 19292 113092 19348 113102
rect 19180 88900 19236 88910
rect 18172 71428 18228 71438
rect 18172 70644 18228 71372
rect 18172 70578 18228 70588
rect 19180 69972 19236 88844
rect 19292 70756 19348 113036
rect 20076 111748 20132 111758
rect 19964 110404 20020 110414
rect 19852 109060 19908 109070
rect 19516 99652 19572 99662
rect 19292 70690 19348 70700
rect 19404 94164 19460 94174
rect 19180 69906 19236 69916
rect 19404 69188 19460 94108
rect 19516 70980 19572 99596
rect 19740 98308 19796 98318
rect 19628 96964 19684 96974
rect 19628 73668 19684 96908
rect 19628 73602 19684 73612
rect 19516 70914 19572 70924
rect 19740 69748 19796 98252
rect 19852 72548 19908 109004
rect 19964 73556 20020 110348
rect 19964 73490 20020 73500
rect 20076 73444 20132 111692
rect 20076 73378 20132 73388
rect 20188 106372 20244 106382
rect 19852 72482 19908 72492
rect 20188 70196 20244 106316
rect 20412 105028 20468 105038
rect 20188 70130 20244 70140
rect 20300 103684 20356 103694
rect 19740 69682 19796 69692
rect 19404 69122 19460 69132
rect 20300 68628 20356 103628
rect 20412 70084 20468 104972
rect 20412 70018 20468 70028
rect 21868 72324 21924 72334
rect 21868 69412 21924 72268
rect 47404 70756 47460 70766
rect 47404 70690 47460 70700
rect 21868 69346 21924 69356
rect 21980 70532 22036 70542
rect 21980 68852 22036 70476
rect 64092 70196 64148 70206
rect 21980 68786 22036 68796
rect 25564 70028 26264 70084
rect 20300 68562 20356 68572
rect 25564 68404 25620 70028
rect 25564 68338 25620 68348
rect 28588 68404 28644 70056
rect 30940 69188 30996 70056
rect 33292 69412 33348 70056
rect 33292 69346 33348 69356
rect 30940 69122 30996 69132
rect 31164 69188 31220 69198
rect 31164 68852 31220 69132
rect 35644 69076 35700 70056
rect 35644 69010 35700 69020
rect 37324 70028 38024 70084
rect 31164 68786 31220 68796
rect 37324 68628 37380 70028
rect 40348 69188 40404 70056
rect 40348 69122 40404 69132
rect 42028 70028 42728 70084
rect 37324 68562 37380 68572
rect 42028 68628 42084 70028
rect 45052 68964 45108 70056
rect 45052 68898 45108 68908
rect 49084 70028 49784 70084
rect 42028 68562 42084 68572
rect 49084 68628 49140 70028
rect 49084 68562 49140 68572
rect 52108 68628 52164 70056
rect 52108 68562 52164 68572
rect 53788 70028 54488 70084
rect 56140 70028 56840 70084
rect 58828 70028 59192 70084
rect 60844 70028 61544 70084
rect 53788 68628 53844 70028
rect 53788 68562 53844 68572
rect 56140 68628 56196 70028
rect 56140 68562 56196 68572
rect 58828 68516 58884 70028
rect 58828 68450 58884 68460
rect 60844 68516 60900 70028
rect 60844 68450 60900 68460
rect 28588 68338 28644 68348
rect 63868 67172 63924 70056
rect 63868 67106 63924 67116
rect 63980 69748 64036 69758
rect 61516 66164 61572 66174
rect 11788 60498 11844 60508
rect 60508 66108 61516 66164
rect 60508 35308 60564 66108
rect 61516 66098 61572 66108
rect 61516 64708 61572 64718
rect 61516 55468 61572 64652
rect 60284 35252 60564 35308
rect 60620 55412 61572 55468
rect 60284 23604 60340 35252
rect 60620 27412 60676 55412
rect 63980 50820 64036 69692
rect 64092 59556 64148 70140
rect 64540 70084 64596 70094
rect 64428 70028 64540 70084
rect 64092 59490 64148 59500
rect 64204 69860 64260 69870
rect 63980 50754 64036 50764
rect 61516 44324 61572 44334
rect 61516 43708 61572 44268
rect 60844 43652 61572 43708
rect 60844 38668 60900 43652
rect 64204 43540 64260 69804
rect 64316 68628 64372 68638
rect 64316 56644 64372 68572
rect 64428 58100 64484 70028
rect 64540 70018 64596 70028
rect 64876 69972 64932 69982
rect 64764 63924 64820 63934
rect 64428 58034 64484 58044
rect 64652 62468 64708 62478
rect 64316 56578 64372 56588
rect 64204 43474 64260 43484
rect 64316 52276 64372 52286
rect 63868 42084 63924 42094
rect 60732 38612 60900 38668
rect 62188 39172 62244 39182
rect 60732 29426 60788 38612
rect 61516 37044 61572 37054
rect 60732 29374 60734 29426
rect 60786 29374 60788 29426
rect 60732 29362 60788 29374
rect 60956 36988 61516 37044
rect 60620 27356 60900 27412
rect 60732 27188 60788 27198
rect 60396 27186 60788 27188
rect 60396 27134 60734 27186
rect 60786 27134 60788 27186
rect 60396 27132 60788 27134
rect 60396 23716 60452 27132
rect 60732 27122 60788 27132
rect 60844 26068 60900 27356
rect 60620 26012 60900 26068
rect 60396 23660 60564 23716
rect 60284 23548 60452 23604
rect 11676 19842 11732 19852
rect 14924 18564 14980 20104
rect 14924 18498 14980 18508
rect 20412 17556 20468 20104
rect 25228 20076 25928 20132
rect 30268 20076 31416 20132
rect 35308 20076 36904 20132
rect 20412 17490 20468 17500
rect 23436 17556 23492 17566
rect 10892 16146 10948 16156
rect 23436 15092 23492 17500
rect 23436 15026 23492 15036
rect 4508 8306 4564 8316
rect 4284 8194 4340 8204
rect 25228 4228 25284 20076
rect 30268 5908 30324 20076
rect 30268 5842 30324 5852
rect 35308 4340 35364 20076
rect 42364 16884 42420 20104
rect 42364 16818 42420 16828
rect 44716 16884 44772 16894
rect 44716 13412 44772 16828
rect 44716 13346 44772 13356
rect 47852 10948 47908 20104
rect 53340 17668 53396 20104
rect 53340 17602 53396 17612
rect 58828 12628 58884 20104
rect 60396 12964 60452 23548
rect 60508 14644 60564 23660
rect 60620 19572 60676 26012
rect 60620 19506 60676 19516
rect 60732 23714 60788 23726
rect 60732 23662 60734 23714
rect 60786 23662 60788 23714
rect 60732 14868 60788 23662
rect 60956 23548 61012 36988
rect 61516 36978 61572 36988
rect 61068 29426 61124 29438
rect 61068 29374 61070 29426
rect 61122 29374 61124 29426
rect 61068 23714 61124 29374
rect 61964 27188 62020 27198
rect 61964 27094 62020 27132
rect 61068 23662 61070 23714
rect 61122 23662 61124 23714
rect 61068 23650 61124 23662
rect 60844 23492 61012 23548
rect 60844 21028 60900 23492
rect 60844 20962 60900 20972
rect 61516 22484 61572 22494
rect 61516 20020 61572 22428
rect 61516 19954 61572 19964
rect 60732 14802 60788 14812
rect 60508 14578 60564 14588
rect 60396 12898 60452 12908
rect 58828 12562 58884 12572
rect 47852 10882 47908 10892
rect 62188 10052 62244 39116
rect 62300 31892 62356 31902
rect 62300 16324 62356 31836
rect 63868 16436 63924 42028
rect 63980 26068 64036 26078
rect 63980 21252 64036 26012
rect 63980 21186 64036 21196
rect 63868 16370 63924 16380
rect 62300 16258 62356 16268
rect 64316 13300 64372 52220
rect 64540 49364 64596 49374
rect 64428 47908 64484 47918
rect 64428 16660 64484 47852
rect 64540 18228 64596 49308
rect 64540 18162 64596 18172
rect 64428 16594 64484 16604
rect 64316 13234 64372 13244
rect 64652 13076 64708 62412
rect 64764 14532 64820 63868
rect 64876 40628 64932 69916
rect 66220 68964 66276 70056
rect 66220 68898 66276 68908
rect 68572 68852 68628 70056
rect 68572 68786 68628 68796
rect 70924 65492 70980 70056
rect 73276 67060 73332 70056
rect 75628 69076 75684 70056
rect 77980 69188 78036 70056
rect 77980 69122 78036 69132
rect 75628 69010 75684 69020
rect 80332 68740 80388 70056
rect 80332 68674 80388 68684
rect 73276 66994 73332 67004
rect 70924 65426 70980 65436
rect 82684 63812 82740 70056
rect 85036 66836 85092 70056
rect 87388 66948 87444 70056
rect 89740 68628 89796 70056
rect 89740 68562 89796 68572
rect 90748 70028 92120 70084
rect 94108 70028 94472 70084
rect 87388 66882 87444 66892
rect 85036 66770 85092 66780
rect 82684 63746 82740 63756
rect 65100 61012 65156 61022
rect 64876 40562 64932 40572
rect 64988 55188 65044 55198
rect 64988 14980 65044 55132
rect 64988 14914 65044 14924
rect 64764 14466 64820 14476
rect 65100 13188 65156 60956
rect 90748 14420 90804 70028
rect 90748 14354 90804 14364
rect 65100 13122 65156 13132
rect 64652 13010 64708 13020
rect 62188 9986 62244 9996
rect 94108 6132 94164 70028
rect 96796 65604 96852 70056
rect 96796 65538 96852 65548
rect 98252 65604 98308 65614
rect 94108 6066 94164 6076
rect 98252 4564 98308 65548
rect 99148 21140 99204 70056
rect 100828 70028 101528 70084
rect 102508 70028 103880 70084
rect 105868 70028 106232 70084
rect 107548 70028 108584 70084
rect 100828 24388 100884 70028
rect 100828 24322 100884 24332
rect 102508 22708 102564 70028
rect 102508 22642 102564 22652
rect 99148 21074 99204 21084
rect 105868 7700 105924 70028
rect 107548 27748 107604 70028
rect 110908 65604 110964 70056
rect 110908 65538 110964 65548
rect 113260 63028 113316 70056
rect 113260 62962 113316 62972
rect 113372 65604 113428 65614
rect 107548 27682 107604 27692
rect 105868 7634 105924 7644
rect 98252 4498 98308 4508
rect 113372 4452 113428 65548
rect 115612 65604 115668 70056
rect 117628 70028 117992 70084
rect 119308 70028 120344 70084
rect 115612 65538 115668 65548
rect 116732 65604 116788 65614
rect 116732 9380 116788 65548
rect 116732 9314 116788 9324
rect 117628 7588 117684 70028
rect 119308 21028 119364 70028
rect 119308 20962 119364 20972
rect 117628 7522 117684 7532
rect 122668 6020 122724 70056
rect 124348 70028 125048 70084
rect 126028 70028 127400 70084
rect 124348 11060 124404 70028
rect 124348 10994 124404 11004
rect 126028 9268 126084 70028
rect 129724 61348 129780 70056
rect 129724 61282 129780 61292
rect 131068 70028 132104 70084
rect 131068 15092 131124 70028
rect 131068 15026 131124 15036
rect 131628 15092 131684 15102
rect 131628 14308 131684 15036
rect 131628 14242 131684 14252
rect 126028 9202 126084 9212
rect 134428 7924 134484 70056
rect 136108 70028 136808 70084
rect 137788 70028 139160 70084
rect 141148 70028 141512 70084
rect 142828 70028 143864 70084
rect 136108 8036 136164 70028
rect 136108 7970 136164 7980
rect 134428 7858 134484 7868
rect 122668 5954 122724 5964
rect 134428 7700 134484 7710
rect 134428 4676 134484 7644
rect 137788 7476 137844 70028
rect 140028 14420 140084 14430
rect 137788 7410 137844 7420
rect 138460 7924 138516 7934
rect 134428 4610 134484 4620
rect 113372 4386 113428 4396
rect 35308 4274 35364 4284
rect 25228 4162 25284 4172
rect 138460 480 138516 7868
rect 19768 -960 19992 480
rect 20888 -960 21112 480
rect 22008 -960 22232 480
rect 23128 -960 23352 480
rect 24248 -960 24472 480
rect 25368 -960 25592 480
rect 26488 -960 26712 480
rect 27608 -960 27832 480
rect 28728 -960 28952 480
rect 29848 -960 30072 480
rect 30968 -960 31192 480
rect 32088 -960 32312 480
rect 33208 -960 33432 480
rect 34328 -960 34552 480
rect 35448 -960 35672 480
rect 36568 -960 36792 480
rect 37688 -960 37912 480
rect 38808 -960 39032 480
rect 39928 -960 40152 480
rect 41048 -960 41272 480
rect 42168 -960 42392 480
rect 43288 -960 43512 480
rect 44408 -960 44632 480
rect 45528 -960 45752 480
rect 46648 -960 46872 480
rect 47768 -960 47992 480
rect 48888 -960 49112 480
rect 50008 -960 50232 480
rect 51128 -960 51352 480
rect 52248 -960 52472 480
rect 53368 -960 53592 480
rect 54488 -960 54712 480
rect 55608 -960 55832 480
rect 56728 -960 56952 480
rect 57848 -960 58072 480
rect 58968 -960 59192 480
rect 60088 -960 60312 480
rect 61208 -960 61432 480
rect 62328 -960 62552 480
rect 63448 -960 63672 480
rect 64568 -960 64792 480
rect 65688 -960 65912 480
rect 66808 -960 67032 480
rect 67928 -960 68152 480
rect 69048 -960 69272 480
rect 70168 -960 70392 480
rect 71288 -960 71512 480
rect 72408 -960 72632 480
rect 73528 -960 73752 480
rect 74648 -960 74872 480
rect 75768 -960 75992 480
rect 76888 -960 77112 480
rect 78008 -960 78232 480
rect 79128 -960 79352 480
rect 80248 -960 80472 480
rect 81368 -960 81592 480
rect 82488 -960 82712 480
rect 83608 -960 83832 480
rect 84728 -960 84952 480
rect 85848 -960 86072 480
rect 86968 -960 87192 480
rect 88088 -960 88312 480
rect 89208 -960 89432 480
rect 90328 -960 90552 480
rect 91448 -960 91672 480
rect 92568 -960 92792 480
rect 93688 -960 93912 480
rect 94808 -960 95032 480
rect 95928 -960 96152 480
rect 97048 -960 97272 480
rect 98168 -960 98392 480
rect 99288 -960 99512 480
rect 100408 -960 100632 480
rect 101528 -960 101752 480
rect 102648 -960 102872 480
rect 103768 -960 103992 480
rect 104888 -960 105112 480
rect 106008 -960 106232 480
rect 107128 -960 107352 480
rect 108248 -960 108472 480
rect 109368 -960 109592 480
rect 110488 -960 110712 480
rect 111608 -960 111832 480
rect 112728 -960 112952 480
rect 113848 -960 114072 480
rect 114968 -960 115192 480
rect 116088 -960 116312 480
rect 117208 -960 117432 480
rect 118328 -960 118552 480
rect 119448 -960 119672 480
rect 120568 -960 120792 480
rect 121688 -960 121912 480
rect 122808 -960 123032 480
rect 123928 -960 124152 480
rect 125048 -960 125272 480
rect 126168 -960 126392 480
rect 127288 -960 127512 480
rect 128408 -960 128632 480
rect 129528 -960 129752 480
rect 130648 -960 130872 480
rect 131768 -960 131992 480
rect 132888 -960 133112 480
rect 134008 -960 134232 480
rect 135128 -960 135352 480
rect 136248 -960 136472 480
rect 137368 -960 137592 480
rect 138460 392 138712 480
rect 138488 -960 138712 392
rect 139608 -960 139832 480
rect 140028 420 140084 14364
rect 141148 6804 141204 70028
rect 142828 8484 142884 70028
rect 146188 65940 146244 70056
rect 146188 65874 146244 65884
rect 147868 70028 148568 70084
rect 149548 70028 150920 70084
rect 152908 70028 153272 70084
rect 147868 22932 147924 70028
rect 147980 65940 148036 65950
rect 147980 64708 148036 65884
rect 147980 64642 148036 64652
rect 147868 22866 147924 22876
rect 142828 8418 142884 8428
rect 145292 22708 145348 22718
rect 141148 6738 141204 6748
rect 141820 8036 141876 8046
rect 140588 480 140756 532
rect 141820 480 141876 7980
rect 145180 7476 145236 7486
rect 144060 6132 144116 6142
rect 144060 480 144116 6076
rect 145180 480 145236 7420
rect 145292 4788 145348 22652
rect 148652 21140 148708 21150
rect 145292 4722 145348 4732
rect 148540 6804 148596 6814
rect 147420 4564 147476 4574
rect 147420 480 147476 4508
rect 148540 480 148596 6748
rect 148652 5012 148708 21084
rect 149548 14644 149604 70028
rect 152908 26852 152964 70028
rect 152908 26786 152964 26796
rect 154588 64708 154644 64718
rect 152908 24388 152964 24398
rect 152908 20188 152964 24332
rect 152908 20132 153524 20188
rect 149548 14578 149604 14588
rect 151900 8484 151956 8494
rect 148652 4946 148708 4956
rect 150780 5012 150836 5022
rect 150780 480 150836 4956
rect 151900 480 151956 8428
rect 140588 476 140952 480
rect 140588 420 140644 476
rect 140028 364 140644 420
rect 140700 392 140952 476
rect 141820 392 142072 480
rect 140728 -960 140952 392
rect 141848 -960 142072 392
rect 142968 -960 143192 480
rect 144060 392 144312 480
rect 145180 392 145432 480
rect 144088 -960 144312 392
rect 145208 -960 145432 392
rect 146328 -960 146552 480
rect 147420 392 147672 480
rect 148540 392 148792 480
rect 147448 -960 147672 392
rect 148568 -960 148792 392
rect 149688 -960 149912 480
rect 150780 392 151032 480
rect 151900 392 152152 480
rect 150808 -960 151032 392
rect 151928 -960 152152 392
rect 153048 -960 153272 480
rect 153468 420 153524 20132
rect 154028 480 154196 532
rect 154028 476 154392 480
rect 154028 420 154084 476
rect 153468 364 154084 420
rect 154140 392 154392 476
rect 154168 -960 154392 392
rect 154588 420 154644 64652
rect 155596 64708 155652 70056
rect 155596 64642 155652 64652
rect 157052 27748 157108 27758
rect 157052 4900 157108 27692
rect 157948 22708 158004 70056
rect 159628 70028 160328 70084
rect 157948 22642 158004 22652
rect 158060 22932 158116 22942
rect 157052 4834 157108 4844
rect 157500 4788 157556 4798
rect 155148 480 155316 532
rect 157500 480 157556 4732
rect 155148 476 155512 480
rect 155148 420 155204 476
rect 154588 364 155204 420
rect 155260 392 155512 476
rect 155288 -960 155512 392
rect 156408 -960 156632 480
rect 157500 392 157752 480
rect 157528 -960 157752 392
rect 158060 420 158116 22876
rect 159628 12852 159684 70028
rect 162652 65604 162708 70056
rect 162652 65538 162708 65548
rect 163772 65604 163828 65614
rect 162092 63028 162148 63038
rect 159628 12786 159684 12796
rect 160412 14644 160468 14654
rect 160412 5012 160468 14588
rect 160412 4946 160468 4956
rect 161980 5012 162036 5022
rect 160860 4676 160916 4686
rect 158508 480 158676 532
rect 160860 480 160916 4620
rect 161980 480 162036 4956
rect 162092 4788 162148 62972
rect 163772 26068 163828 65548
rect 165004 64820 165060 70056
rect 165004 64754 165060 64764
rect 166348 70028 167384 70084
rect 163772 26002 163828 26012
rect 163996 26852 164052 26862
rect 162092 4722 162148 4732
rect 163996 4452 164052 26796
rect 166348 7700 166404 70028
rect 169708 11172 169764 70056
rect 171500 64708 171556 64718
rect 169708 11106 169764 11116
rect 171388 22708 171444 22718
rect 166348 7634 166404 7644
rect 170268 11060 170324 11070
rect 163996 4386 164052 4396
rect 164220 4900 164276 4910
rect 164220 480 164276 4844
rect 167580 4564 167636 4574
rect 165340 4452 165396 4462
rect 165340 480 165396 4396
rect 167580 480 167636 4508
rect 170268 4452 170324 11004
rect 170268 4386 170324 4396
rect 170940 4788 170996 4798
rect 168924 4116 168980 4126
rect 168924 480 168980 4060
rect 170940 480 170996 4732
rect 158508 476 158872 480
rect 158508 420 158564 476
rect 158060 364 158564 420
rect 158620 392 158872 476
rect 158648 -960 158872 392
rect 159768 -960 159992 480
rect 160860 392 161112 480
rect 161980 392 162232 480
rect 160888 -960 161112 392
rect 162008 -960 162232 392
rect 163128 -960 163352 480
rect 164220 392 164472 480
rect 165340 392 165592 480
rect 164248 -960 164472 392
rect 165368 -960 165592 392
rect 166488 -960 166712 480
rect 167580 392 167832 480
rect 167608 -960 167832 392
rect 168728 392 168980 480
rect 168728 -960 168952 392
rect 169848 -960 170072 480
rect 170940 392 171192 480
rect 170968 -960 171192 392
rect 171388 420 171444 22652
rect 171500 4116 171556 64652
rect 172060 63028 172116 70056
rect 172060 62962 172116 62972
rect 173068 70028 174440 70084
rect 173068 13412 173124 70028
rect 176764 55468 176820 70056
rect 175532 55412 177268 55468
rect 175532 18564 175588 55412
rect 175532 18498 175588 18508
rect 173068 13346 173124 13356
rect 174636 13412 174692 13422
rect 174636 12740 174692 13356
rect 174636 12674 174692 12684
rect 174748 12852 174804 12862
rect 171500 4050 171556 4060
rect 174300 9380 174356 9390
rect 171948 480 172116 532
rect 174300 480 174356 9324
rect 171948 476 172312 480
rect 171948 420 172004 476
rect 171388 364 172004 420
rect 172060 392 172312 476
rect 172088 -960 172312 392
rect 173208 -960 173432 480
rect 174300 392 174552 480
rect 174328 -960 174552 392
rect 174748 420 174804 12796
rect 177212 9716 177268 55412
rect 177212 9650 177268 9660
rect 178108 26068 178164 26078
rect 177660 7588 177716 7598
rect 175308 480 175476 532
rect 177660 480 177716 7532
rect 175308 476 175672 480
rect 175308 420 175364 476
rect 174748 364 175364 420
rect 175420 392 175672 476
rect 175448 -960 175672 392
rect 176568 -960 176792 480
rect 177660 392 177912 480
rect 177688 -960 177912 392
rect 178108 420 178164 26012
rect 179788 21028 179844 21038
rect 179788 20188 179844 20972
rect 179788 20132 180404 20188
rect 178668 480 178836 532
rect 178668 476 179032 480
rect 178668 420 178724 476
rect 178108 364 178724 420
rect 178780 392 179032 476
rect 178808 -960 179032 392
rect 179928 -960 180152 480
rect 180348 420 180404 20132
rect 180460 2548 180516 115388
rect 180572 64820 180628 64830
rect 180572 4116 180628 64764
rect 188860 11172 188916 11182
rect 182364 7700 182420 7710
rect 180572 4050 180628 4060
rect 181468 6020 181524 6030
rect 181468 3556 181524 5964
rect 181468 3490 181524 3500
rect 182140 4116 182196 4126
rect 180460 2482 180516 2492
rect 180908 480 181076 532
rect 182140 480 182196 4060
rect 182364 4116 182420 7644
rect 187740 4452 187796 4462
rect 182364 4050 182420 4060
rect 185500 4116 185556 4126
rect 184380 3556 184436 3566
rect 184380 480 184436 3500
rect 185500 480 185556 4060
rect 187740 480 187796 4396
rect 188860 480 188916 11116
rect 188972 10276 189028 129388
rect 188972 10210 189028 10220
rect 189308 118020 189364 118030
rect 189308 5796 189364 117964
rect 189868 67172 189924 587132
rect 192332 583044 192388 583054
rect 191548 317380 191604 317390
rect 191212 313684 191268 313694
rect 190988 313572 191044 313582
rect 190652 313460 190708 313470
rect 189980 313348 190036 313358
rect 189980 157892 190036 313292
rect 189980 156996 190036 157836
rect 190092 302036 190148 302046
rect 190092 157220 190148 301980
rect 190652 158116 190708 313404
rect 190652 157668 190708 158060
rect 190652 157602 190708 157612
rect 190764 309988 190820 309998
rect 190764 305060 190820 309932
rect 190764 157444 190820 305004
rect 190764 157378 190820 157388
rect 190876 303268 190932 303278
rect 190876 158228 190932 303212
rect 190092 157154 190148 157164
rect 189980 156930 190036 156940
rect 189868 67106 189924 67116
rect 190652 124404 190708 124414
rect 189308 5730 189364 5740
rect 190652 2996 190708 124348
rect 190876 124180 190932 158172
rect 190988 301924 191044 313516
rect 190988 156884 191044 301868
rect 191212 301700 191268 313628
rect 191212 157556 191268 301644
rect 191436 307076 191492 307086
rect 191436 301812 191492 307020
rect 191436 159796 191492 301756
rect 191436 159730 191492 159740
rect 191212 157490 191268 157500
rect 190988 156818 191044 156828
rect 190876 124114 190932 124124
rect 191436 151172 191492 151182
rect 191436 149604 191492 151116
rect 191324 121268 191380 121278
rect 190764 61348 190820 61358
rect 190764 4116 190820 61292
rect 190764 4050 190820 4060
rect 191100 9268 191156 9278
rect 190652 2930 190708 2940
rect 191100 480 191156 9212
rect 191324 3108 191380 121212
rect 191324 3042 191380 3052
rect 191436 2884 191492 149548
rect 191548 128548 191604 317324
rect 191548 128482 191604 128492
rect 191660 306964 191716 306974
rect 191660 121940 191716 306908
rect 191884 306740 191940 306750
rect 191884 305844 191940 306684
rect 191884 154308 191940 305788
rect 191884 154242 191940 154252
rect 191660 121268 191716 121884
rect 191660 121202 191716 121212
rect 192332 69076 192388 582988
rect 194012 561204 194068 561214
rect 192332 69010 192388 69020
rect 192444 461188 192500 461198
rect 192444 67060 192500 461132
rect 192556 317604 192612 317614
rect 192556 68628 192612 317548
rect 193116 306852 193172 306862
rect 193116 305172 193172 306796
rect 193116 305106 193172 305116
rect 193900 304164 193956 304174
rect 192668 302148 192724 302158
rect 192668 151172 192724 302092
rect 193900 153748 193956 304108
rect 194012 156212 194068 561148
rect 194124 517524 194180 517534
rect 194124 159572 194180 517468
rect 196476 319172 196532 587356
rect 222236 587412 222292 591560
rect 222236 587346 222292 587356
rect 402108 587300 402164 591560
rect 402108 587234 402164 587244
rect 467516 587188 467572 591560
rect 467516 587122 467572 587132
rect 532588 461188 532644 591612
rect 532812 591556 532868 591612
rect 532924 591560 533176 591640
rect 549304 591560 549528 593000
rect 565656 591560 565880 593000
rect 582008 591560 582232 593000
rect 532924 591556 532980 591560
rect 532812 591500 532980 591556
rect 532588 461122 532644 461132
rect 589820 484372 589876 484382
rect 587132 451108 587188 451118
rect 202300 319284 202356 320040
rect 202300 319218 202356 319228
rect 196476 319106 196532 319116
rect 206108 319172 206164 320040
rect 206108 319106 206164 319116
rect 208348 320012 209944 320068
rect 213388 320012 213752 320068
rect 216748 320012 217560 320068
rect 220108 320012 221368 320068
rect 194684 317044 194740 317054
rect 194124 159506 194180 159516
rect 194236 311668 194292 311678
rect 194012 156146 194068 156156
rect 193900 153682 193956 153692
rect 193228 152964 193284 152974
rect 193228 152292 193284 152908
rect 193228 152226 193284 152236
rect 192668 151106 192724 151116
rect 194012 127764 194068 127774
rect 193004 126308 193060 126318
rect 192556 68562 192612 68572
rect 192668 126196 192724 126206
rect 192444 66994 192500 67004
rect 191436 2818 191492 2828
rect 191548 63028 191604 63038
rect 180908 476 181272 480
rect 180908 420 180964 476
rect 180348 364 180964 420
rect 181020 392 181272 476
rect 182140 392 182392 480
rect 181048 -960 181272 392
rect 182168 -960 182392 392
rect 183288 -960 183512 480
rect 184380 392 184632 480
rect 185500 392 185752 480
rect 184408 -960 184632 392
rect 185528 -960 185752 392
rect 186648 -960 186872 480
rect 187740 392 187992 480
rect 188860 392 189112 480
rect 187768 -960 187992 392
rect 188888 -960 189112 392
rect 190008 -960 190232 480
rect 191100 392 191352 480
rect 191128 -960 191352 392
rect 191548 420 191604 62972
rect 192668 756 192724 126140
rect 192892 124516 192948 124526
rect 192892 1540 192948 124460
rect 193004 6580 193060 126252
rect 193004 6514 193060 6524
rect 193116 119364 193172 119374
rect 192892 1474 192948 1484
rect 193116 1428 193172 119308
rect 193900 117684 193956 117694
rect 193900 7924 193956 117628
rect 193900 7858 193956 7868
rect 193116 1362 193172 1372
rect 194012 1204 194068 127708
rect 194124 118132 194180 118142
rect 194124 7140 194180 118076
rect 194236 66948 194292 311612
rect 194572 303268 194628 303278
rect 194236 66882 194292 66892
rect 194348 301588 194404 301598
rect 194348 63812 194404 301532
rect 194348 63746 194404 63756
rect 194460 124404 194516 124414
rect 194460 13300 194516 124348
rect 194572 118692 194628 303212
rect 194684 121828 194740 316988
rect 195692 315028 195748 315038
rect 194908 159236 194964 159246
rect 194908 158340 194964 159180
rect 195692 159012 195748 314972
rect 197932 313908 197988 313918
rect 197036 313460 197092 313470
rect 196364 306852 196420 306862
rect 196252 306740 196308 306750
rect 195692 158946 195748 158956
rect 195916 168644 195972 168654
rect 195916 159124 195972 168588
rect 194908 158274 194964 158284
rect 195804 154420 195860 154430
rect 195692 153636 195748 153646
rect 195468 151172 195524 151182
rect 194908 148260 194964 148270
rect 194908 147924 194964 148204
rect 194908 147858 194964 147868
rect 194684 121762 194740 121772
rect 194908 122612 194964 122622
rect 194908 121380 194964 122556
rect 194908 121314 194964 121324
rect 194572 118626 194628 118636
rect 194684 121156 194740 121166
rect 194460 13234 194516 13244
rect 194572 116788 194628 116798
rect 194572 9940 194628 116732
rect 194572 9874 194628 9884
rect 194124 7074 194180 7084
rect 194012 1138 194068 1148
rect 194460 4116 194516 4126
rect 192668 690 192724 700
rect 192108 480 192276 532
rect 194460 480 194516 4060
rect 194684 1316 194740 121100
rect 194796 120036 194852 120046
rect 194796 119700 194852 119980
rect 195468 120036 195524 151116
rect 195468 119970 195524 119980
rect 195692 149716 195748 153580
rect 194796 4788 194852 119644
rect 195468 116452 195524 116462
rect 194796 4722 194852 4732
rect 194908 12740 194964 12750
rect 194684 1250 194740 1260
rect 192108 476 192472 480
rect 192108 420 192164 476
rect 191548 364 192164 420
rect 192220 392 192472 476
rect 192248 -960 192472 392
rect 193368 -960 193592 480
rect 194460 392 194712 480
rect 194488 -960 194712 392
rect 194908 420 194964 12684
rect 195468 7252 195524 116396
rect 195468 7186 195524 7196
rect 195692 4452 195748 149660
rect 195804 124404 195860 154364
rect 195804 124338 195860 124348
rect 195804 122724 195860 122734
rect 195804 9828 195860 122668
rect 195804 9762 195860 9772
rect 195916 6468 195972 159068
rect 196028 155876 196084 155886
rect 196028 138852 196084 155820
rect 196252 154420 196308 306684
rect 196252 154354 196308 154364
rect 196364 151172 196420 306796
rect 196364 151106 196420 151116
rect 196476 169092 196532 169102
rect 196476 158340 196532 169036
rect 196028 138786 196084 138796
rect 196140 148036 196196 148046
rect 196028 121380 196084 121390
rect 196028 10500 196084 121324
rect 196140 13412 196196 147980
rect 196364 147924 196420 147934
rect 196140 13346 196196 13356
rect 196252 146468 196308 146478
rect 196028 10434 196084 10444
rect 196252 8708 196308 146412
rect 196252 8642 196308 8652
rect 196364 7588 196420 147868
rect 196364 7522 196420 7532
rect 195916 6402 195972 6412
rect 195692 4386 195748 4396
rect 196476 2772 196532 158284
rect 197036 152516 197092 313404
rect 197484 310436 197540 310446
rect 197372 309988 197428 309998
rect 197372 168084 197428 309932
rect 197372 168018 197428 168028
rect 197484 159796 197540 310380
rect 197820 310324 197876 310334
rect 197708 303716 197764 303726
rect 197372 158452 197428 158462
rect 197036 152450 197092 152460
rect 197148 157220 197204 157230
rect 196588 152292 196644 152302
rect 196588 142212 196644 152236
rect 196588 142146 196644 142156
rect 197148 141988 197204 157164
rect 197148 141922 197204 141932
rect 197260 154532 197316 154542
rect 197260 153076 197316 154476
rect 197260 122612 197316 153020
rect 197260 122546 197316 122556
rect 197372 146356 197428 158396
rect 196588 14308 196644 14318
rect 196588 4116 196644 14252
rect 197372 6244 197428 146300
rect 197484 142884 197540 159740
rect 197596 303492 197652 303502
rect 197596 154532 197652 303436
rect 197596 154466 197652 154476
rect 197484 137788 197540 142828
rect 197708 151396 197764 303660
rect 197820 153636 197876 310268
rect 197820 153570 197876 153580
rect 197932 156100 197988 313852
rect 208348 313908 208404 320012
rect 208348 313842 208404 313852
rect 197484 137732 197652 137788
rect 197372 6178 197428 6188
rect 197484 131236 197540 131246
rect 196588 4050 196644 4060
rect 197484 3220 197540 131180
rect 197596 6132 197652 137732
rect 197596 6066 197652 6076
rect 197708 119588 197764 151340
rect 197484 3154 197540 3164
rect 196476 2706 196532 2716
rect 197708 868 197764 119532
rect 197820 151060 197876 151070
rect 197820 118468 197876 151004
rect 197932 147924 197988 156044
rect 197932 147858 197988 147868
rect 198044 313796 198100 313806
rect 198044 152852 198100 313740
rect 213388 313796 213444 320012
rect 213388 313730 213444 313740
rect 199164 313684 199220 313694
rect 199052 310212 199108 310222
rect 198828 306964 198884 306974
rect 198716 302260 198772 302270
rect 198156 178052 198212 178062
rect 198156 160132 198212 177996
rect 198716 178052 198772 302204
rect 198716 177986 198772 177996
rect 198156 159684 198212 160076
rect 198156 159618 198212 159628
rect 198268 161364 198324 161374
rect 198268 157332 198324 161308
rect 198268 157266 198324 157276
rect 198716 159684 198772 159694
rect 198044 146468 198100 152796
rect 198380 152404 198436 152414
rect 198380 148932 198436 152348
rect 198380 148866 198436 148876
rect 198716 148036 198772 159628
rect 198716 147970 198772 147980
rect 198828 156548 198884 306908
rect 198940 303604 198996 303614
rect 198940 156548 198996 303548
rect 199052 159460 199108 310156
rect 199164 159684 199220 313628
rect 216748 313684 216804 320012
rect 216748 313618 216804 313628
rect 199388 313572 199444 313582
rect 199164 159618 199220 159628
rect 199276 311892 199332 311902
rect 199276 159908 199332 311836
rect 199052 158452 199108 159404
rect 199052 158386 199108 158396
rect 198940 156492 199220 156548
rect 198044 146402 198100 146412
rect 198156 142996 198212 143006
rect 197820 118402 197876 118412
rect 197932 119476 197988 119486
rect 197820 116228 197876 116238
rect 197820 8428 197876 116172
rect 197932 9268 197988 119420
rect 197932 9202 197988 9212
rect 198044 104132 198100 104142
rect 197820 8372 197988 8428
rect 197708 802 197764 812
rect 197820 4116 197876 4126
rect 195468 480 195636 532
rect 197820 480 197876 4060
rect 197932 2660 197988 8372
rect 197932 2594 197988 2604
rect 198044 1092 198100 104076
rect 198156 8484 198212 142940
rect 198828 142996 198884 156492
rect 198828 142930 198884 142940
rect 199052 156324 199108 156334
rect 199052 146244 199108 156268
rect 198492 13412 198548 13422
rect 198156 8418 198212 8428
rect 198268 10276 198324 10286
rect 198268 1652 198324 10220
rect 198492 8596 198548 13356
rect 198828 13300 198884 13310
rect 198492 8530 198548 8540
rect 198604 12628 198660 12638
rect 198604 4564 198660 12572
rect 198604 4498 198660 4508
rect 198828 2548 198884 13244
rect 198828 2482 198884 2492
rect 198940 10948 198996 10958
rect 198268 1586 198324 1596
rect 198044 1026 198100 1036
rect 198940 480 198996 10892
rect 199052 3892 199108 146188
rect 199164 153188 199220 156492
rect 199164 122836 199220 153132
rect 199276 149548 199332 159852
rect 199388 157668 199444 313516
rect 220108 313572 220164 320012
rect 220108 313506 220164 313516
rect 225148 310436 225204 320040
rect 225148 310370 225204 310380
rect 228508 320012 228984 320068
rect 231868 320012 232792 320068
rect 235228 320012 236600 320068
rect 228508 310324 228564 320012
rect 228508 310258 228564 310268
rect 231868 310212 231924 320012
rect 231868 310146 231924 310156
rect 235228 306964 235284 320012
rect 240380 314188 240436 320040
rect 240268 314132 240436 314188
rect 243628 320012 244216 320068
rect 246988 320012 248024 320068
rect 250348 320012 251832 320068
rect 255388 320012 255640 320068
rect 258748 320012 259448 320068
rect 262108 320012 263256 320068
rect 265468 320012 267064 320068
rect 270508 320012 270872 320068
rect 273868 320012 274680 320068
rect 277228 320012 278488 320068
rect 240268 311892 240324 314132
rect 240268 311826 240324 311836
rect 235228 306898 235284 306908
rect 243628 303716 243684 320012
rect 243628 303650 243684 303660
rect 246988 303604 247044 320012
rect 246988 303538 247044 303548
rect 250348 303492 250404 320012
rect 255388 313460 255444 320012
rect 255388 313394 255444 313404
rect 250348 303426 250404 303436
rect 258748 302260 258804 320012
rect 262108 306852 262164 320012
rect 262108 306786 262164 306796
rect 265468 306740 265524 320012
rect 270508 310100 270564 320012
rect 270508 310034 270564 310044
rect 273868 309988 273924 320012
rect 273868 309922 273924 309932
rect 265468 306674 265524 306684
rect 258748 302194 258804 302204
rect 277228 302148 277284 320012
rect 282268 313348 282324 320040
rect 282268 313282 282324 313292
rect 285628 320012 286104 320068
rect 285628 305284 285684 320012
rect 289884 315140 289940 320040
rect 289884 315074 289940 315084
rect 292348 320012 293720 320068
rect 285628 305218 285684 305228
rect 292348 305172 292404 320012
rect 297500 314188 297556 320040
rect 297388 314132 297556 314188
rect 300748 320012 301336 320068
rect 304108 320012 305144 320068
rect 297388 309988 297444 314132
rect 300748 310100 300804 320012
rect 304108 310212 304164 320012
rect 308924 317044 308980 320040
rect 308924 316978 308980 316988
rect 312508 320012 312760 320068
rect 315868 320012 316568 320068
rect 319228 320012 320376 320068
rect 322588 320012 324184 320068
rect 327628 320012 327992 320068
rect 330988 320012 331800 320068
rect 334348 320012 335608 320068
rect 304108 310146 304164 310156
rect 300748 310034 300804 310044
rect 297388 309922 297444 309932
rect 312508 306740 312564 320012
rect 312508 306674 312564 306684
rect 292348 305106 292404 305116
rect 315868 303492 315924 320012
rect 319228 313348 319284 320012
rect 319228 313282 319284 313292
rect 315868 303426 315924 303436
rect 322588 303380 322644 320012
rect 327628 313460 327684 320012
rect 330988 313572 331044 320012
rect 330988 313506 331044 313516
rect 327628 313394 327684 313404
rect 334348 303604 334404 320012
rect 339388 316932 339444 320040
rect 339388 316866 339444 316876
rect 342748 320012 343224 320068
rect 342748 313684 342804 320012
rect 347004 317044 347060 320040
rect 347004 316978 347060 316988
rect 350812 316932 350868 320040
rect 354620 317156 354676 320040
rect 354620 317090 354676 317100
rect 357868 320012 358456 320068
rect 350812 316866 350868 316876
rect 342748 313618 342804 313628
rect 357868 312564 357924 320012
rect 357868 308420 357924 312508
rect 361228 315924 361284 315934
rect 361228 311780 361284 315868
rect 362236 315924 362292 320040
rect 366044 316820 366100 320040
rect 366044 316754 366100 316764
rect 369628 320012 369880 320068
rect 372988 320012 373688 320068
rect 403368 320012 404068 320068
rect 407176 320012 407764 320068
rect 362236 315858 362292 315868
rect 361228 311714 361284 311724
rect 357868 308354 357924 308364
rect 334348 303538 334404 303548
rect 322588 303314 322644 303324
rect 277228 302082 277284 302092
rect 369628 302036 369684 320012
rect 372988 303268 373044 320012
rect 404012 319172 404068 320012
rect 404012 319106 404068 319116
rect 397852 317268 397908 317278
rect 378140 317156 378196 317166
rect 372988 303202 373044 303212
rect 376348 313572 376404 313582
rect 376348 302596 376404 313516
rect 378028 313460 378084 313470
rect 376348 302530 376404 302540
rect 377020 313348 377076 313358
rect 369628 301970 369684 301980
rect 301308 160244 301364 160254
rect 218204 160132 218260 160142
rect 202300 159572 202356 160104
rect 202300 159506 202356 159516
rect 199388 156324 199444 157612
rect 199388 156258 199444 156268
rect 199948 159012 200004 159022
rect 199388 151284 199444 151294
rect 199388 150388 199444 151228
rect 199948 151284 200004 158956
rect 202524 156436 202580 156446
rect 201180 153076 201236 153086
rect 201180 152740 201236 153020
rect 201180 152674 201236 152684
rect 199948 151218 200004 151228
rect 202524 151060 202580 156380
rect 206108 156212 206164 160104
rect 206892 158340 206948 158350
rect 206108 156146 206164 156156
rect 206668 158228 206724 158238
rect 206668 156212 206724 158172
rect 206668 156146 206724 156156
rect 206780 156324 206836 156334
rect 206780 154420 206836 156268
rect 206780 154354 206836 154364
rect 202524 150994 202580 151004
rect 203308 154196 203364 154206
rect 203308 150612 203364 154140
rect 204988 152964 205044 152974
rect 204988 151956 205044 152908
rect 204988 151890 205044 151900
rect 206892 150836 206948 158284
rect 207004 156548 207060 156558
rect 207004 154532 207060 156492
rect 209916 156100 209972 160104
rect 213724 156884 213780 160104
rect 217532 159572 217588 160104
rect 217532 159506 217588 159516
rect 269388 160132 269444 160142
rect 218204 159572 218260 160076
rect 218204 159506 218260 159516
rect 213724 156818 213780 156828
rect 213948 158228 214004 158238
rect 209916 156034 209972 156044
rect 213052 156324 213108 156334
rect 207004 154466 207060 154476
rect 209356 154532 209412 154542
rect 209356 150948 209412 154476
rect 209916 154308 209972 154318
rect 209916 151172 209972 154252
rect 213052 154084 213108 156268
rect 213052 154018 213108 154028
rect 209916 151106 209972 151116
rect 213948 151060 214004 158172
rect 221340 157668 221396 160104
rect 225148 159796 225204 160104
rect 225148 159730 225204 159740
rect 226828 160020 226884 160030
rect 221340 157602 221396 157612
rect 225260 159684 225316 159694
rect 223804 157332 223860 157342
rect 215068 153972 215124 153982
rect 215068 152852 215124 153916
rect 213948 150994 214004 151004
rect 214956 152796 215124 152852
rect 209356 150882 209412 150892
rect 206892 150770 206948 150780
rect 214956 150836 215012 152796
rect 223356 152740 223412 152750
rect 215068 152628 215124 152638
rect 215068 151060 215124 152572
rect 216748 152628 216804 152638
rect 216748 151172 216804 152572
rect 216748 151106 216804 151116
rect 223356 151172 223412 152684
rect 223804 152740 223860 157276
rect 223804 152674 223860 152684
rect 223356 151106 223412 151116
rect 215068 150994 215124 151004
rect 225260 150948 225316 159628
rect 226828 157332 226884 159964
rect 226828 157266 226884 157276
rect 228508 159796 228564 159806
rect 225260 150882 225316 150892
rect 225484 151956 225540 151966
rect 225484 150948 225540 151900
rect 228508 151060 228564 159740
rect 228956 153636 229012 160104
rect 232764 159460 232820 160104
rect 236572 159684 236628 160104
rect 240380 159908 240436 160104
rect 240380 159842 240436 159852
rect 236572 159618 236628 159628
rect 232764 159394 232820 159404
rect 230300 159124 230356 159134
rect 230188 158228 230244 158238
rect 230188 154420 230244 158172
rect 230188 154354 230244 154364
rect 230300 154196 230356 159068
rect 238812 158228 238868 158238
rect 230300 154130 230356 154140
rect 238700 154196 238756 154206
rect 228956 153570 229012 153580
rect 238588 154084 238644 154094
rect 238588 151172 238644 154028
rect 238588 151106 238644 151116
rect 228508 150994 228564 151004
rect 238700 151060 238756 154140
rect 238700 150994 238756 151004
rect 225484 150882 225540 150892
rect 238812 150948 238868 158172
rect 244188 152628 244244 160104
rect 247996 152852 248052 160104
rect 251804 154084 251860 160104
rect 251804 154018 251860 154028
rect 252028 158116 252084 158126
rect 247996 152786 248052 152796
rect 244188 152562 244244 152572
rect 252028 151172 252084 158060
rect 253820 158116 253876 158126
rect 253708 154308 253764 154318
rect 253708 152852 253764 154252
rect 253708 152786 253764 152796
rect 253820 152740 253876 158060
rect 253820 152674 253876 152684
rect 252028 151106 252084 151116
rect 253708 152628 253764 152638
rect 253708 151060 253764 152572
rect 255612 152516 255668 160104
rect 259420 159572 259476 160104
rect 259420 159506 259476 159516
rect 260764 154644 260820 154654
rect 260764 152740 260820 154588
rect 262108 154644 262164 154654
rect 262108 153860 262164 154588
rect 262108 153794 262164 153804
rect 263228 152852 263284 160104
rect 263788 159236 263844 159246
rect 263788 153972 263844 159180
rect 263788 153906 263844 153916
rect 263900 158228 263956 158238
rect 263228 152786 263284 152796
rect 263900 152852 263956 158172
rect 263900 152786 263956 152796
rect 260764 152674 260820 152684
rect 267036 152628 267092 160104
rect 274652 160132 274708 160142
rect 269276 158116 269332 158126
rect 269276 154308 269332 158060
rect 269388 155988 269444 160076
rect 270844 157668 270900 160104
rect 297500 160132 297556 160142
rect 274652 160066 274708 160076
rect 270844 157602 270900 157612
rect 269388 155922 269444 155932
rect 270396 156436 270452 156446
rect 269276 154242 269332 154252
rect 270396 154084 270452 156380
rect 270396 154018 270452 154028
rect 278460 153860 278516 160104
rect 282268 159236 282324 160104
rect 286076 159796 286132 160104
rect 286076 159730 286132 159740
rect 282268 159170 282324 159180
rect 285628 158228 285684 158238
rect 283836 158116 283892 158126
rect 283836 157668 283892 158060
rect 283836 157602 283892 157612
rect 282156 156100 282212 156110
rect 282156 154308 282212 156044
rect 285628 156100 285684 158172
rect 285628 156034 285684 156044
rect 289884 154420 289940 160104
rect 293692 157444 293748 160104
rect 297500 160066 297556 160076
rect 300748 159796 300804 159806
rect 300748 157780 300804 159740
rect 300748 157714 300804 157724
rect 301308 157556 301364 160188
rect 301308 157490 301364 157500
rect 304444 160132 304500 160142
rect 293692 157378 293748 157388
rect 289884 154354 289940 154364
rect 294252 156324 294308 156334
rect 294252 154420 294308 156268
rect 294252 154354 294308 154364
rect 282156 154242 282212 154252
rect 304444 154308 304500 160076
rect 305116 157892 305172 160104
rect 308924 159124 308980 160104
rect 312760 160076 313460 160132
rect 313404 159684 313460 160076
rect 313404 159618 313460 159628
rect 308924 159058 308980 159068
rect 305116 157668 305172 157836
rect 309148 158228 309204 158238
rect 309148 157892 309204 158172
rect 309148 157826 309204 157836
rect 315420 158228 315476 158238
rect 305116 157602 305172 157612
rect 304444 154242 304500 154252
rect 278460 153794 278516 153804
rect 283388 153860 283444 153870
rect 267036 152562 267092 152572
rect 255612 152450 255668 152460
rect 283388 152516 283444 153804
rect 283388 152450 283444 152460
rect 315420 151172 315476 158172
rect 316540 154420 316596 160104
rect 320348 157892 320404 160104
rect 320348 157826 320404 157836
rect 320012 157556 320068 157566
rect 320012 155988 320068 157500
rect 320012 155922 320068 155932
rect 316540 154354 316596 154364
rect 319116 154644 319172 154654
rect 319116 154196 319172 154588
rect 319116 154130 319172 154140
rect 315420 151106 315476 151116
rect 317212 153412 317268 153422
rect 317212 151172 317268 153356
rect 324156 152628 324212 160104
rect 327964 159460 328020 160104
rect 327964 159394 328020 159404
rect 330652 159908 330708 159918
rect 329756 158116 329812 158126
rect 329756 156100 329812 158060
rect 330652 157668 330708 159852
rect 330876 159684 330932 159694
rect 330876 159124 330932 159628
rect 331772 159684 331828 160104
rect 335580 159796 335636 160104
rect 335580 159730 335636 159740
rect 331772 159618 331828 159628
rect 330876 159058 330932 159068
rect 330652 157602 330708 157612
rect 339388 157220 339444 160104
rect 343196 158228 343252 160104
rect 346108 160020 346164 160030
rect 346108 159460 346164 159964
rect 347004 159572 347060 160104
rect 347004 159506 347060 159516
rect 346108 159394 346164 159404
rect 350812 159236 350868 160104
rect 350812 159170 350868 159180
rect 343196 157780 343252 158172
rect 343196 157714 343252 157724
rect 354620 157668 354676 160104
rect 354620 157602 354676 157612
rect 358428 157556 358484 160104
rect 358428 157490 358484 157500
rect 359548 157444 359604 157454
rect 339388 157154 339444 157164
rect 356188 157332 356244 157342
rect 329756 156034 329812 156044
rect 332668 156436 332724 156446
rect 324156 152562 324212 152572
rect 332668 152628 332724 156380
rect 348012 156436 348068 156446
rect 344652 156324 344708 156334
rect 343308 156100 343364 156110
rect 343196 155988 343252 155998
rect 342188 154644 342244 154654
rect 342188 154196 342244 154588
rect 342188 154130 342244 154140
rect 343196 154196 343252 155932
rect 343196 154130 343252 154140
rect 343308 153972 343364 156044
rect 344652 154308 344708 156268
rect 347900 156212 347956 156222
rect 348012 156212 348068 156380
rect 347956 156156 348068 156212
rect 356188 156212 356244 157276
rect 357980 157220 358036 157230
rect 347900 156146 347956 156156
rect 356188 156146 356244 156156
rect 357868 156436 357924 156446
rect 357868 156100 357924 156380
rect 357868 156034 357924 156044
rect 357980 155876 358036 157164
rect 357980 155810 358036 155820
rect 359548 155876 359604 157388
rect 362236 157444 362292 160104
rect 366044 159012 366100 160104
rect 366044 158946 366100 158956
rect 362236 157378 362292 157388
rect 369852 156996 369908 160104
rect 369852 156930 369908 156940
rect 359548 155810 359604 155820
rect 344652 154242 344708 154252
rect 343308 153906 343364 153916
rect 359548 153860 359604 153870
rect 359548 152740 359604 153804
rect 359548 152674 359604 152684
rect 362796 153300 362852 153310
rect 362796 152740 362852 153244
rect 362796 152674 362852 152684
rect 332668 152562 332724 152572
rect 317212 151106 317268 151116
rect 363356 152516 363412 152526
rect 253708 150994 253764 151004
rect 238812 150882 238868 150892
rect 214956 150770 215012 150780
rect 203308 150546 203364 150556
rect 363356 150612 363412 152460
rect 373660 152404 373716 160104
rect 377020 157892 377076 313292
rect 377020 156324 377076 157836
rect 377020 156258 377076 156268
rect 377132 310100 377188 310110
rect 373660 152338 373716 152348
rect 377132 154196 377188 310044
rect 377468 303604 377524 303614
rect 377244 303380 377300 303390
rect 377244 156100 377300 303324
rect 377356 302596 377412 302606
rect 377356 159684 377412 302540
rect 377356 156884 377412 159628
rect 377468 159796 377524 303548
rect 378028 302484 378084 313404
rect 378140 305732 378196 317100
rect 378140 305666 378196 305676
rect 378252 317044 378308 317054
rect 378028 302418 378084 302428
rect 378252 301924 378308 316988
rect 383068 316932 383124 316942
rect 379708 315924 379764 315934
rect 379036 313684 379092 313694
rect 378252 300916 378308 301868
rect 378252 300850 378308 300860
rect 378364 310212 378420 310222
rect 378364 160916 378420 310156
rect 378364 160850 378420 160860
rect 378588 305732 378644 305742
rect 378588 305060 378644 305676
rect 377468 157332 377524 159740
rect 378140 160020 378196 160030
rect 378140 159684 378196 159964
rect 377468 157266 377524 157276
rect 378028 159124 378084 159134
rect 378028 158116 378084 159068
rect 377356 156828 377636 156884
rect 377244 156034 377300 156044
rect 377356 156324 377412 156334
rect 363356 150546 363412 150556
rect 199388 150322 199444 150332
rect 377132 149548 377188 154140
rect 199276 149492 199444 149548
rect 377132 149492 377300 149548
rect 199164 7812 199220 122780
rect 199388 144564 199444 149492
rect 199164 7746 199220 7756
rect 199276 17668 199332 17678
rect 199276 4340 199332 17612
rect 199388 6804 199444 144508
rect 203196 10500 203252 10510
rect 200172 10388 200228 10398
rect 200172 7476 200228 10332
rect 202300 8372 202356 10136
rect 202300 8306 202356 8316
rect 200172 7410 200228 7420
rect 203196 6916 203252 10444
rect 203196 6850 203252 6860
rect 205100 9604 205156 9614
rect 199388 6738 199444 6748
rect 199948 6804 200004 6814
rect 199948 4676 200004 6748
rect 199948 4610 200004 4620
rect 204540 5908 204596 5918
rect 199276 4274 199332 4284
rect 202300 4340 202356 4350
rect 199052 3826 199108 3836
rect 201180 4116 201236 4126
rect 201180 480 201236 4060
rect 202300 480 202356 4284
rect 204540 480 204596 5852
rect 205100 5908 205156 9548
rect 206108 8260 206164 10136
rect 206108 8194 206164 8204
rect 209916 7588 209972 10136
rect 213724 8708 213780 10136
rect 213724 8642 213780 8652
rect 217532 8596 217588 10136
rect 217532 8530 217588 8540
rect 209916 7522 209972 7532
rect 206780 6916 206836 6926
rect 205100 5842 205156 5852
rect 206668 6804 206724 6814
rect 206668 5796 206724 6748
rect 206668 5730 206724 5740
rect 206780 4676 206836 6860
rect 206780 4610 206836 4620
rect 205660 4564 205716 4574
rect 204988 4228 205044 4238
rect 204988 3220 205044 4172
rect 204988 3154 205044 3164
rect 205212 3220 205268 3230
rect 205212 2660 205268 3164
rect 205548 2660 205604 2670
rect 205212 2594 205268 2604
rect 205324 2604 205548 2660
rect 205324 2548 205380 2604
rect 205548 2594 205604 2604
rect 205324 2482 205380 2492
rect 205660 480 205716 4508
rect 221340 3892 221396 10136
rect 225148 6132 225204 10136
rect 225148 6066 225204 6076
rect 223356 5908 223412 5918
rect 223356 5012 223412 5852
rect 223356 4946 223412 4956
rect 224924 5124 224980 5134
rect 221340 3826 221396 3836
rect 207900 3780 207956 3790
rect 207900 480 207956 3724
rect 224924 1652 224980 5068
rect 228956 4452 229012 10136
rect 232764 6244 232820 10136
rect 236572 8484 236628 10136
rect 236572 8418 236628 8428
rect 232764 6178 232820 6188
rect 228956 4386 229012 4396
rect 230188 6020 230244 6030
rect 230188 4452 230244 5964
rect 230300 5236 230356 5246
rect 230300 5012 230356 5180
rect 230300 4946 230356 4956
rect 240380 4564 240436 10136
rect 240380 4498 240436 4508
rect 230188 4386 230244 4396
rect 224924 1586 224980 1596
rect 244188 868 244244 10136
rect 247996 7812 248052 10136
rect 247996 7746 248052 7756
rect 251804 4676 251860 10136
rect 251804 4610 251860 4620
rect 255612 4452 255668 10136
rect 259420 6356 259476 10136
rect 259420 6290 259476 6300
rect 263228 4788 263284 10136
rect 263228 4722 263284 4732
rect 255612 4386 255668 4396
rect 267036 2660 267092 10136
rect 270844 6468 270900 10136
rect 270844 6402 270900 6412
rect 274652 4900 274708 10136
rect 274652 4834 274708 4844
rect 277228 4900 277284 4910
rect 277228 2884 277284 4844
rect 278460 4900 278516 10136
rect 278460 4834 278516 4844
rect 277228 2818 277284 2828
rect 282268 2772 282324 10136
rect 286076 2996 286132 10136
rect 286076 2930 286132 2940
rect 282268 2706 282324 2716
rect 267036 2594 267092 2604
rect 289884 980 289940 10136
rect 293692 2996 293748 10136
rect 297500 8428 297556 10136
rect 297388 8372 297556 8428
rect 297388 6356 297444 8372
rect 297388 6020 297444 6300
rect 297276 5964 297444 6020
rect 297276 3108 297332 5964
rect 301308 4788 301364 10136
rect 301308 4722 301364 4732
rect 305116 4676 305172 10136
rect 308924 7924 308980 10136
rect 308924 7858 308980 7868
rect 312732 6244 312788 10136
rect 312732 6178 312788 6188
rect 316540 6132 316596 10136
rect 320348 8596 320404 10136
rect 320348 8530 320404 8540
rect 316540 6066 316596 6076
rect 305116 4610 305172 4620
rect 314972 5236 315028 5246
rect 297276 3042 297332 3052
rect 314972 3108 315028 5180
rect 324156 4564 324212 10136
rect 327964 8260 328020 10136
rect 327964 8194 328020 8204
rect 324156 4498 324212 4508
rect 331772 4452 331828 10136
rect 335580 9716 335636 10136
rect 335580 8484 335636 9660
rect 335580 8418 335636 8428
rect 339388 7476 339444 10136
rect 339388 7410 339444 7420
rect 343196 6020 343252 10136
rect 347004 7924 347060 10136
rect 347004 7858 347060 7868
rect 347788 9268 347844 9278
rect 343196 5954 343252 5964
rect 331772 4386 331828 4396
rect 341628 5124 341684 5134
rect 314972 3042 315028 3052
rect 330204 3444 330260 3454
rect 293692 1092 293748 2940
rect 330204 2884 330260 3388
rect 330204 2818 330260 2828
rect 293692 1026 293748 1036
rect 341628 1092 341684 5068
rect 347788 2772 347844 9212
rect 350812 8708 350868 10136
rect 350812 8642 350868 8652
rect 354620 7812 354676 10136
rect 358428 8036 358484 10136
rect 362236 8148 362292 10136
rect 362236 8082 362292 8092
rect 358428 7970 358484 7980
rect 354620 7746 354676 7756
rect 366044 7140 366100 10136
rect 369852 8372 369908 10136
rect 369852 8306 369908 8316
rect 373660 7252 373716 10136
rect 373660 7186 373716 7196
rect 366044 7074 366100 7084
rect 356188 6804 356244 6814
rect 347788 2706 347844 2716
rect 352604 5908 352660 5918
rect 341628 1026 341684 1036
rect 289884 914 289940 924
rect 244188 802 244244 812
rect 352604 480 352660 5852
rect 356188 2660 356244 6748
rect 377244 4788 377300 149492
rect 377356 8596 377412 156268
rect 377356 8530 377412 8540
rect 377468 156100 377524 156110
rect 377244 4722 377300 4732
rect 377468 4564 377524 156044
rect 377468 4498 377524 4508
rect 377580 4452 377636 156828
rect 378028 6244 378084 158060
rect 378140 8260 378196 159628
rect 378476 159236 378532 159246
rect 378364 158228 378420 158238
rect 378140 8194 378196 8204
rect 378252 156436 378308 156446
rect 378028 6178 378084 6188
rect 378252 6020 378308 156380
rect 378364 7924 378420 158172
rect 378476 8708 378532 159180
rect 378476 8642 378532 8652
rect 378588 157668 378644 305004
rect 378812 302484 378868 302494
rect 378700 300916 378756 300926
rect 378700 159572 378756 300860
rect 378812 159684 378868 302428
rect 378812 159618 378868 159628
rect 378924 302036 378980 302046
rect 378700 158228 378756 159516
rect 378700 158162 378756 158172
rect 378364 7858 378420 7868
rect 378588 7812 378644 157612
rect 378924 156996 378980 301980
rect 378588 7746 378644 7756
rect 378700 154420 378756 154430
rect 378700 6132 378756 154364
rect 378812 153972 378868 153982
rect 378812 6468 378868 153916
rect 378924 152628 378980 156940
rect 379036 157780 379092 313628
rect 379036 156436 379092 157724
rect 379036 156370 379092 156380
rect 379148 312564 379204 312574
rect 379148 157556 379204 312508
rect 379148 156100 379204 157500
rect 379148 156034 379204 156044
rect 379260 303492 379316 303502
rect 379260 154420 379316 303436
rect 379260 154354 379316 154364
rect 379708 157444 379764 315868
rect 379820 306740 379876 306750
rect 379820 301812 379876 306684
rect 379820 158116 379876 301756
rect 383068 301700 383124 316876
rect 397628 313796 397684 313806
rect 397516 313684 397572 313694
rect 397404 310436 397460 310446
rect 383068 159236 383124 301644
rect 383068 159170 383124 159180
rect 396396 306740 396452 306750
rect 379820 158050 379876 158060
rect 379708 154420 379764 157388
rect 388892 157332 388948 157342
rect 379708 154354 379764 154364
rect 383068 156100 383124 156110
rect 378924 152562 378980 152572
rect 379708 152628 379764 152638
rect 378812 6402 378868 6412
rect 378924 150612 378980 150622
rect 378700 6066 378756 6076
rect 378252 5954 378308 5964
rect 378924 4900 378980 150556
rect 379708 8372 379764 152572
rect 379708 8306 379764 8316
rect 383068 8036 383124 156044
rect 386428 154420 386484 154430
rect 386428 8148 386484 154364
rect 388892 67284 388948 157276
rect 388892 67218 388948 67228
rect 395612 104132 395668 104142
rect 386428 8082 386484 8092
rect 383068 7970 383124 7980
rect 378924 4834 378980 4844
rect 377580 4386 377636 4396
rect 356188 2594 356244 2604
rect 395612 1204 395668 104076
rect 396396 104132 396452 306684
rect 397180 303604 397236 303614
rect 397180 161308 397236 303548
rect 396396 104066 396452 104076
rect 397068 161252 397236 161308
rect 397292 303492 397348 303502
rect 397068 159684 397124 161252
rect 395612 1138 395668 1148
rect 397068 1092 397124 159628
rect 397292 159348 397348 303436
rect 397292 149548 397348 159292
rect 397404 155652 397460 310380
rect 397404 155586 397460 155596
rect 397516 157556 397572 313628
rect 397180 149492 397348 149548
rect 397180 3108 397236 149492
rect 397180 3042 397236 3052
rect 397516 2884 397572 157500
rect 397628 155540 397684 313740
rect 397628 155474 397684 155484
rect 397740 310324 397796 310334
rect 397740 152180 397796 310268
rect 397740 152114 397796 152124
rect 397852 157332 397908 317212
rect 397852 152068 397908 157276
rect 397964 317156 398020 317166
rect 397964 157444 398020 317100
rect 399532 317044 399588 317054
rect 397964 152292 398020 157388
rect 397964 152226 398020 152236
rect 398076 313572 398132 313582
rect 397852 152002 397908 152012
rect 398076 151060 398132 313516
rect 399420 313460 399476 313470
rect 398972 311780 399028 311790
rect 398860 306964 398916 306974
rect 398860 161308 398916 306908
rect 398748 161252 398916 161308
rect 398636 158450 398692 158462
rect 398636 158398 398638 158450
rect 398690 158398 398692 158450
rect 398636 156100 398692 158398
rect 398636 156034 398692 156044
rect 398748 157892 398804 161252
rect 398972 158452 399028 311724
rect 399308 310212 399364 310222
rect 399196 310100 399252 310110
rect 398076 126028 398132 151004
rect 398748 149548 398804 157836
rect 398860 158396 399028 158452
rect 399084 309988 399140 309998
rect 399084 158450 399140 309932
rect 399084 158398 399086 158450
rect 399138 158398 399140 158450
rect 398860 157668 398916 158396
rect 399084 158386 399140 158398
rect 399196 158452 399252 310044
rect 399196 158386 399252 158396
rect 398860 154980 398916 157612
rect 398972 158228 399028 158238
rect 399308 158228 399364 310156
rect 398972 155092 399028 158172
rect 399196 158172 399364 158228
rect 399420 158228 399476 313404
rect 398972 155036 399140 155092
rect 398860 154924 399028 154980
rect 398748 149492 398916 149548
rect 397516 2818 397572 2828
rect 397740 125972 398132 126028
rect 397740 2772 397796 125972
rect 397740 2706 397796 2716
rect 398860 1428 398916 149492
rect 398972 1540 399028 154924
rect 399084 154420 399140 155036
rect 399084 4004 399140 154364
rect 399196 154196 399252 158172
rect 399420 158162 399476 158172
rect 399532 158114 399588 316988
rect 399532 158062 399534 158114
rect 399586 158062 399588 158114
rect 399532 158050 399588 158062
rect 399644 316932 399700 316942
rect 399308 158002 399364 158014
rect 399308 157950 399310 158002
rect 399362 157950 399364 158002
rect 399308 157556 399364 157950
rect 399532 157890 399588 157902
rect 399532 157838 399534 157890
rect 399586 157838 399588 157890
rect 399308 157500 399476 157556
rect 399196 149548 399252 154140
rect 399420 155876 399476 157500
rect 399196 149492 399364 149548
rect 399308 6580 399364 149492
rect 399420 9828 399476 155820
rect 399420 9762 399476 9772
rect 399532 154308 399588 157838
rect 399308 6514 399364 6524
rect 399084 3938 399140 3948
rect 399532 2660 399588 154252
rect 399644 155988 399700 316876
rect 399756 316820 399812 316830
rect 399756 158002 399812 316764
rect 407708 315812 407764 320012
rect 410172 320012 410872 320068
rect 413980 320012 414680 320068
rect 418348 320012 418488 320068
rect 421708 320012 422296 320068
rect 425068 320012 426104 320068
rect 428428 320012 429912 320068
rect 433468 320012 433720 320068
rect 436828 320012 437528 320068
rect 440188 320012 441336 320068
rect 445256 320012 445396 320068
rect 410172 317268 410228 320012
rect 410172 317202 410228 317212
rect 413980 317156 414036 320012
rect 413980 317090 414036 317100
rect 407708 315746 407764 315756
rect 418348 313796 418404 320012
rect 418348 313730 418404 313740
rect 421708 313684 421764 320012
rect 421708 313618 421764 313628
rect 425068 313572 425124 320012
rect 425068 313506 425124 313516
rect 400316 313348 400372 313358
rect 400204 306852 400260 306862
rect 399756 157950 399758 158002
rect 399810 157950 399812 158002
rect 399756 157938 399812 157950
rect 399868 158228 399924 158238
rect 399756 157780 399812 157790
rect 399868 157780 399924 158172
rect 399812 157724 399924 157780
rect 399756 157220 399812 157724
rect 399756 157154 399812 157164
rect 399644 153860 399700 155932
rect 399644 153794 399700 153804
rect 400204 151172 400260 306796
rect 400316 154532 400372 313292
rect 428428 310436 428484 320012
rect 428428 310370 428484 310380
rect 433468 310324 433524 320012
rect 433468 310258 433524 310268
rect 436828 310212 436884 320012
rect 440188 311780 440244 320012
rect 445340 314188 445396 320012
rect 448588 320012 448952 320068
rect 452060 320012 452760 320068
rect 455980 320012 456568 320068
rect 460488 320012 460628 320068
rect 448588 317044 448644 320012
rect 448588 316978 448644 316988
rect 452060 316932 452116 320012
rect 452060 316866 452116 316876
rect 455980 316820 456036 320012
rect 455980 316754 456036 316764
rect 460572 314188 460628 320012
rect 445228 314132 445396 314188
rect 460348 314132 460628 314188
rect 463708 320012 464184 320068
rect 467068 320012 467992 320068
rect 470428 320012 471800 320068
rect 475468 320012 475608 320068
rect 478828 320012 479416 320068
rect 482188 320012 483224 320068
rect 485548 320012 487032 320068
rect 490588 320012 490840 320068
rect 493948 320012 494648 320068
rect 497308 320012 498456 320068
rect 502376 320012 502516 320068
rect 445228 313460 445284 314132
rect 445228 313394 445284 313404
rect 460348 313348 460404 314132
rect 460348 313282 460404 313292
rect 440188 311714 440244 311724
rect 436828 310146 436884 310156
rect 463708 310100 463764 320012
rect 463708 310034 463764 310044
rect 467068 309988 467124 320012
rect 467068 309922 467124 309932
rect 470428 306964 470484 320012
rect 470428 306898 470484 306908
rect 475468 306852 475524 320012
rect 475468 306786 475524 306796
rect 478828 303604 478884 320012
rect 482188 306740 482244 320012
rect 482188 306674 482244 306684
rect 478828 303538 478884 303548
rect 485548 303492 485604 320012
rect 485548 303426 485604 303436
rect 490588 303380 490644 320012
rect 490588 303314 490644 303324
rect 400316 154466 400372 154476
rect 400428 303268 400484 303278
rect 400204 151106 400260 151116
rect 400428 114268 400484 303212
rect 493948 303268 494004 320012
rect 497308 309988 497364 320012
rect 502460 314188 502516 320012
rect 502348 314132 502516 314188
rect 505708 320012 506072 320068
rect 509180 320012 509880 320068
rect 512428 320012 513688 320068
rect 517608 320012 517748 320068
rect 521416 320012 522116 320068
rect 525224 320012 525476 320068
rect 502348 313348 502404 314132
rect 502348 313282 502404 313292
rect 505708 310100 505764 320012
rect 509180 315028 509236 320012
rect 509180 314962 509236 314972
rect 505708 310034 505764 310044
rect 497308 309922 497364 309932
rect 493948 303202 494004 303212
rect 512428 303268 512484 320012
rect 517692 314188 517748 320012
rect 522060 316820 522116 320012
rect 525420 316932 525476 320012
rect 525420 316866 525476 316876
rect 527548 320012 528920 320068
rect 532588 320012 532728 320068
rect 536648 320012 537236 320068
rect 522060 316754 522116 316764
rect 517468 314132 517748 314188
rect 517468 310212 517524 314132
rect 527548 313460 527604 320012
rect 532588 313572 532644 320012
rect 537180 317044 537236 320012
rect 537180 316978 537236 316988
rect 539644 320012 540344 320068
rect 542668 320012 544152 320068
rect 547708 320012 547960 320068
rect 551880 320012 552580 320068
rect 539644 316708 539700 320012
rect 539644 316642 539700 316652
rect 542668 313684 542724 320012
rect 542668 313618 542724 313628
rect 532588 313506 532644 313516
rect 527548 313394 527604 313404
rect 517468 310146 517524 310156
rect 547708 303380 547764 320012
rect 552524 316708 552580 320012
rect 552524 316642 552580 316652
rect 554428 320012 555576 320068
rect 559496 320012 560196 320068
rect 547708 303314 547764 303324
rect 512428 303202 512484 303212
rect 554428 301700 554484 320012
rect 560140 317156 560196 320012
rect 560140 317090 560196 317100
rect 562828 320012 563192 320068
rect 566188 320012 567000 320068
rect 570920 320012 571172 320068
rect 574728 320012 574868 320068
rect 562828 313796 562884 320012
rect 562828 313730 562884 313740
rect 566188 308308 566244 320012
rect 571116 317268 571172 320012
rect 571116 317202 571172 317212
rect 574812 314188 574868 320012
rect 579740 317268 579796 317278
rect 578060 317044 578116 317054
rect 566188 308242 566244 308252
rect 574588 314132 574868 314188
rect 577948 316932 578004 316942
rect 574588 304948 574644 314132
rect 577948 305732 578004 316876
rect 577948 305666 578004 305676
rect 574588 304882 574644 304892
rect 554428 301634 554484 301644
rect 400652 154532 400708 154542
rect 400652 149380 400708 154476
rect 403228 149492 403284 160104
rect 407148 159572 407204 160104
rect 407148 159506 407204 159516
rect 410844 157332 410900 160104
rect 414652 157444 414708 160104
rect 414652 157378 414708 157388
rect 410844 157266 410900 157276
rect 418460 155540 418516 160104
rect 422268 157556 422324 160104
rect 422268 157490 422324 157500
rect 418460 155474 418516 155484
rect 426076 151060 426132 160104
rect 429884 155652 429940 160104
rect 429884 155586 429940 155596
rect 433692 152628 433748 160104
rect 437500 154196 437556 160104
rect 441308 157668 441364 160104
rect 445228 157780 445284 160104
rect 445228 157714 445284 157724
rect 441308 157602 441364 157612
rect 448924 155876 448980 160104
rect 452732 155988 452788 160104
rect 452732 155922 452788 155932
rect 448924 155810 448980 155820
rect 456540 154308 456596 160104
rect 456540 154242 456596 154252
rect 459452 154868 459508 154878
rect 437500 154130 437556 154140
rect 433692 152562 433748 152572
rect 426076 150994 426132 151004
rect 403228 149426 403284 149436
rect 400652 149314 400708 149324
rect 459452 149380 459508 154812
rect 460348 154868 460404 160104
rect 460348 154802 460404 154812
rect 464156 154420 464212 160104
rect 467964 155988 468020 160104
rect 471772 157892 471828 160104
rect 471772 157826 471828 157836
rect 467964 155922 468020 155932
rect 464156 154354 464212 154364
rect 475580 151172 475636 160104
rect 479388 159684 479444 160104
rect 479388 159618 479444 159628
rect 475580 151106 475636 151116
rect 481292 154868 481348 154878
rect 459452 149314 459508 149324
rect 400428 114212 400708 114268
rect 399532 2594 399588 2604
rect 400652 102452 400708 114212
rect 481292 104132 481348 154812
rect 483196 154868 483252 160104
rect 487004 159348 487060 160104
rect 490812 159460 490868 160104
rect 490812 159394 490868 159404
rect 487004 159282 487060 159292
rect 483196 154802 483252 154812
rect 493052 154868 493108 154878
rect 481292 104066 481348 104076
rect 398972 1474 399028 1484
rect 398860 1362 398916 1372
rect 400652 1316 400708 102396
rect 493052 102452 493108 154812
rect 494620 154868 494676 160104
rect 494620 154802 494676 154812
rect 493052 102386 493108 102396
rect 496412 151172 496468 151182
rect 496412 7364 496468 151116
rect 498428 151172 498484 160104
rect 502376 160076 503188 160132
rect 498428 151106 498484 151116
rect 503132 152628 503188 160076
rect 506044 157332 506100 160104
rect 509852 158900 509908 160104
rect 509852 158834 509908 158844
rect 513212 160076 513688 160132
rect 517608 160076 518308 160132
rect 513212 159460 513268 160076
rect 506044 153748 506100 157276
rect 506044 153682 506100 153692
rect 496412 7298 496468 7308
rect 503132 6692 503188 152572
rect 513212 9940 513268 159404
rect 518252 154420 518308 160076
rect 521276 156212 521332 160104
rect 521276 156146 521332 156156
rect 525196 156100 525252 160104
rect 525196 156034 525252 156044
rect 528332 160076 528920 160132
rect 528332 155988 528388 160076
rect 528332 155204 528388 155932
rect 528332 155138 528388 155148
rect 532700 157780 532756 160104
rect 517356 138628 517412 138638
rect 517356 101556 517412 138572
rect 513212 9874 513268 9884
rect 516572 100884 516628 100894
rect 516572 8484 516628 100828
rect 517356 100884 517412 101500
rect 517356 100818 517412 100828
rect 518252 10052 518308 154364
rect 519036 153748 519092 153758
rect 519036 84980 519092 153692
rect 532700 152852 532756 157724
rect 532700 152786 532756 152796
rect 535948 160076 536536 160132
rect 535948 138628 536004 160076
rect 540316 157108 540372 160104
rect 540316 157042 540372 157052
rect 544124 155876 544180 160104
rect 544124 150500 544180 155820
rect 547708 160076 547960 160132
rect 551068 160076 551768 160132
rect 547708 157668 547764 160076
rect 547708 154084 547764 157612
rect 551068 159348 551124 160076
rect 551068 156324 551124 159292
rect 551068 156258 551124 156268
rect 555548 157556 555604 160104
rect 555548 155428 555604 157500
rect 555548 155362 555604 155372
rect 559468 159236 559524 160104
rect 563304 160076 563668 160132
rect 547708 154018 547764 154028
rect 559468 152740 559524 159180
rect 563612 157444 563668 160076
rect 566972 158788 567028 160104
rect 566972 158722 567028 158732
rect 570780 157892 570836 160104
rect 570780 157826 570836 157836
rect 563612 156324 563668 157388
rect 563612 156258 563668 156268
rect 559468 152674 559524 152684
rect 544124 150434 544180 150444
rect 535948 138562 536004 138572
rect 519036 84914 519092 84924
rect 530908 60060 532504 60116
rect 556108 60060 557480 60116
rect 530908 12628 530964 60060
rect 530908 12562 530964 12572
rect 518252 9986 518308 9996
rect 516572 8418 516628 8428
rect 503132 6626 503188 6636
rect 556108 5908 556164 60060
rect 556108 5842 556164 5852
rect 567868 12628 567924 12638
rect 400652 1250 400708 1260
rect 397068 1026 397124 1036
rect 195468 476 195832 480
rect 195468 420 195524 476
rect 194908 364 195524 420
rect 195580 392 195832 476
rect 195608 -960 195832 392
rect 196728 -960 196952 480
rect 197820 392 198072 480
rect 198940 392 199192 480
rect 197848 -960 198072 392
rect 198968 -960 199192 392
rect 200088 -960 200312 480
rect 201180 392 201432 480
rect 202300 392 202552 480
rect 201208 -960 201432 392
rect 202328 -960 202552 392
rect 203448 -960 203672 480
rect 204540 392 204792 480
rect 205660 392 205912 480
rect 204568 -960 204792 392
rect 205688 -960 205912 392
rect 206808 -960 207032 480
rect 207900 392 208152 480
rect 207928 -960 208152 392
rect 209048 -960 209272 480
rect 210168 -960 210392 480
rect 211288 -960 211512 480
rect 212408 -960 212632 480
rect 213528 -960 213752 480
rect 214648 -960 214872 480
rect 215768 -960 215992 480
rect 216888 -960 217112 480
rect 218008 -960 218232 480
rect 219128 -960 219352 480
rect 220248 -960 220472 480
rect 221368 -960 221592 480
rect 222488 -960 222712 480
rect 223608 -960 223832 480
rect 224728 -960 224952 480
rect 225848 -960 226072 480
rect 226968 -960 227192 480
rect 228088 -960 228312 480
rect 229208 -960 229432 480
rect 230328 -960 230552 480
rect 231448 -960 231672 480
rect 232568 -960 232792 480
rect 233688 -960 233912 480
rect 234808 -960 235032 480
rect 235928 -960 236152 480
rect 237048 -960 237272 480
rect 238168 -960 238392 480
rect 239288 -960 239512 480
rect 240408 -960 240632 480
rect 241528 -960 241752 480
rect 242648 -960 242872 480
rect 243768 -960 243992 480
rect 244888 -960 245112 480
rect 246008 -960 246232 480
rect 247128 -960 247352 480
rect 248248 -960 248472 480
rect 249368 -960 249592 480
rect 250488 -960 250712 480
rect 251608 -960 251832 480
rect 252728 -960 252952 480
rect 253848 -960 254072 480
rect 254968 -960 255192 480
rect 256088 -960 256312 480
rect 257208 -960 257432 480
rect 258328 -960 258552 480
rect 259448 -960 259672 480
rect 260568 -960 260792 480
rect 261688 -960 261912 480
rect 262808 -960 263032 480
rect 263928 -960 264152 480
rect 265048 -960 265272 480
rect 266168 -960 266392 480
rect 267288 -960 267512 480
rect 268408 -960 268632 480
rect 269528 -960 269752 480
rect 270648 -960 270872 480
rect 271768 -960 271992 480
rect 272888 -960 273112 480
rect 274008 -960 274232 480
rect 275128 -960 275352 480
rect 276248 -960 276472 480
rect 277368 -960 277592 480
rect 278488 -960 278712 480
rect 279608 -960 279832 480
rect 280728 -960 280952 480
rect 281848 -960 282072 480
rect 282968 -960 283192 480
rect 284088 -960 284312 480
rect 285208 -960 285432 480
rect 286328 -960 286552 480
rect 287448 -960 287672 480
rect 288568 -960 288792 480
rect 289688 -960 289912 480
rect 290808 -960 291032 480
rect 291928 -960 292152 480
rect 293048 -960 293272 480
rect 294168 -960 294392 480
rect 295288 -960 295512 480
rect 296408 -960 296632 480
rect 297528 -960 297752 480
rect 298648 -960 298872 480
rect 299768 -960 299992 480
rect 300888 -960 301112 480
rect 302008 -960 302232 480
rect 303128 -960 303352 480
rect 304248 -960 304472 480
rect 305368 -960 305592 480
rect 306488 -960 306712 480
rect 307608 -960 307832 480
rect 308728 -960 308952 480
rect 309848 -960 310072 480
rect 310968 -960 311192 480
rect 312088 -960 312312 480
rect 313208 -960 313432 480
rect 314328 -960 314552 480
rect 315448 -960 315672 480
rect 316568 -960 316792 480
rect 317688 -960 317912 480
rect 318808 -960 319032 480
rect 319928 -960 320152 480
rect 321048 -960 321272 480
rect 322168 -960 322392 480
rect 323288 -960 323512 480
rect 324408 -960 324632 480
rect 325528 -960 325752 480
rect 326648 -960 326872 480
rect 327768 -960 327992 480
rect 328888 -960 329112 480
rect 330008 -960 330232 480
rect 331128 -960 331352 480
rect 332248 -960 332472 480
rect 333368 -960 333592 480
rect 334488 -960 334712 480
rect 335608 -960 335832 480
rect 336728 -960 336952 480
rect 337848 -960 338072 480
rect 338968 -960 339192 480
rect 340088 -960 340312 480
rect 341208 -960 341432 480
rect 342328 -960 342552 480
rect 343448 -960 343672 480
rect 344568 -960 344792 480
rect 345688 -960 345912 480
rect 346808 -960 347032 480
rect 347928 -960 348152 480
rect 349048 -960 349272 480
rect 350168 -960 350392 480
rect 351288 -960 351512 480
rect 352408 392 352660 480
rect 352408 -960 352632 392
rect 353528 -960 353752 480
rect 354648 -960 354872 480
rect 355768 -960 355992 480
rect 356888 -960 357112 480
rect 358008 -960 358232 480
rect 359128 -960 359352 480
rect 360248 -960 360472 480
rect 361368 -960 361592 480
rect 362488 -960 362712 480
rect 363608 -960 363832 480
rect 364728 -960 364952 480
rect 365848 -960 366072 480
rect 366968 -960 367192 480
rect 368088 -960 368312 480
rect 369208 -960 369432 480
rect 370328 -960 370552 480
rect 371448 -960 371672 480
rect 372568 -960 372792 480
rect 373688 -960 373912 480
rect 374808 -960 375032 480
rect 375928 -960 376152 480
rect 377048 -960 377272 480
rect 378168 -960 378392 480
rect 379288 -960 379512 480
rect 380408 -960 380632 480
rect 381528 -960 381752 480
rect 382648 -960 382872 480
rect 383768 -960 383992 480
rect 384888 -960 385112 480
rect 386008 -960 386232 480
rect 387128 -960 387352 480
rect 388248 -960 388472 480
rect 389368 -960 389592 480
rect 390488 -960 390712 480
rect 391608 -960 391832 480
rect 392728 -960 392952 480
rect 393848 -960 394072 480
rect 394968 -960 395192 480
rect 396088 -960 396312 480
rect 397208 -960 397432 480
rect 398328 -960 398552 480
rect 399448 -960 399672 480
rect 400568 -960 400792 480
rect 401688 -960 401912 480
rect 402808 -960 403032 480
rect 403928 -960 404152 480
rect 405048 -960 405272 480
rect 406168 -960 406392 480
rect 407288 -960 407512 480
rect 408408 -960 408632 480
rect 409528 -960 409752 480
rect 410648 -960 410872 480
rect 411768 -960 411992 480
rect 412888 -960 413112 480
rect 414008 -960 414232 480
rect 415128 -960 415352 480
rect 416248 -960 416472 480
rect 417368 -960 417592 480
rect 418488 -960 418712 480
rect 419608 -960 419832 480
rect 420728 -960 420952 480
rect 421848 -960 422072 480
rect 422968 -960 423192 480
rect 424088 -960 424312 480
rect 425208 -960 425432 480
rect 426328 -960 426552 480
rect 427448 -960 427672 480
rect 428568 -960 428792 480
rect 429688 -960 429912 480
rect 430808 -960 431032 480
rect 431928 -960 432152 480
rect 433048 -960 433272 480
rect 434168 -960 434392 480
rect 435288 -960 435512 480
rect 436408 -960 436632 480
rect 437528 -960 437752 480
rect 438648 -960 438872 480
rect 439768 -960 439992 480
rect 440888 -960 441112 480
rect 442008 -960 442232 480
rect 443128 -960 443352 480
rect 444248 -960 444472 480
rect 445368 -960 445592 480
rect 446488 -960 446712 480
rect 447608 -960 447832 480
rect 448728 -960 448952 480
rect 449848 -960 450072 480
rect 450968 -960 451192 480
rect 452088 -960 452312 480
rect 453208 -960 453432 480
rect 454328 -960 454552 480
rect 455448 -960 455672 480
rect 456568 -960 456792 480
rect 457688 -960 457912 480
rect 458808 -960 459032 480
rect 459928 -960 460152 480
rect 461048 -960 461272 480
rect 462168 -960 462392 480
rect 463288 -960 463512 480
rect 464408 -960 464632 480
rect 465528 -960 465752 480
rect 466648 -960 466872 480
rect 467768 -960 467992 480
rect 468888 -960 469112 480
rect 470008 -960 470232 480
rect 471128 -960 471352 480
rect 472248 -960 472472 480
rect 473368 -960 473592 480
rect 474488 -960 474712 480
rect 475608 -960 475832 480
rect 476728 -960 476952 480
rect 477848 -960 478072 480
rect 478968 -960 479192 480
rect 480088 -960 480312 480
rect 481208 -960 481432 480
rect 482328 -960 482552 480
rect 483448 -960 483672 480
rect 484568 -960 484792 480
rect 485688 -960 485912 480
rect 486808 -960 487032 480
rect 487928 -960 488152 480
rect 489048 -960 489272 480
rect 490168 -960 490392 480
rect 491288 -960 491512 480
rect 492408 -960 492632 480
rect 493528 -960 493752 480
rect 494648 -960 494872 480
rect 495768 -960 495992 480
rect 496888 -960 497112 480
rect 498008 -960 498232 480
rect 499128 -960 499352 480
rect 500248 -960 500472 480
rect 501368 -960 501592 480
rect 502488 -960 502712 480
rect 503608 -960 503832 480
rect 504728 -960 504952 480
rect 505848 -960 506072 480
rect 506968 -960 507192 480
rect 508088 -960 508312 480
rect 509208 -960 509432 480
rect 510328 -960 510552 480
rect 511448 -960 511672 480
rect 512568 -960 512792 480
rect 513688 -960 513912 480
rect 514808 -960 515032 480
rect 515928 -960 516152 480
rect 517048 -960 517272 480
rect 518168 -960 518392 480
rect 519288 -960 519512 480
rect 520408 -960 520632 480
rect 521528 -960 521752 480
rect 522648 -960 522872 480
rect 523768 -960 523992 480
rect 524888 -960 525112 480
rect 526008 -960 526232 480
rect 527128 -960 527352 480
rect 528248 -960 528472 480
rect 529368 -960 529592 480
rect 530488 -960 530712 480
rect 531608 -960 531832 480
rect 532728 -960 532952 480
rect 533848 -960 534072 480
rect 534968 -960 535192 480
rect 536088 -960 536312 480
rect 537208 -960 537432 480
rect 538328 -960 538552 480
rect 539448 -960 539672 480
rect 540568 -960 540792 480
rect 541688 -960 541912 480
rect 542808 -960 543032 480
rect 543928 -960 544152 480
rect 545048 -960 545272 480
rect 546168 -960 546392 480
rect 547288 -960 547512 480
rect 548408 -960 548632 480
rect 549528 -960 549752 480
rect 550648 -960 550872 480
rect 551768 -960 551992 480
rect 552888 -960 553112 480
rect 554008 -960 554232 480
rect 555128 -960 555352 480
rect 556248 -960 556472 480
rect 557368 -960 557592 480
rect 558488 -960 558712 480
rect 559608 -960 559832 480
rect 560728 -960 560952 480
rect 561848 -960 562072 480
rect 562968 -960 563192 480
rect 564088 -960 564312 480
rect 565208 -960 565432 480
rect 566328 -960 566552 480
rect 567448 -960 567672 480
rect 567868 420 567924 12572
rect 574588 2548 574644 160104
rect 578060 153748 578116 316988
rect 578284 316820 578340 316830
rect 578060 153682 578116 153692
rect 578172 313348 578228 313358
rect 578172 152628 578228 313292
rect 578284 156212 578340 316764
rect 578508 313684 578564 313694
rect 578284 156146 578340 156156
rect 578396 313460 578452 313470
rect 578396 155988 578452 313404
rect 578396 155922 578452 155932
rect 578508 155876 578564 313628
rect 579628 309988 579684 309998
rect 578620 305732 578676 305742
rect 578620 304164 578676 305676
rect 578620 156100 578676 304108
rect 578732 301700 578788 301710
rect 578732 157556 578788 301644
rect 578732 157490 578788 157500
rect 578620 156034 578676 156044
rect 578508 155810 578564 155820
rect 578172 152562 578228 152572
rect 579628 151172 579684 309932
rect 579740 157892 579796 317212
rect 581420 317156 581476 317166
rect 581308 316708 581364 316718
rect 579964 313572 580020 313582
rect 579740 157826 579796 157836
rect 579852 310212 579908 310222
rect 579852 154420 579908 310156
rect 579964 157780 580020 313516
rect 579964 157714 580020 157724
rect 580076 310100 580132 310110
rect 580076 157332 580132 310044
rect 580188 303380 580244 303390
rect 580188 157668 580244 303324
rect 580300 303268 580356 303278
rect 580300 159460 580356 303212
rect 580300 159394 580356 159404
rect 581308 159348 581364 316652
rect 581308 159282 581364 159292
rect 581420 159236 581476 317100
rect 581420 159170 581476 159180
rect 584668 313796 584724 313806
rect 580188 157602 580244 157612
rect 584668 157444 584724 313740
rect 587132 301588 587188 451052
rect 587244 406756 587300 406766
rect 587244 306628 587300 406700
rect 589708 395668 589764 395678
rect 587356 362404 587412 362414
rect 587356 311668 587412 362348
rect 587356 311602 587412 311612
rect 587244 306562 587300 306572
rect 587132 301522 587188 301532
rect 584668 157378 584724 157388
rect 580076 157266 580132 157276
rect 579852 154354 579908 154364
rect 579628 151106 579684 151116
rect 589708 149492 589764 395612
rect 589820 319172 589876 484316
rect 590044 440020 590100 440030
rect 589820 319106 589876 319116
rect 589932 351316 589988 351326
rect 589708 149426 589764 149436
rect 589820 295876 589876 295886
rect 589820 84084 589876 295820
rect 589932 159572 589988 351260
rect 590044 315812 590100 439964
rect 590044 315746 590100 315756
rect 589932 159506 589988 159516
rect 589820 84018 589876 84028
rect 574588 2482 574644 2492
rect 568428 480 568596 532
rect 568428 476 568792 480
rect 568428 420 568484 476
rect 567868 364 568484 420
rect 568540 392 568792 476
rect 568568 -960 568792 392
rect 569688 -960 569912 480
rect 570808 -960 571032 480
rect 571928 -960 572152 480
<< via2 >>
rect 9884 587916 9940 587972
rect 3276 587356 3332 587412
rect 3164 320908 3220 320964
rect 2492 268828 2548 268884
rect 28 225148 84 225204
rect 28 47068 84 47124
rect 2604 181804 2660 181860
rect 26012 587356 26068 587412
rect 8316 587244 8372 587300
rect 7532 507724 7588 507780
rect 5852 475132 5908 475188
rect 3388 431788 3444 431844
rect 3388 321020 3444 321076
rect 4172 420812 4228 420868
rect 3276 319228 3332 319284
rect 3164 157276 3220 157332
rect 2604 35308 2660 35364
rect 3276 75628 3332 75684
rect 2492 21868 2548 21924
rect 3276 19404 3332 19460
rect 4172 12796 4228 12852
rect 4284 388220 4340 388276
rect 4396 377356 4452 377412
rect 4396 70812 4452 70868
rect 4508 344764 4564 344820
rect 4732 333900 4788 333956
rect 4620 290444 4676 290500
rect 4844 301308 4900 301364
rect 6636 316652 6692 316708
rect 6524 310044 6580 310100
rect 6412 303212 6468 303268
rect 6300 301532 6356 301588
rect 5852 159628 5908 159684
rect 6076 160076 6132 160132
rect 4844 70700 4900 70756
rect 4956 78988 5012 79044
rect 4732 68908 4788 68964
rect 6300 157612 6356 157668
rect 6524 159516 6580 159572
rect 6412 155372 6468 155428
rect 7420 301756 7476 301812
rect 7420 157724 7476 157780
rect 6636 148652 6692 148708
rect 6076 40460 6132 40516
rect 6524 73948 6580 74004
rect 4956 21420 5012 21476
rect 6524 21308 6580 21364
rect 6636 72380 6692 72436
rect 6636 19964 6692 20020
rect 7868 464268 7924 464324
rect 7644 313516 7700 313572
rect 7644 159404 7700 159460
rect 7756 310156 7812 310212
rect 7756 152796 7812 152852
rect 7532 19740 7588 19796
rect 4620 17948 4676 18004
rect 8204 317100 8260 317156
rect 8092 316988 8148 317044
rect 7980 316876 8036 316932
rect 7980 157388 8036 157444
rect 8092 156940 8148 156996
rect 8204 154140 8260 154196
rect 75068 587244 75124 587300
rect 9996 587132 10052 587188
rect 91420 587132 91476 587188
rect 205884 587468 205940 587524
rect 196476 587356 196532 587412
rect 157052 587244 157108 587300
rect 188972 587244 189028 587300
rect 140700 587132 140756 587188
rect 13244 319228 13300 319284
rect 9996 319116 10052 319172
rect 17052 319116 17108 319172
rect 9660 317324 9716 317380
rect 9548 309932 9604 309988
rect 9436 303436 9492 303492
rect 9100 301644 9156 301700
rect 9100 157836 9156 157892
rect 9212 246988 9268 247044
rect 9324 203532 9380 203588
rect 9772 317212 9828 317268
rect 9996 313740 10052 313796
rect 9772 159292 9828 159348
rect 9884 313628 9940 313684
rect 9660 159180 9716 159236
rect 9548 158732 9604 158788
rect 9436 157500 9492 157556
rect 9884 154364 9940 154420
rect 10444 313292 10500 313348
rect 20188 301756 20244 301812
rect 32284 317324 32340 317380
rect 26908 303436 26964 303492
rect 23548 301644 23604 301700
rect 39900 317212 39956 317268
rect 43708 317100 43764 317156
rect 47068 313740 47124 313796
rect 50428 313628 50484 313684
rect 58940 316988 58996 317044
rect 62748 316876 62804 316932
rect 53788 313516 53844 313572
rect 65548 313404 65604 313460
rect 68908 313292 68964 313348
rect 73948 310156 74004 310212
rect 77308 310044 77364 310100
rect 85596 316764 85652 316820
rect 89404 316652 89460 316708
rect 80668 303324 80724 303380
rect 97020 316652 97076 316708
rect 112252 316764 112308 316820
rect 115948 313292 116004 313348
rect 119308 309932 119364 309988
rect 122668 307020 122724 307076
rect 107548 306908 107604 306964
rect 104188 306796 104244 306852
rect 100828 306684 100884 306740
rect 92428 303212 92484 303268
rect 131292 316876 131348 316932
rect 150332 317100 150388 317156
rect 146524 316988 146580 317044
rect 161308 313628 161364 313684
rect 157948 313516 158004 313572
rect 152908 313404 152964 313460
rect 164668 309932 164724 309988
rect 176988 317212 177044 317268
rect 173068 311724 173124 311780
rect 168028 308252 168084 308308
rect 141148 303548 141204 303604
rect 137788 303436 137844 303492
rect 134428 303324 134484 303380
rect 126028 303212 126084 303268
rect 188972 319228 189028 319284
rect 189868 587132 189924 587188
rect 184604 317324 184660 317380
rect 188300 317212 188356 317268
rect 188188 317100 188244 317156
rect 179788 301980 179844 302036
rect 188076 316764 188132 316820
rect 35308 301532 35364 301588
rect 188076 160188 188132 160244
rect 17052 159628 17108 159684
rect 24668 157836 24724 157892
rect 20860 157724 20916 157780
rect 22652 157724 22708 157780
rect 13244 157276 13300 157332
rect 10444 156156 10500 156212
rect 9996 154252 10052 154308
rect 21868 145292 21924 145348
rect 11788 126028 11844 126084
rect 10892 116620 10948 116676
rect 9324 54796 9380 54852
rect 9996 74396 10052 74452
rect 9212 30156 9268 30212
rect 10108 69020 10164 69076
rect 11676 77308 11732 77364
rect 10892 66892 10948 66948
rect 11564 70588 11620 70644
rect 10108 62524 10164 62580
rect 9996 21196 10052 21252
rect 10892 40572 10948 40628
rect 8316 21084 8372 21140
rect 7868 16492 7924 16548
rect 11004 29708 11060 29764
rect 11564 20188 11620 20244
rect 11004 20076 11060 20132
rect 32284 159180 32340 159236
rect 33292 159180 33348 159236
rect 28476 157500 28532 157556
rect 28476 157164 28532 157220
rect 31948 158844 32004 158900
rect 24668 156268 24724 156324
rect 27692 156268 27748 156324
rect 22652 120092 22708 120148
rect 26908 138572 26964 138628
rect 25564 119308 25620 119364
rect 24220 119196 24276 119252
rect 27692 135212 27748 135268
rect 29372 143612 29428 143668
rect 27468 129388 27524 129444
rect 28812 127708 28868 127764
rect 29372 119196 29428 119252
rect 30940 120988 30996 121044
rect 33292 156380 33348 156436
rect 36092 157612 36148 157668
rect 39900 159292 39956 159348
rect 39900 157052 39956 157108
rect 41132 156380 41188 156436
rect 36092 156268 36148 156324
rect 37772 156268 37828 156324
rect 36988 133532 37044 133588
rect 34188 126028 34244 126084
rect 33628 121100 33684 121156
rect 36876 115948 36932 116004
rect 37772 132636 37828 132692
rect 46172 157164 46228 157220
rect 43708 154140 43764 154196
rect 44492 154140 44548 154196
rect 41132 122556 41188 122612
rect 43820 150332 43876 150388
rect 41692 119196 41748 119252
rect 40348 118412 40404 118468
rect 39004 118076 39060 118132
rect 43036 118636 43092 118692
rect 44492 129276 44548 129332
rect 45388 148764 45444 148820
rect 43820 118076 43876 118132
rect 44380 123564 44436 123620
rect 48748 155596 48804 155652
rect 47516 154252 47572 154308
rect 47852 154252 47908 154308
rect 46172 127596 46228 127652
rect 47068 137788 47124 137844
rect 47852 136892 47908 136948
rect 47068 120652 47124 120708
rect 47180 126924 47236 126980
rect 45388 119196 45444 119252
rect 47740 120652 47796 120708
rect 45724 118524 45780 118580
rect 55132 159404 55188 159460
rect 56364 159404 56420 159460
rect 55468 158732 55524 158788
rect 51212 154364 51268 154420
rect 50428 140252 50484 140308
rect 48748 118636 48804 118692
rect 49756 118972 49812 119028
rect 51212 124236 51268 124292
rect 52892 155484 52948 155540
rect 53788 150556 53844 150612
rect 56364 157164 56420 157220
rect 59724 156940 59780 156996
rect 59612 143836 59668 143892
rect 52892 118972 52948 119028
rect 53788 118636 53844 118692
rect 52444 117628 52500 117684
rect 57820 121772 57876 121828
rect 62300 158956 62356 159012
rect 63084 157388 63140 157444
rect 62972 152012 63028 152068
rect 59724 131852 59780 131908
rect 59612 118636 59668 118692
rect 66332 154476 66388 154532
rect 63084 128492 63140 128548
rect 63868 148652 63924 148708
rect 62972 118524 63028 118580
rect 65548 146972 65604 147028
rect 69692 156156 69748 156212
rect 68908 145404 68964 145460
rect 67228 141932 67284 141988
rect 66332 133644 66388 133700
rect 65548 118412 65604 118468
rect 67228 119196 67284 119252
rect 66556 116060 66612 116116
rect 70364 156156 70420 156212
rect 71372 157052 71428 157108
rect 69692 130956 69748 131012
rect 70588 142044 70644 142100
rect 77980 159516 78036 159572
rect 78876 159516 78932 159572
rect 78876 157052 78932 157108
rect 81788 159068 81844 159124
rect 74172 156380 74228 156436
rect 74172 152796 74228 152852
rect 78988 150444 79044 150500
rect 71372 135996 71428 136052
rect 73052 146972 73108 147028
rect 75628 145516 75684 145572
rect 77308 138684 77364 138740
rect 73052 119196 73108 119252
rect 84812 156044 84868 156100
rect 81788 150332 81844 150388
rect 82348 155372 82404 155428
rect 84028 153244 84084 153300
rect 80668 118412 80724 118468
rect 82012 116172 82068 116228
rect 84812 147084 84868 147140
rect 86492 157164 86548 157220
rect 85708 126140 85764 126196
rect 86716 157052 86772 157108
rect 93212 159180 93268 159236
rect 89068 149548 89124 149604
rect 89068 148764 89124 148820
rect 90636 157052 90692 157108
rect 87388 143724 87444 143780
rect 86716 130172 86772 130228
rect 86492 120316 86548 120372
rect 87388 118300 87444 118356
rect 89068 125916 89124 125972
rect 90636 125916 90692 125972
rect 91532 156268 91588 156324
rect 89068 123564 89124 123620
rect 90076 125244 90132 125300
rect 89180 123452 89236 123508
rect 89180 118300 89236 118356
rect 91420 125132 91476 125188
rect 97020 157052 97076 157108
rect 97468 159964 97524 160020
rect 93212 155596 93268 155652
rect 96012 131068 96068 131124
rect 91532 123564 91588 123620
rect 94108 126812 94164 126868
rect 92764 120204 92820 120260
rect 95452 117852 95508 117908
rect 100940 154476 100996 154532
rect 99148 153692 99204 153748
rect 100828 152236 100884 152292
rect 100940 152012 100996 152068
rect 100828 120652 100884 120708
rect 101052 131180 101108 131236
rect 107436 153804 107492 153860
rect 107324 139356 107380 139412
rect 104188 129164 104244 129220
rect 104972 139020 105028 139076
rect 104860 122668 104916 122724
rect 101500 120652 101556 120708
rect 103516 119196 103572 119252
rect 107324 137788 107380 137844
rect 105532 129164 105588 129220
rect 105532 126924 105588 126980
rect 107436 124124 107492 124180
rect 107436 122668 107492 122724
rect 107548 147084 107604 147140
rect 107324 121884 107380 121940
rect 104972 119196 105028 119252
rect 106204 119084 106260 119140
rect 112252 159516 112308 159572
rect 116732 156940 116788 156996
rect 112252 155484 112308 155540
rect 114268 155484 114324 155540
rect 110012 153916 110068 153972
rect 107660 139356 107716 139412
rect 109228 148092 109284 148148
rect 107660 138908 107716 138964
rect 110012 119084 110068 119140
rect 110908 152012 110964 152068
rect 112588 142156 112644 142212
rect 116732 140252 116788 140308
rect 117628 155596 117684 155652
rect 116956 119420 117012 119476
rect 115612 117740 115668 117796
rect 119308 152124 119364 152180
rect 123676 159740 123732 159796
rect 131292 154364 131348 154420
rect 131292 153916 131348 153972
rect 127484 153804 127540 153860
rect 127708 153804 127764 153860
rect 119420 143836 119476 143892
rect 126028 152348 126084 152404
rect 122668 139020 122724 139076
rect 122668 138796 122724 138852
rect 120988 126252 121044 126308
rect 122332 124348 122388 124404
rect 125020 122668 125076 122724
rect 134428 149436 134484 149492
rect 136892 147980 136948 148036
rect 134428 147084 134484 147140
rect 135212 147868 135268 147924
rect 127708 117964 127764 118020
rect 131068 137004 131124 137060
rect 130396 116284 130452 116340
rect 135212 127596 135268 127652
rect 135324 135212 135380 135268
rect 133084 120092 133140 120148
rect 133084 119084 133140 119140
rect 134428 119196 134484 119252
rect 135324 119196 135380 119252
rect 137004 146188 137060 146244
rect 140252 149660 140308 149716
rect 137788 139356 137844 139412
rect 138572 142828 138628 142884
rect 136892 119084 136948 119140
rect 137116 122556 137172 122612
rect 137788 132636 137844 132692
rect 138572 132636 138628 132692
rect 139468 135996 139524 136052
rect 141036 148092 141092 148148
rect 146188 147756 146244 147812
rect 149548 146972 149604 147028
rect 153692 157612 153748 157668
rect 148652 146412 148708 146468
rect 141036 137676 141092 137732
rect 142044 146300 142100 146356
rect 140252 135996 140308 136052
rect 141932 136892 141988 136948
rect 141932 136444 141988 136500
rect 141148 129276 141204 129332
rect 143724 144508 143780 144564
rect 143612 142940 143668 142996
rect 143612 136444 143668 136500
rect 142044 129276 142100 129332
rect 143836 124236 143892 124292
rect 145292 131852 145348 131908
rect 147868 128492 147924 128548
rect 145292 122780 145348 122836
rect 146524 122780 146580 122836
rect 145180 120316 145236 120372
rect 145180 119532 145236 119588
rect 147868 121212 147924 121268
rect 150332 144620 150388 144676
rect 148652 119196 148708 119252
rect 148876 133644 148932 133700
rect 148876 119196 148932 119252
rect 149772 130956 149828 131012
rect 150332 130956 150388 131012
rect 151900 123564 151956 123620
rect 158732 156828 158788 156884
rect 156268 150332 156324 150388
rect 157948 148764 158004 148820
rect 153692 123452 153748 123508
rect 153804 130172 153860 130228
rect 153804 124460 153860 124516
rect 151900 119644 151956 119700
rect 155932 123452 155988 123508
rect 154588 118076 154644 118132
rect 162092 157500 162148 157556
rect 158732 143724 158788 143780
rect 160412 152460 160468 152516
rect 159628 140252 159684 140308
rect 165564 157388 165620 157444
rect 162092 125244 162148 125300
rect 163772 156268 163828 156324
rect 165564 156268 165620 156324
rect 166348 158732 166404 158788
rect 163772 125132 163828 125188
rect 160412 119196 160468 119252
rect 165340 118524 165396 118580
rect 169372 157836 169428 157892
rect 167132 156268 167188 156324
rect 169372 156268 169428 156324
rect 173852 157276 173908 157332
rect 168028 153916 168084 153972
rect 169708 148876 169764 148932
rect 167132 120204 167188 120260
rect 168028 116396 168084 116452
rect 171388 128492 171444 128548
rect 173852 126812 173908 126868
rect 175532 156268 175588 156324
rect 176988 156268 177044 156324
rect 180572 157164 180628 157220
rect 188076 159516 188132 159572
rect 184604 153916 184660 153972
rect 188972 316988 189028 317044
rect 188748 311724 188804 311780
rect 188300 148764 188356 148820
rect 188412 303548 188468 303604
rect 188412 302540 188468 302596
rect 188188 145404 188244 145460
rect 180572 143612 180628 143668
rect 188524 303436 188580 303492
rect 188524 302428 188580 302484
rect 188636 303324 188692 303380
rect 188860 308364 188916 308420
rect 188860 157836 188916 157892
rect 188748 157276 188804 157332
rect 188972 157724 189028 157780
rect 188636 149436 188692 149492
rect 189644 316876 189700 316932
rect 189644 161308 189700 161364
rect 189644 154364 189700 154420
rect 188972 147756 189028 147812
rect 188524 139356 188580 139412
rect 188412 137676 188468 137732
rect 175532 123452 175588 123508
rect 188972 129388 189028 129444
rect 178780 118748 178836 118804
rect 173404 118636 173460 118692
rect 176876 117852 176932 117908
rect 176876 116732 176932 116788
rect 19292 113036 19348 113092
rect 19180 88844 19236 88900
rect 18172 71372 18228 71428
rect 18172 70588 18228 70644
rect 20076 111692 20132 111748
rect 19964 110348 20020 110404
rect 19852 109004 19908 109060
rect 19516 99596 19572 99652
rect 19292 70700 19348 70756
rect 19404 94108 19460 94164
rect 19180 69916 19236 69972
rect 19740 98252 19796 98308
rect 19628 96908 19684 96964
rect 19628 73612 19684 73668
rect 19516 70924 19572 70980
rect 19964 73500 20020 73556
rect 20076 73388 20132 73444
rect 20188 106316 20244 106372
rect 19852 72492 19908 72548
rect 20412 104972 20468 105028
rect 20188 70140 20244 70196
rect 20300 103628 20356 103684
rect 19740 69692 19796 69748
rect 19404 69132 19460 69188
rect 20412 70028 20468 70084
rect 21868 72268 21924 72324
rect 47404 70700 47460 70756
rect 21868 69356 21924 69412
rect 21980 70476 22036 70532
rect 64092 70140 64148 70196
rect 21980 68796 22036 68852
rect 20300 68572 20356 68628
rect 25564 68348 25620 68404
rect 33292 69356 33348 69412
rect 30940 69132 30996 69188
rect 31164 69132 31220 69188
rect 35644 69020 35700 69076
rect 31164 68796 31220 68852
rect 40348 69132 40404 69188
rect 37324 68572 37380 68628
rect 45052 68908 45108 68964
rect 42028 68572 42084 68628
rect 49084 68572 49140 68628
rect 52108 68572 52164 68628
rect 53788 68572 53844 68628
rect 56140 68572 56196 68628
rect 58828 68460 58884 68516
rect 60844 68460 60900 68516
rect 28588 68348 28644 68404
rect 63868 67116 63924 67172
rect 63980 69692 64036 69748
rect 11788 60508 11844 60564
rect 61516 66108 61572 66164
rect 61516 64652 61572 64708
rect 64540 70028 64596 70084
rect 64092 59500 64148 59556
rect 64204 69804 64260 69860
rect 63980 50764 64036 50820
rect 61516 44268 61572 44324
rect 64316 68572 64372 68628
rect 64876 69916 64932 69972
rect 64764 63868 64820 63924
rect 64428 58044 64484 58100
rect 64652 62412 64708 62468
rect 64316 56588 64372 56644
rect 64204 43484 64260 43540
rect 64316 52220 64372 52276
rect 63868 42028 63924 42084
rect 62188 39116 62244 39172
rect 61516 36988 61572 37044
rect 11676 19852 11732 19908
rect 14924 18508 14980 18564
rect 20412 17500 20468 17556
rect 23436 17500 23492 17556
rect 10892 16156 10948 16212
rect 23436 15036 23492 15092
rect 4508 8316 4564 8372
rect 4284 8204 4340 8260
rect 30268 5852 30324 5908
rect 42364 16828 42420 16884
rect 44716 16828 44772 16884
rect 44716 13356 44772 13412
rect 53340 17612 53396 17668
rect 60620 19516 60676 19572
rect 61964 27186 62020 27188
rect 61964 27134 61966 27186
rect 61966 27134 62018 27186
rect 62018 27134 62020 27186
rect 61964 27132 62020 27134
rect 60844 20972 60900 21028
rect 61516 22428 61572 22484
rect 61516 19964 61572 20020
rect 60732 14812 60788 14868
rect 60508 14588 60564 14644
rect 60396 12908 60452 12964
rect 58828 12572 58884 12628
rect 47852 10892 47908 10948
rect 62300 31836 62356 31892
rect 63980 26012 64036 26068
rect 63980 21196 64036 21252
rect 63868 16380 63924 16436
rect 62300 16268 62356 16324
rect 64540 49308 64596 49364
rect 64428 47852 64484 47908
rect 64540 18172 64596 18228
rect 64428 16604 64484 16660
rect 64316 13244 64372 13300
rect 66220 68908 66276 68964
rect 68572 68796 68628 68852
rect 77980 69132 78036 69188
rect 75628 69020 75684 69076
rect 80332 68684 80388 68740
rect 73276 67004 73332 67060
rect 70924 65436 70980 65492
rect 89740 68572 89796 68628
rect 87388 66892 87444 66948
rect 85036 66780 85092 66836
rect 82684 63756 82740 63812
rect 65100 60956 65156 61012
rect 64876 40572 64932 40628
rect 64988 55132 65044 55188
rect 64988 14924 65044 14980
rect 64764 14476 64820 14532
rect 90748 14364 90804 14420
rect 65100 13132 65156 13188
rect 64652 13020 64708 13076
rect 62188 9996 62244 10052
rect 96796 65548 96852 65604
rect 98252 65548 98308 65604
rect 94108 6076 94164 6132
rect 100828 24332 100884 24388
rect 102508 22652 102564 22708
rect 99148 21084 99204 21140
rect 110908 65548 110964 65604
rect 113260 62972 113316 63028
rect 113372 65548 113428 65604
rect 107548 27692 107604 27748
rect 105868 7644 105924 7700
rect 98252 4508 98308 4564
rect 115612 65548 115668 65604
rect 116732 65548 116788 65604
rect 116732 9324 116788 9380
rect 119308 20972 119364 21028
rect 117628 7532 117684 7588
rect 124348 11004 124404 11060
rect 129724 61292 129780 61348
rect 131068 15036 131124 15092
rect 131628 15036 131684 15092
rect 131628 14252 131684 14308
rect 126028 9212 126084 9268
rect 136108 7980 136164 8036
rect 134428 7868 134484 7924
rect 122668 5964 122724 6020
rect 134428 7644 134484 7700
rect 140028 14364 140084 14420
rect 137788 7420 137844 7476
rect 138460 7868 138516 7924
rect 134428 4620 134484 4676
rect 113372 4396 113428 4452
rect 35308 4284 35364 4340
rect 25228 4172 25284 4228
rect 146188 65884 146244 65940
rect 147980 65884 148036 65940
rect 147980 64652 148036 64708
rect 147868 22876 147924 22932
rect 142828 8428 142884 8484
rect 145292 22652 145348 22708
rect 141148 6748 141204 6804
rect 141820 7980 141876 8036
rect 145180 7420 145236 7476
rect 144060 6076 144116 6132
rect 148652 21084 148708 21140
rect 145292 4732 145348 4788
rect 148540 6748 148596 6804
rect 147420 4508 147476 4564
rect 152908 26796 152964 26852
rect 154588 64652 154644 64708
rect 152908 24332 152964 24388
rect 149548 14588 149604 14644
rect 151900 8428 151956 8484
rect 148652 4956 148708 5012
rect 150780 4956 150836 5012
rect 155596 64652 155652 64708
rect 157052 27692 157108 27748
rect 157948 22652 158004 22708
rect 158060 22876 158116 22932
rect 157052 4844 157108 4900
rect 157500 4732 157556 4788
rect 162652 65548 162708 65604
rect 163772 65548 163828 65604
rect 162092 62972 162148 63028
rect 159628 12796 159684 12852
rect 160412 14588 160468 14644
rect 160412 4956 160468 5012
rect 161980 4956 162036 5012
rect 160860 4620 160916 4676
rect 165004 64764 165060 64820
rect 163772 26012 163828 26068
rect 163996 26796 164052 26852
rect 162092 4732 162148 4788
rect 171500 64652 171556 64708
rect 169708 11116 169764 11172
rect 171388 22652 171444 22708
rect 166348 7644 166404 7700
rect 170268 11004 170324 11060
rect 163996 4396 164052 4452
rect 164220 4844 164276 4900
rect 167580 4508 167636 4564
rect 165340 4396 165396 4452
rect 170268 4396 170324 4452
rect 170940 4732 170996 4788
rect 168924 4060 168980 4116
rect 172060 62972 172116 63028
rect 175532 18508 175588 18564
rect 173068 13356 173124 13412
rect 174636 13356 174692 13412
rect 174636 12684 174692 12740
rect 174748 12796 174804 12852
rect 171500 4060 171556 4116
rect 174300 9324 174356 9380
rect 177212 9660 177268 9716
rect 178108 26012 178164 26068
rect 177660 7532 177716 7588
rect 179788 20972 179844 21028
rect 180572 64764 180628 64820
rect 188860 11116 188916 11172
rect 182364 7644 182420 7700
rect 180572 4060 180628 4116
rect 181468 5964 181524 6020
rect 181468 3500 181524 3556
rect 182140 4060 182196 4116
rect 180460 2492 180516 2548
rect 187740 4396 187796 4452
rect 182364 4060 182420 4116
rect 185500 4060 185556 4116
rect 184380 3500 184436 3556
rect 188972 10220 189028 10276
rect 189308 117964 189364 118020
rect 192332 582988 192388 583044
rect 191548 317324 191604 317380
rect 191212 313628 191268 313684
rect 190988 313516 191044 313572
rect 190652 313404 190708 313460
rect 189980 313292 190036 313348
rect 189980 157836 190036 157892
rect 190092 301980 190148 302036
rect 190652 158060 190708 158116
rect 190652 157612 190708 157668
rect 190764 309932 190820 309988
rect 190764 305004 190820 305060
rect 190764 157388 190820 157444
rect 190876 303212 190932 303268
rect 190876 158172 190932 158228
rect 190092 157164 190148 157220
rect 189980 156940 190036 156996
rect 189868 67116 189924 67172
rect 190652 124348 190708 124404
rect 189308 5740 189364 5796
rect 190988 301868 191044 301924
rect 191212 301644 191268 301700
rect 191436 307020 191492 307076
rect 191436 301756 191492 301812
rect 191436 159740 191492 159796
rect 191212 157500 191268 157556
rect 190988 156828 191044 156884
rect 190876 124124 190932 124180
rect 191436 151116 191492 151172
rect 191436 149548 191492 149604
rect 191324 121212 191380 121268
rect 190764 61292 190820 61348
rect 190764 4060 190820 4116
rect 191100 9212 191156 9268
rect 190652 2940 190708 2996
rect 191324 3052 191380 3108
rect 191548 128492 191604 128548
rect 191660 306908 191716 306964
rect 191884 306684 191940 306740
rect 191884 305788 191940 305844
rect 191884 154252 191940 154308
rect 191660 121884 191716 121940
rect 191660 121212 191716 121268
rect 194012 561148 194068 561204
rect 192332 69020 192388 69076
rect 192444 461132 192500 461188
rect 192556 317548 192612 317604
rect 193116 306796 193172 306852
rect 193116 305116 193172 305172
rect 193900 304108 193956 304164
rect 192668 302092 192724 302148
rect 194124 517468 194180 517524
rect 222236 587356 222292 587412
rect 402108 587244 402164 587300
rect 467516 587132 467572 587188
rect 532588 461132 532644 461188
rect 589820 484316 589876 484372
rect 587132 451052 587188 451108
rect 202300 319228 202356 319284
rect 196476 319116 196532 319172
rect 206108 319116 206164 319172
rect 194684 316988 194740 317044
rect 194124 159516 194180 159572
rect 194236 311612 194292 311668
rect 194012 156156 194068 156212
rect 193900 153692 193956 153748
rect 193228 152908 193284 152964
rect 193228 152236 193284 152292
rect 192668 151116 192724 151172
rect 194012 127708 194068 127764
rect 193004 126252 193060 126308
rect 192556 68572 192612 68628
rect 192668 126140 192724 126196
rect 192444 67004 192500 67060
rect 191436 2828 191492 2884
rect 191548 62972 191604 63028
rect 192892 124460 192948 124516
rect 193004 6524 193060 6580
rect 193116 119308 193172 119364
rect 192892 1484 192948 1540
rect 193900 117628 193956 117684
rect 193900 7868 193956 7924
rect 193116 1372 193172 1428
rect 194124 118076 194180 118132
rect 194572 303212 194628 303268
rect 194236 66892 194292 66948
rect 194348 301532 194404 301588
rect 194348 63756 194404 63812
rect 194460 124348 194516 124404
rect 195692 314972 195748 315028
rect 194908 159180 194964 159236
rect 197932 313852 197988 313908
rect 197036 313404 197092 313460
rect 196364 306796 196420 306852
rect 196252 306684 196308 306740
rect 195692 158956 195748 159012
rect 195916 168588 195972 168644
rect 195916 159068 195972 159124
rect 194908 158284 194964 158340
rect 195804 154364 195860 154420
rect 195692 153580 195748 153636
rect 195468 151116 195524 151172
rect 194908 148204 194964 148260
rect 194908 147868 194964 147924
rect 194684 121772 194740 121828
rect 194908 122556 194964 122612
rect 194908 121324 194964 121380
rect 194572 118636 194628 118692
rect 194684 121100 194740 121156
rect 194460 13244 194516 13300
rect 194572 116732 194628 116788
rect 194572 9884 194628 9940
rect 194124 7084 194180 7140
rect 194012 1148 194068 1204
rect 194460 4060 194516 4116
rect 192668 700 192724 756
rect 194796 119980 194852 120036
rect 195468 119980 195524 120036
rect 195692 149660 195748 149716
rect 194796 119644 194852 119700
rect 195468 116396 195524 116452
rect 194796 4732 194852 4788
rect 194908 12684 194964 12740
rect 194684 1260 194740 1316
rect 195468 7196 195524 7252
rect 195804 124348 195860 124404
rect 195804 122668 195860 122724
rect 195804 9772 195860 9828
rect 196028 155820 196084 155876
rect 196252 154364 196308 154420
rect 196364 151116 196420 151172
rect 196476 169036 196532 169092
rect 196476 158284 196532 158340
rect 196028 138796 196084 138852
rect 196140 147980 196196 148036
rect 196028 121324 196084 121380
rect 196364 147868 196420 147924
rect 196140 13356 196196 13412
rect 196252 146412 196308 146468
rect 196028 10444 196084 10500
rect 196252 8652 196308 8708
rect 196364 7532 196420 7588
rect 195916 6412 195972 6468
rect 195692 4396 195748 4452
rect 197484 310380 197540 310436
rect 197372 309932 197428 309988
rect 197372 168028 197428 168084
rect 197820 310268 197876 310324
rect 197708 303660 197764 303716
rect 197484 159740 197540 159796
rect 197372 158396 197428 158452
rect 197036 152460 197092 152516
rect 197148 157164 197204 157220
rect 196588 152236 196644 152292
rect 196588 142156 196644 142212
rect 197148 141932 197204 141988
rect 197260 154476 197316 154532
rect 197260 153020 197316 153076
rect 197260 122556 197316 122612
rect 197372 146300 197428 146356
rect 196588 14252 196644 14308
rect 197596 303436 197652 303492
rect 197596 154476 197652 154532
rect 197484 142828 197540 142884
rect 197820 153580 197876 153636
rect 208348 313852 208404 313908
rect 197932 156044 197988 156100
rect 197708 151340 197764 151396
rect 197372 6188 197428 6244
rect 197484 131180 197540 131236
rect 196588 4060 196644 4116
rect 197596 6076 197652 6132
rect 197708 119532 197764 119588
rect 197484 3164 197540 3220
rect 196476 2716 196532 2772
rect 197820 151004 197876 151060
rect 197932 147868 197988 147924
rect 198044 313740 198100 313796
rect 213388 313740 213444 313796
rect 199164 313628 199220 313684
rect 199052 310156 199108 310212
rect 198828 306908 198884 306964
rect 198716 302204 198772 302260
rect 198156 177996 198212 178052
rect 198716 177996 198772 178052
rect 198156 160076 198212 160132
rect 198156 159628 198212 159684
rect 198268 161308 198324 161364
rect 198268 157276 198324 157332
rect 198716 159628 198772 159684
rect 198044 152796 198100 152852
rect 198380 152348 198436 152404
rect 198380 148876 198436 148932
rect 198716 147980 198772 148036
rect 198828 156492 198884 156548
rect 198940 303548 198996 303604
rect 216748 313628 216804 313684
rect 199388 313516 199444 313572
rect 199164 159628 199220 159684
rect 199276 311836 199332 311892
rect 199276 159852 199332 159908
rect 199052 159404 199108 159460
rect 199052 158396 199108 158452
rect 198044 146412 198100 146468
rect 198156 142940 198212 142996
rect 197820 118412 197876 118468
rect 197932 119420 197988 119476
rect 197820 116172 197876 116228
rect 197932 9212 197988 9268
rect 198044 104076 198100 104132
rect 197708 812 197764 868
rect 197820 4060 197876 4116
rect 197932 2604 197988 2660
rect 198828 142940 198884 142996
rect 199052 156268 199108 156324
rect 199052 146188 199108 146244
rect 198492 13356 198548 13412
rect 198156 8428 198212 8484
rect 198268 10220 198324 10276
rect 198828 13244 198884 13300
rect 198492 8540 198548 8596
rect 198604 12572 198660 12628
rect 198604 4508 198660 4564
rect 198828 2492 198884 2548
rect 198940 10892 198996 10948
rect 198268 1596 198324 1652
rect 198044 1036 198100 1092
rect 199164 153132 199220 153188
rect 220108 313516 220164 313572
rect 225148 310380 225204 310436
rect 228508 310268 228564 310324
rect 231868 310156 231924 310212
rect 240268 311836 240324 311892
rect 235228 306908 235284 306964
rect 243628 303660 243684 303716
rect 246988 303548 247044 303604
rect 255388 313404 255444 313460
rect 250348 303436 250404 303492
rect 262108 306796 262164 306852
rect 270508 310044 270564 310100
rect 273868 309932 273924 309988
rect 265468 306684 265524 306740
rect 258748 302204 258804 302260
rect 282268 313292 282324 313348
rect 289884 315084 289940 315140
rect 285628 305228 285684 305284
rect 308924 316988 308980 317044
rect 304108 310156 304164 310212
rect 300748 310044 300804 310100
rect 297388 309932 297444 309988
rect 312508 306684 312564 306740
rect 292348 305116 292404 305172
rect 319228 313292 319284 313348
rect 315868 303436 315924 303492
rect 330988 313516 331044 313572
rect 327628 313404 327684 313460
rect 339388 316876 339444 316932
rect 347004 316988 347060 317044
rect 354620 317100 354676 317156
rect 350812 316876 350868 316932
rect 342748 313628 342804 313684
rect 357868 312508 357924 312564
rect 361228 315868 361284 315924
rect 366044 316764 366100 316820
rect 362236 315868 362292 315924
rect 361228 311724 361284 311780
rect 357868 308364 357924 308420
rect 334348 303548 334404 303604
rect 322588 303324 322644 303380
rect 277228 302092 277284 302148
rect 404012 319116 404068 319172
rect 397852 317212 397908 317268
rect 378140 317100 378196 317156
rect 372988 303212 373044 303268
rect 376348 313516 376404 313572
rect 378028 313404 378084 313460
rect 376348 302540 376404 302596
rect 377020 313292 377076 313348
rect 369628 301980 369684 302036
rect 301308 160188 301364 160244
rect 202300 159516 202356 159572
rect 199388 157612 199444 157668
rect 199388 156268 199444 156324
rect 199948 158956 200004 159012
rect 199388 151228 199444 151284
rect 202524 156380 202580 156436
rect 201180 153020 201236 153076
rect 201180 152684 201236 152740
rect 199948 151228 200004 151284
rect 206892 158284 206948 158340
rect 206108 156156 206164 156212
rect 206668 158172 206724 158228
rect 206668 156156 206724 156212
rect 206780 156268 206836 156324
rect 206780 154364 206836 154420
rect 202524 151004 202580 151060
rect 203308 154140 203364 154196
rect 204988 152908 205044 152964
rect 204988 151900 205044 151956
rect 207004 156492 207060 156548
rect 217532 159516 217588 159572
rect 218204 160076 218260 160132
rect 218204 159516 218260 159572
rect 213724 156828 213780 156884
rect 213948 158172 214004 158228
rect 209916 156044 209972 156100
rect 213052 156268 213108 156324
rect 207004 154476 207060 154532
rect 209356 154476 209412 154532
rect 209916 154252 209972 154308
rect 213052 154028 213108 154084
rect 209916 151116 209972 151172
rect 225148 159740 225204 159796
rect 226828 159964 226884 160020
rect 221340 157612 221396 157668
rect 225260 159628 225316 159684
rect 223804 157276 223860 157332
rect 215068 153916 215124 153972
rect 213948 151004 214004 151060
rect 209356 150892 209412 150948
rect 206892 150780 206948 150836
rect 223356 152684 223412 152740
rect 215068 152572 215124 152628
rect 216748 152572 216804 152628
rect 216748 151116 216804 151172
rect 223804 152684 223860 152740
rect 223356 151116 223412 151172
rect 215068 151004 215124 151060
rect 226828 157276 226884 157332
rect 228508 159740 228564 159796
rect 225260 150892 225316 150948
rect 225484 151900 225540 151956
rect 240380 159852 240436 159908
rect 236572 159628 236628 159684
rect 232764 159404 232820 159460
rect 230300 159068 230356 159124
rect 230188 158172 230244 158228
rect 230188 154364 230244 154420
rect 238812 158172 238868 158228
rect 230300 154140 230356 154196
rect 238700 154140 238756 154196
rect 228956 153580 229012 153636
rect 238588 154028 238644 154084
rect 238588 151116 238644 151172
rect 228508 151004 228564 151060
rect 238700 151004 238756 151060
rect 225484 150892 225540 150948
rect 251804 154028 251860 154084
rect 252028 158060 252084 158116
rect 247996 152796 248052 152852
rect 244188 152572 244244 152628
rect 253820 158060 253876 158116
rect 253708 154252 253764 154308
rect 253708 152796 253764 152852
rect 253820 152684 253876 152740
rect 252028 151116 252084 151172
rect 253708 152572 253764 152628
rect 259420 159516 259476 159572
rect 260764 154588 260820 154644
rect 262108 154588 262164 154644
rect 262108 153804 262164 153860
rect 263788 159180 263844 159236
rect 263788 153916 263844 153972
rect 263900 158172 263956 158228
rect 263228 152796 263284 152852
rect 263900 152796 263956 152852
rect 260764 152684 260820 152740
rect 269388 160076 269444 160132
rect 269276 158060 269332 158116
rect 274652 160076 274708 160132
rect 270844 157612 270900 157668
rect 269388 155932 269444 155988
rect 270396 156380 270452 156436
rect 269276 154252 269332 154308
rect 270396 154028 270452 154084
rect 286076 159740 286132 159796
rect 282268 159180 282324 159236
rect 285628 158172 285684 158228
rect 283836 158060 283892 158116
rect 283836 157612 283892 157668
rect 282156 156044 282212 156100
rect 285628 156044 285684 156100
rect 297500 160076 297556 160132
rect 300748 159740 300804 159796
rect 300748 157724 300804 157780
rect 301308 157500 301364 157556
rect 304444 160076 304500 160132
rect 293692 157388 293748 157444
rect 289884 154364 289940 154420
rect 294252 156268 294308 156324
rect 294252 154364 294308 154420
rect 282156 154252 282212 154308
rect 313404 159628 313460 159684
rect 308924 159068 308980 159124
rect 305116 157836 305172 157892
rect 309148 158172 309204 158228
rect 309148 157836 309204 157892
rect 315420 158172 315476 158228
rect 305116 157612 305172 157668
rect 304444 154252 304500 154308
rect 278460 153804 278516 153860
rect 283388 153804 283444 153860
rect 267036 152572 267092 152628
rect 255612 152460 255668 152516
rect 283388 152460 283444 152516
rect 320348 157836 320404 157892
rect 320012 157500 320068 157556
rect 320012 155932 320068 155988
rect 316540 154364 316596 154420
rect 319116 154588 319172 154644
rect 319116 154140 319172 154196
rect 315420 151116 315476 151172
rect 317212 153356 317268 153412
rect 327964 159404 328020 159460
rect 330652 159852 330708 159908
rect 329756 158060 329812 158116
rect 330876 159628 330932 159684
rect 335580 159740 335636 159796
rect 331772 159628 331828 159684
rect 330876 159068 330932 159124
rect 330652 157612 330708 157668
rect 346108 159964 346164 160020
rect 347004 159516 347060 159572
rect 346108 159404 346164 159460
rect 350812 159180 350868 159236
rect 343196 158172 343252 158228
rect 343196 157724 343252 157780
rect 354620 157612 354676 157668
rect 358428 157500 358484 157556
rect 359548 157388 359604 157444
rect 339388 157164 339444 157220
rect 356188 157276 356244 157332
rect 329756 156044 329812 156100
rect 332668 156380 332724 156436
rect 324156 152572 324212 152628
rect 348012 156380 348068 156436
rect 344652 156268 344708 156324
rect 343308 156044 343364 156100
rect 343196 155932 343252 155988
rect 342188 154588 342244 154644
rect 342188 154140 342244 154196
rect 343196 154140 343252 154196
rect 347900 156156 347956 156212
rect 357980 157164 358036 157220
rect 356188 156156 356244 156212
rect 357868 156380 357924 156436
rect 357868 156044 357924 156100
rect 357980 155820 358036 155876
rect 366044 158956 366100 159012
rect 362236 157388 362292 157444
rect 369852 156940 369908 156996
rect 359548 155820 359604 155876
rect 344652 154252 344708 154308
rect 343308 153916 343364 153972
rect 359548 153804 359604 153860
rect 359548 152684 359604 152740
rect 362796 153244 362852 153300
rect 362796 152684 362852 152740
rect 332668 152572 332724 152628
rect 317212 151116 317268 151172
rect 363356 152460 363412 152516
rect 253708 151004 253764 151060
rect 238812 150892 238868 150948
rect 214956 150780 215012 150836
rect 203308 150556 203364 150612
rect 377020 157836 377076 157892
rect 377020 156268 377076 156324
rect 377132 310044 377188 310100
rect 373660 152348 373716 152404
rect 377468 303548 377524 303604
rect 377244 303324 377300 303380
rect 377356 302540 377412 302596
rect 377356 159628 377412 159684
rect 378140 305676 378196 305732
rect 378252 316988 378308 317044
rect 378028 302428 378084 302484
rect 383068 316876 383124 316932
rect 379708 315868 379764 315924
rect 379036 313628 379092 313684
rect 378252 301868 378308 301924
rect 378252 300860 378308 300916
rect 378364 310156 378420 310212
rect 378364 160860 378420 160916
rect 378588 305676 378644 305732
rect 378588 305004 378644 305060
rect 377468 159740 377524 159796
rect 378140 159964 378196 160020
rect 378140 159628 378196 159684
rect 377468 157276 377524 157332
rect 378028 159068 378084 159124
rect 378028 158060 378084 158116
rect 377244 156044 377300 156100
rect 377356 156268 377412 156324
rect 377132 154140 377188 154196
rect 363356 150556 363412 150612
rect 199388 150332 199444 150388
rect 199164 122780 199220 122836
rect 199388 144508 199444 144564
rect 199164 7756 199220 7812
rect 199276 17612 199332 17668
rect 203196 10444 203252 10500
rect 200172 10332 200228 10388
rect 202300 8316 202356 8372
rect 200172 7420 200228 7476
rect 203196 6860 203252 6916
rect 205100 9548 205156 9604
rect 199388 6748 199444 6804
rect 199948 6748 200004 6804
rect 199948 4620 200004 4676
rect 204540 5852 204596 5908
rect 199276 4284 199332 4340
rect 202300 4284 202356 4340
rect 199052 3836 199108 3892
rect 201180 4060 201236 4116
rect 206108 8204 206164 8260
rect 213724 8652 213780 8708
rect 217532 8540 217588 8596
rect 209916 7532 209972 7588
rect 206780 6860 206836 6916
rect 205100 5852 205156 5908
rect 206668 6748 206724 6804
rect 206668 5740 206724 5796
rect 206780 4620 206836 4676
rect 205660 4508 205716 4564
rect 204988 4172 205044 4228
rect 204988 3164 205044 3220
rect 205212 3164 205268 3220
rect 205212 2604 205268 2660
rect 205548 2604 205604 2660
rect 205324 2492 205380 2548
rect 225148 6076 225204 6132
rect 223356 5852 223412 5908
rect 223356 4956 223412 5012
rect 224924 5068 224980 5124
rect 221340 3836 221396 3892
rect 207900 3724 207956 3780
rect 236572 8428 236628 8484
rect 232764 6188 232820 6244
rect 228956 4396 229012 4452
rect 230188 5964 230244 6020
rect 230300 5180 230356 5236
rect 230300 4956 230356 5012
rect 240380 4508 240436 4564
rect 230188 4396 230244 4452
rect 224924 1596 224980 1652
rect 247996 7756 248052 7812
rect 251804 4620 251860 4676
rect 259420 6300 259476 6356
rect 263228 4732 263284 4788
rect 255612 4396 255668 4452
rect 270844 6412 270900 6468
rect 274652 4844 274708 4900
rect 277228 4844 277284 4900
rect 278460 4844 278516 4900
rect 277228 2828 277284 2884
rect 286076 2940 286132 2996
rect 282268 2716 282324 2772
rect 267036 2604 267092 2660
rect 297388 6300 297444 6356
rect 301308 4732 301364 4788
rect 308924 7868 308980 7924
rect 312732 6188 312788 6244
rect 320348 8540 320404 8596
rect 316540 6076 316596 6132
rect 305116 4620 305172 4676
rect 314972 5180 315028 5236
rect 297276 3052 297332 3108
rect 327964 8204 328020 8260
rect 324156 4508 324212 4564
rect 335580 9660 335636 9716
rect 335580 8428 335636 8484
rect 339388 7420 339444 7476
rect 347004 7868 347060 7924
rect 347788 9212 347844 9268
rect 343196 5964 343252 6020
rect 331772 4396 331828 4452
rect 341628 5068 341684 5124
rect 314972 3052 315028 3108
rect 330204 3388 330260 3444
rect 293692 2940 293748 2996
rect 330204 2828 330260 2884
rect 293692 1036 293748 1092
rect 350812 8652 350868 8708
rect 362236 8092 362292 8148
rect 358428 7980 358484 8036
rect 354620 7756 354676 7812
rect 369852 8316 369908 8372
rect 373660 7196 373716 7252
rect 366044 7084 366100 7140
rect 356188 6748 356244 6804
rect 347788 2716 347844 2772
rect 352604 5852 352660 5908
rect 341628 1036 341684 1092
rect 289884 924 289940 980
rect 244188 812 244244 868
rect 377356 8540 377412 8596
rect 377468 156044 377524 156100
rect 377244 4732 377300 4788
rect 377468 4508 377524 4564
rect 378476 159180 378532 159236
rect 378364 158172 378420 158228
rect 378140 8204 378196 8260
rect 378252 156380 378308 156436
rect 378028 6188 378084 6244
rect 378476 8652 378532 8708
rect 378812 302428 378868 302484
rect 378700 300860 378756 300916
rect 378812 159628 378868 159684
rect 378924 301980 378980 302036
rect 378700 159516 378756 159572
rect 378700 158172 378756 158228
rect 378588 157612 378644 157668
rect 378364 7868 378420 7924
rect 378924 156940 378980 156996
rect 378588 7756 378644 7812
rect 378700 154364 378756 154420
rect 378812 153916 378868 153972
rect 379036 157724 379092 157780
rect 379036 156380 379092 156436
rect 379148 312508 379204 312564
rect 379148 157500 379204 157556
rect 379148 156044 379204 156100
rect 379260 303436 379316 303492
rect 379260 154364 379316 154420
rect 379820 306684 379876 306740
rect 379820 301756 379876 301812
rect 397628 313740 397684 313796
rect 397516 313628 397572 313684
rect 397404 310380 397460 310436
rect 383068 301644 383124 301700
rect 383068 159180 383124 159236
rect 396396 306684 396452 306740
rect 379820 158060 379876 158116
rect 379708 157388 379764 157444
rect 388892 157276 388948 157332
rect 379708 154364 379764 154420
rect 383068 156044 383124 156100
rect 378924 152572 378980 152628
rect 379708 152572 379764 152628
rect 378812 6412 378868 6468
rect 378924 150556 378980 150612
rect 378700 6076 378756 6132
rect 378252 5964 378308 6020
rect 379708 8316 379764 8372
rect 386428 154364 386484 154420
rect 388892 67228 388948 67284
rect 395612 104076 395668 104132
rect 386428 8092 386484 8148
rect 383068 7980 383124 8036
rect 378924 4844 378980 4900
rect 377580 4396 377636 4452
rect 356188 2604 356244 2660
rect 397180 303548 397236 303604
rect 396396 104076 396452 104132
rect 397292 303436 397348 303492
rect 397068 159628 397124 159684
rect 395612 1148 395668 1204
rect 397292 159292 397348 159348
rect 397404 155596 397460 155652
rect 397516 157500 397572 157556
rect 397180 3052 397236 3108
rect 397628 155484 397684 155540
rect 397740 310268 397796 310324
rect 397740 152124 397796 152180
rect 397852 157276 397908 157332
rect 397964 317100 398020 317156
rect 399532 316988 399588 317044
rect 397964 157388 398020 157444
rect 397964 152236 398020 152292
rect 398076 313516 398132 313572
rect 397852 152012 397908 152068
rect 399420 313404 399476 313460
rect 398972 311724 399028 311780
rect 398860 306908 398916 306964
rect 398636 156044 398692 156100
rect 399308 310156 399364 310212
rect 399196 310044 399252 310100
rect 398748 157836 398804 157892
rect 398076 151004 398132 151060
rect 399084 309932 399140 309988
rect 399196 158396 399252 158452
rect 398860 157612 398916 157668
rect 398972 158172 399028 158228
rect 399420 158172 399476 158228
rect 397516 2828 397572 2884
rect 397740 2716 397796 2772
rect 399084 154364 399140 154420
rect 399644 316876 399700 316932
rect 399196 154140 399252 154196
rect 399420 155820 399476 155876
rect 399420 9772 399476 9828
rect 399532 154252 399588 154308
rect 399308 6524 399364 6580
rect 399084 3948 399140 4004
rect 399756 316764 399812 316820
rect 410172 317212 410228 317268
rect 413980 317100 414036 317156
rect 407708 315756 407764 315812
rect 418348 313740 418404 313796
rect 421708 313628 421764 313684
rect 425068 313516 425124 313572
rect 400316 313292 400372 313348
rect 400204 306796 400260 306852
rect 399868 158172 399924 158228
rect 399756 157724 399812 157780
rect 399756 157164 399812 157220
rect 399644 155932 399700 155988
rect 399644 153804 399700 153860
rect 428428 310380 428484 310436
rect 433468 310268 433524 310324
rect 448588 316988 448644 317044
rect 452060 316876 452116 316932
rect 455980 316764 456036 316820
rect 445228 313404 445284 313460
rect 460348 313292 460404 313348
rect 440188 311724 440244 311780
rect 436828 310156 436884 310212
rect 463708 310044 463764 310100
rect 467068 309932 467124 309988
rect 470428 306908 470484 306964
rect 475468 306796 475524 306852
rect 482188 306684 482244 306740
rect 478828 303548 478884 303604
rect 485548 303436 485604 303492
rect 490588 303324 490644 303380
rect 400316 154476 400372 154532
rect 400428 303212 400484 303268
rect 400204 151116 400260 151172
rect 502348 313292 502404 313348
rect 509180 314972 509236 315028
rect 505708 310044 505764 310100
rect 497308 309932 497364 309988
rect 493948 303212 494004 303268
rect 525420 316876 525476 316932
rect 522060 316764 522116 316820
rect 537180 316988 537236 317044
rect 539644 316652 539700 316708
rect 542668 313628 542724 313684
rect 532588 313516 532644 313572
rect 527548 313404 527604 313460
rect 517468 310156 517524 310212
rect 552524 316652 552580 316708
rect 547708 303324 547764 303380
rect 512428 303212 512484 303268
rect 560140 317100 560196 317156
rect 562828 313740 562884 313796
rect 571116 317212 571172 317268
rect 579740 317212 579796 317268
rect 578060 316988 578116 317044
rect 566188 308252 566244 308308
rect 577948 316876 578004 316932
rect 577948 305676 578004 305732
rect 574588 304892 574644 304948
rect 554428 301644 554484 301700
rect 400652 154476 400708 154532
rect 407148 159516 407204 159572
rect 414652 157388 414708 157444
rect 410844 157276 410900 157332
rect 422268 157500 422324 157556
rect 418460 155484 418516 155540
rect 429884 155596 429940 155652
rect 445228 157724 445284 157780
rect 441308 157612 441364 157668
rect 452732 155932 452788 155988
rect 448924 155820 448980 155876
rect 456540 154252 456596 154308
rect 459452 154812 459508 154868
rect 437500 154140 437556 154196
rect 433692 152572 433748 152628
rect 426076 151004 426132 151060
rect 403228 149436 403284 149492
rect 400652 149324 400708 149380
rect 460348 154812 460404 154868
rect 471772 157836 471828 157892
rect 467964 155932 468020 155988
rect 464156 154364 464212 154420
rect 479388 159628 479444 159684
rect 475580 151116 475636 151172
rect 481292 154812 481348 154868
rect 459452 149324 459508 149380
rect 399532 2604 399588 2660
rect 490812 159404 490868 159460
rect 487004 159292 487060 159348
rect 483196 154812 483252 154868
rect 493052 154812 493108 154868
rect 481292 104076 481348 104132
rect 400652 102396 400708 102452
rect 398972 1484 399028 1540
rect 398860 1372 398916 1428
rect 494620 154812 494676 154868
rect 493052 102396 493108 102452
rect 496412 151116 496468 151172
rect 498428 151116 498484 151172
rect 509852 158844 509908 158900
rect 513212 159404 513268 159460
rect 506044 157276 506100 157332
rect 506044 153692 506100 153748
rect 503132 152572 503188 152628
rect 496412 7308 496468 7364
rect 521276 156156 521332 156212
rect 525196 156044 525252 156100
rect 528332 155932 528388 155988
rect 528332 155148 528388 155204
rect 532700 157724 532756 157780
rect 518252 154364 518308 154420
rect 517356 138572 517412 138628
rect 517356 101500 517412 101556
rect 513212 9884 513268 9940
rect 516572 100828 516628 100884
rect 517356 100828 517412 100884
rect 519036 153692 519092 153748
rect 532700 152796 532756 152852
rect 540316 157052 540372 157108
rect 544124 155820 544180 155876
rect 547708 157612 547764 157668
rect 551068 159292 551124 159348
rect 551068 156268 551124 156324
rect 555548 157500 555604 157556
rect 555548 155372 555604 155428
rect 559468 159180 559524 159236
rect 547708 154028 547764 154084
rect 566972 158732 567028 158788
rect 570780 157836 570836 157892
rect 563612 157388 563668 157444
rect 563612 156268 563668 156324
rect 559468 152684 559524 152740
rect 544124 150444 544180 150500
rect 535948 138572 536004 138628
rect 519036 84924 519092 84980
rect 530908 12572 530964 12628
rect 518252 9996 518308 10052
rect 516572 8428 516628 8484
rect 503132 6636 503188 6692
rect 556108 5852 556164 5908
rect 567868 12572 567924 12628
rect 400652 1260 400708 1316
rect 397068 1036 397124 1092
rect 578284 316764 578340 316820
rect 578060 153692 578116 153748
rect 578172 313292 578228 313348
rect 578508 313628 578564 313684
rect 578284 156156 578340 156212
rect 578396 313404 578452 313460
rect 578396 155932 578452 155988
rect 579628 309932 579684 309988
rect 578620 305676 578676 305732
rect 578620 304108 578676 304164
rect 578732 301644 578788 301700
rect 578732 157500 578788 157556
rect 578620 156044 578676 156100
rect 578508 155820 578564 155876
rect 578172 152572 578228 152628
rect 581420 317100 581476 317156
rect 581308 316652 581364 316708
rect 579964 313516 580020 313572
rect 579740 157836 579796 157892
rect 579852 310156 579908 310212
rect 579964 157724 580020 157780
rect 580076 310044 580132 310100
rect 580188 303324 580244 303380
rect 580300 303212 580356 303268
rect 580300 159404 580356 159460
rect 581308 159292 581364 159348
rect 581420 159180 581476 159236
rect 584668 313740 584724 313796
rect 580188 157612 580244 157668
rect 587244 406700 587300 406756
rect 589708 395612 589764 395668
rect 587356 362348 587412 362404
rect 587356 311612 587412 311668
rect 587244 306572 587300 306628
rect 587132 301532 587188 301588
rect 584668 157388 584724 157444
rect 580076 157276 580132 157332
rect 579852 154364 579908 154420
rect 579628 151116 579684 151172
rect 590044 439964 590100 440020
rect 589820 319116 589876 319172
rect 589932 351260 589988 351316
rect 589708 149436 589764 149492
rect 589820 295820 589876 295876
rect 590044 315756 590100 315812
rect 589932 159516 589988 159572
rect 589820 84028 589876 84084
rect 574588 2492 574644 2548
<< metal3 >>
rect 9874 587916 9884 587972
rect 9940 587916 9996 587972
rect 10052 587916 10062 587972
rect 190642 587468 190652 587524
rect 190708 587468 205884 587524
rect 205940 587468 205950 587524
rect 3266 587356 3276 587412
rect 3332 587356 26012 587412
rect 26068 587356 26078 587412
rect 196466 587356 196476 587412
rect 196532 587356 222236 587412
rect 222292 587356 222302 587412
rect 8306 587244 8316 587300
rect 8372 587244 75068 587300
rect 75124 587244 75134 587300
rect 157042 587244 157052 587300
rect 157108 587244 188972 587300
rect 189028 587244 189038 587300
rect 197362 587244 197372 587300
rect 197428 587244 402108 587300
rect 402164 587244 402174 587300
rect 9986 587132 9996 587188
rect 10052 587132 91420 587188
rect 91476 587132 91486 587188
rect 140690 587132 140700 587188
rect 140756 587132 189868 587188
rect 189924 587132 189934 587188
rect 194002 587132 194012 587188
rect 194068 587132 467516 587188
rect 467572 587132 467582 587188
rect 591560 584164 593000 584360
rect 591500 584136 593000 584164
rect 591500 584108 591640 584136
rect 591500 584052 591556 584108
rect -960 583800 480 584024
rect 591500 583996 591668 584052
rect 591612 583044 591668 583996
rect 192322 582988 192332 583044
rect 192388 582988 591668 583044
rect -960 572936 480 573160
rect 591560 573048 593000 573272
rect -960 562100 480 562296
rect -960 562072 532 562100
rect 392 562044 532 562072
rect 476 561988 532 562044
rect 364 561932 532 561988
rect 591560 561960 593000 562184
rect 364 561204 420 561932
rect 364 561148 194012 561204
rect 194068 561148 194078 561204
rect -960 551236 480 551432
rect -960 551208 7644 551236
rect 392 551180 7644 551208
rect 7700 551180 7710 551236
rect 591560 550872 593000 551096
rect -960 540344 480 540568
rect 591560 539812 593000 540008
rect 591500 539784 593000 539812
rect 591500 539756 591640 539784
rect 591500 539700 591556 539756
rect 591500 539644 591668 539700
rect 591612 539364 591668 539644
rect 190866 539308 190876 539364
rect 190932 539308 591668 539364
rect -960 529480 480 529704
rect 591560 528696 593000 528920
rect -960 518644 480 518840
rect -960 518616 532 518644
rect 392 518588 532 518616
rect 476 518532 532 518588
rect 364 518476 532 518532
rect 364 517524 420 518476
rect 591560 517608 593000 517832
rect 364 517468 194124 517524
rect 194180 517468 194190 517524
rect -960 507780 480 507976
rect -960 507752 7532 507780
rect 392 507724 7532 507752
rect 7588 507724 7598 507780
rect 591560 506520 593000 506744
rect -960 496888 480 497112
rect 591560 495460 593000 495656
rect 591500 495432 593000 495460
rect 591500 495404 591640 495432
rect 591500 495348 591556 495404
rect 591500 495292 591668 495348
rect 591612 494004 591668 495292
rect 197586 493948 197596 494004
rect 197652 493948 591668 494004
rect -960 486024 480 486248
rect 591560 484372 593000 484568
rect 589810 484316 589820 484372
rect 589876 484344 593000 484372
rect 589876 484316 591640 484344
rect -960 475188 480 475384
rect -960 475160 5852 475188
rect 392 475132 5852 475160
rect 5908 475132 5918 475188
rect 591560 473256 593000 473480
rect -960 464324 480 464520
rect -960 464296 7868 464324
rect 392 464268 7868 464296
rect 7924 464268 7934 464324
rect 591560 462168 593000 462392
rect 192434 461132 192444 461188
rect 192500 461132 532588 461188
rect 532644 461132 532654 461188
rect -960 453432 480 453656
rect 591560 451108 593000 451304
rect 587122 451052 587132 451108
rect 587188 451080 593000 451108
rect 587188 451052 591640 451080
rect -960 442568 480 442792
rect 591560 440020 593000 440216
rect 590034 439964 590044 440020
rect 590100 439992 593000 440020
rect 590100 439964 591640 439992
rect -960 431844 480 431928
rect -960 431788 3388 431844
rect 3444 431788 3454 431844
rect -960 431704 480 431788
rect 591560 428904 593000 429128
rect -960 420868 480 421064
rect -960 420840 4172 420868
rect 392 420812 4172 420840
rect 4228 420812 4238 420868
rect 591560 417816 593000 418040
rect -960 409976 480 410200
rect 591560 406756 593000 406952
rect 587234 406700 587244 406756
rect 587300 406728 593000 406756
rect 587300 406700 591640 406728
rect -960 399112 480 399336
rect 591560 395668 593000 395864
rect 589698 395612 589708 395668
rect 589764 395640 593000 395668
rect 589764 395612 591640 395640
rect -960 388276 480 388472
rect -960 388248 4284 388276
rect 392 388220 4284 388248
rect 4340 388220 4350 388276
rect 591560 384552 593000 384776
rect -960 377412 480 377608
rect -960 377384 4396 377412
rect 392 377356 4396 377384
rect 4452 377356 4462 377412
rect 591560 373464 593000 373688
rect -960 366520 480 366744
rect 591560 362404 593000 362600
rect 587346 362348 587356 362404
rect 587412 362376 593000 362404
rect 587412 362348 591640 362376
rect -960 355656 480 355880
rect 591560 351316 593000 351512
rect 589922 351260 589932 351316
rect 589988 351288 593000 351316
rect 589988 351260 591640 351288
rect -960 344820 480 345016
rect -960 344792 4508 344820
rect 392 344764 4508 344792
rect 4564 344764 4574 344820
rect 591560 340200 593000 340424
rect -960 333956 480 334152
rect -960 333928 4732 333956
rect 392 333900 4732 333928
rect 4788 333900 4798 333956
rect 591560 329112 593000 329336
rect -960 323064 480 323288
rect 3164 321020 3388 321076
rect 3444 321020 3454 321076
rect 3164 320964 3220 321020
rect 3154 320908 3164 320964
rect 3220 320908 3230 320964
rect 3266 319228 3276 319284
rect 3332 319228 13244 319284
rect 13300 319228 13310 319284
rect 188962 319228 188972 319284
rect 189028 319228 202300 319284
rect 202356 319228 202366 319284
rect 9986 319116 9996 319172
rect 10052 319116 17052 319172
rect 17108 319116 17118 319172
rect 196466 319116 196476 319172
rect 196532 319116 206108 319172
rect 206164 319116 206174 319172
rect 404002 319116 404012 319172
rect 404068 319116 589820 319172
rect 589876 319116 589886 319172
rect 591560 318052 593000 318248
rect 591500 318024 593000 318052
rect 591500 317996 591640 318024
rect 591500 317940 591556 317996
rect 591500 317884 591668 317940
rect 591612 317604 591668 317884
rect 192546 317548 192556 317604
rect 192612 317548 591668 317604
rect 9650 317324 9660 317380
rect 9716 317324 32284 317380
rect 32340 317324 32350 317380
rect 184594 317324 184604 317380
rect 184660 317324 191548 317380
rect 191604 317324 191614 317380
rect 9762 317212 9772 317268
rect 9828 317212 39900 317268
rect 39956 317212 39966 317268
rect 176978 317212 176988 317268
rect 177044 317212 188300 317268
rect 188356 317212 188366 317268
rect 397842 317212 397852 317268
rect 397908 317212 410172 317268
rect 410228 317212 410238 317268
rect 571106 317212 571116 317268
rect 571172 317212 579740 317268
rect 579796 317212 579806 317268
rect 8194 317100 8204 317156
rect 8260 317100 43708 317156
rect 43764 317100 43774 317156
rect 150322 317100 150332 317156
rect 150388 317100 188188 317156
rect 188244 317100 188254 317156
rect 354610 317100 354620 317156
rect 354676 317100 378140 317156
rect 378196 317100 378206 317156
rect 397954 317100 397964 317156
rect 398020 317100 413980 317156
rect 414036 317100 414046 317156
rect 560130 317100 560140 317156
rect 560196 317100 581420 317156
rect 581476 317100 581486 317156
rect 8082 316988 8092 317044
rect 8148 316988 58940 317044
rect 58996 316988 59006 317044
rect 146514 316988 146524 317044
rect 146580 316988 188972 317044
rect 189028 316988 189038 317044
rect 194674 316988 194684 317044
rect 194740 316988 308924 317044
rect 308980 316988 308990 317044
rect 346994 316988 347004 317044
rect 347060 316988 378252 317044
rect 378308 316988 378318 317044
rect 399522 316988 399532 317044
rect 399588 316988 448588 317044
rect 448644 316988 448654 317044
rect 537170 316988 537180 317044
rect 537236 316988 578060 317044
rect 578116 316988 578126 317044
rect 7970 316876 7980 316932
rect 8036 316876 62748 316932
rect 62804 316876 62814 316932
rect 131282 316876 131292 316932
rect 131348 316876 189644 316932
rect 189700 316876 189710 316932
rect 197474 316876 197484 316932
rect 197540 316876 339388 316932
rect 339444 316876 339454 316932
rect 350802 316876 350812 316932
rect 350868 316876 383068 316932
rect 383124 316876 383134 316932
rect 399634 316876 399644 316932
rect 399700 316876 452060 316932
rect 452116 316876 452126 316932
rect 525410 316876 525420 316932
rect 525476 316876 577948 316932
rect 578004 316876 578014 316932
rect 9874 316764 9884 316820
rect 9940 316764 85596 316820
rect 85652 316764 85662 316820
rect 112242 316764 112252 316820
rect 112308 316764 188076 316820
rect 188132 316764 188142 316820
rect 189186 316764 189196 316820
rect 189252 316764 366044 316820
rect 366100 316764 366110 316820
rect 399746 316764 399756 316820
rect 399812 316764 455980 316820
rect 456036 316764 456046 316820
rect 522050 316764 522060 316820
rect 522116 316764 578284 316820
rect 578340 316764 578350 316820
rect 6626 316652 6636 316708
rect 6692 316652 89404 316708
rect 89460 316652 89470 316708
rect 97010 316652 97020 316708
rect 97076 316652 189420 316708
rect 189476 316652 189486 316708
rect 190754 316652 190764 316708
rect 190820 316652 539644 316708
rect 539700 316652 539710 316708
rect 552514 316652 552524 316708
rect 552580 316652 581308 316708
rect 581364 316652 581374 316708
rect 361218 315868 361228 315924
rect 361284 315868 362236 315924
rect 362292 315868 379708 315924
rect 379764 315868 379774 315924
rect 407698 315756 407708 315812
rect 407764 315756 590044 315812
rect 590100 315756 590110 315812
rect 198146 315084 198156 315140
rect 198212 315084 289884 315140
rect 289940 315084 289950 315140
rect 195682 314972 195692 315028
rect 195748 314972 509180 315028
rect 509236 314972 509246 315028
rect 197922 313852 197932 313908
rect 197988 313852 208348 313908
rect 208404 313852 208414 313908
rect 9986 313740 9996 313796
rect 10052 313740 47068 313796
rect 47124 313740 47134 313796
rect 198034 313740 198044 313796
rect 198100 313740 213388 313796
rect 213444 313740 213454 313796
rect 397618 313740 397628 313796
rect 397684 313740 418348 313796
rect 418404 313740 418414 313796
rect 562818 313740 562828 313796
rect 562884 313740 584668 313796
rect 584724 313740 584734 313796
rect 9874 313628 9884 313684
rect 9940 313628 50428 313684
rect 50484 313628 50494 313684
rect 161298 313628 161308 313684
rect 161364 313628 191212 313684
rect 191268 313628 191278 313684
rect 199154 313628 199164 313684
rect 199220 313628 216748 313684
rect 216804 313628 216814 313684
rect 342738 313628 342748 313684
rect 342804 313628 379036 313684
rect 379092 313628 379102 313684
rect 397506 313628 397516 313684
rect 397572 313628 421708 313684
rect 421764 313628 421774 313684
rect 542658 313628 542668 313684
rect 542724 313628 578508 313684
rect 578564 313628 578574 313684
rect 7634 313516 7644 313572
rect 7700 313516 53788 313572
rect 53844 313516 53854 313572
rect 157938 313516 157948 313572
rect 158004 313516 190988 313572
rect 191044 313516 191054 313572
rect 199378 313516 199388 313572
rect 199444 313516 220108 313572
rect 220164 313516 220174 313572
rect 330978 313516 330988 313572
rect 331044 313516 376348 313572
rect 376404 313516 376414 313572
rect 398066 313516 398076 313572
rect 398132 313516 425068 313572
rect 425124 313516 425134 313572
rect 532578 313516 532588 313572
rect 532644 313516 579964 313572
rect 580020 313516 580030 313572
rect 9762 313404 9772 313460
rect 9828 313404 65548 313460
rect 65604 313404 65614 313460
rect 152898 313404 152908 313460
rect 152964 313404 190652 313460
rect 190708 313404 190718 313460
rect 197026 313404 197036 313460
rect 197092 313404 255388 313460
rect 255444 313404 255454 313460
rect 327618 313404 327628 313460
rect 327684 313404 378028 313460
rect 378084 313404 378094 313460
rect 399410 313404 399420 313460
rect 399476 313404 445228 313460
rect 445284 313404 445294 313460
rect 527538 313404 527548 313460
rect 527604 313404 578396 313460
rect 578452 313404 578462 313460
rect 10434 313292 10444 313348
rect 10500 313292 68908 313348
rect 68964 313292 68974 313348
rect 115938 313292 115948 313348
rect 116004 313292 189980 313348
rect 190036 313292 190046 313348
rect 199602 313292 199612 313348
rect 199668 313292 282268 313348
rect 282324 313292 282334 313348
rect 319218 313292 319228 313348
rect 319284 313292 377020 313348
rect 377076 313292 377086 313348
rect 400306 313292 400316 313348
rect 400372 313292 460348 313348
rect 460404 313292 460414 313348
rect 502338 313292 502348 313348
rect 502404 313292 578172 313348
rect 578228 313292 578238 313348
rect 357858 312508 357868 312564
rect 357924 312508 379148 312564
rect 379204 312508 379214 312564
rect -960 312200 480 312424
rect 199266 311836 199276 311892
rect 199332 311836 240268 311892
rect 240324 311836 240334 311892
rect 173058 311724 173068 311780
rect 173124 311724 188748 311780
rect 188804 311724 361228 311780
rect 361284 311724 361294 311780
rect 398962 311724 398972 311780
rect 399028 311724 440188 311780
rect 440244 311724 440254 311780
rect 194226 311612 194236 311668
rect 194292 311612 587356 311668
rect 587412 311612 587422 311668
rect 197474 310380 197484 310436
rect 197540 310380 225148 310436
rect 225204 310380 225214 310436
rect 397394 310380 397404 310436
rect 397460 310380 428428 310436
rect 428484 310380 428494 310436
rect 197810 310268 197820 310324
rect 197876 310268 228508 310324
rect 228564 310268 228574 310324
rect 397730 310268 397740 310324
rect 397796 310268 433468 310324
rect 433524 310268 433534 310324
rect 7746 310156 7756 310212
rect 7812 310156 73948 310212
rect 74004 310156 74014 310212
rect 199042 310156 199052 310212
rect 199108 310156 231868 310212
rect 231924 310156 231934 310212
rect 304098 310156 304108 310212
rect 304164 310156 378364 310212
rect 378420 310156 378430 310212
rect 399298 310156 399308 310212
rect 399364 310156 436828 310212
rect 436884 310156 436894 310212
rect 517458 310156 517468 310212
rect 517524 310156 579852 310212
rect 579908 310156 579918 310212
rect 6514 310044 6524 310100
rect 6580 310044 77308 310100
rect 77364 310044 77374 310100
rect 198034 310044 198044 310100
rect 198100 310044 270508 310100
rect 270564 310044 270574 310100
rect 300738 310044 300748 310100
rect 300804 310044 377132 310100
rect 377188 310044 377198 310100
rect 399186 310044 399196 310100
rect 399252 310044 463708 310100
rect 463764 310044 463774 310100
rect 505698 310044 505708 310100
rect 505764 310044 580076 310100
rect 580132 310044 580142 310100
rect 9538 309932 9548 309988
rect 9604 309932 119308 309988
rect 119364 309932 119374 309988
rect 164658 309932 164668 309988
rect 164724 309932 190764 309988
rect 190820 309932 190830 309988
rect 197362 309932 197372 309988
rect 197428 309932 273868 309988
rect 273924 309932 273934 309988
rect 297378 309932 297388 309988
rect 297444 309932 376348 309988
rect 376404 309932 376414 309988
rect 399074 309932 399084 309988
rect 399140 309932 467068 309988
rect 467124 309932 467134 309988
rect 497298 309932 497308 309988
rect 497364 309932 579628 309988
rect 579684 309932 579694 309988
rect 173012 308364 188860 308420
rect 188916 308364 357868 308420
rect 357924 308364 357934 308420
rect 173012 308308 173068 308364
rect 168018 308252 168028 308308
rect 168084 308252 173068 308308
rect 189074 308252 189084 308308
rect 189140 308252 566188 308308
rect 566244 308252 566254 308308
rect 122658 307020 122668 307076
rect 122724 307020 191436 307076
rect 191492 307020 191502 307076
rect 107538 306908 107548 306964
rect 107604 306908 191660 306964
rect 191716 306908 191726 306964
rect 198818 306908 198828 306964
rect 198884 306908 235228 306964
rect 235284 306908 235294 306964
rect 398850 306908 398860 306964
rect 398916 306908 470428 306964
rect 470484 306908 470494 306964
rect 591560 306936 593000 307160
rect 104178 306796 104188 306852
rect 104244 306796 193116 306852
rect 193172 306796 193182 306852
rect 196354 306796 196364 306852
rect 196420 306796 262108 306852
rect 262164 306796 262174 306852
rect 400194 306796 400204 306852
rect 400260 306796 475468 306852
rect 475524 306796 475534 306852
rect 100818 306684 100828 306740
rect 100884 306684 191884 306740
rect 191940 306684 191950 306740
rect 196242 306684 196252 306740
rect 196308 306684 265468 306740
rect 265524 306684 265534 306740
rect 312498 306684 312508 306740
rect 312564 306684 379820 306740
rect 379876 306684 379886 306740
rect 396386 306684 396396 306740
rect 396452 306684 482188 306740
rect 482244 306684 482254 306740
rect 188962 306572 188972 306628
rect 189028 306572 587244 306628
rect 587300 306572 587310 306628
rect 191874 305788 191884 305844
rect 191940 305788 198156 305844
rect 198212 305788 198222 305844
rect 378130 305676 378140 305732
rect 378196 305676 378588 305732
rect 378644 305676 378654 305732
rect 577938 305676 577948 305732
rect 578004 305676 578620 305732
rect 578676 305676 578686 305732
rect 189410 305228 189420 305284
rect 189476 305228 285628 305284
rect 285684 305228 285694 305284
rect 193106 305116 193116 305172
rect 193172 305116 199052 305172
rect 199108 305116 292348 305172
rect 292404 305116 292414 305172
rect 190754 305004 190764 305060
rect 190820 305004 378588 305060
rect 378644 305004 378654 305060
rect 195682 304892 195692 304948
rect 195748 304892 574588 304948
rect 574644 304892 574654 304948
rect 193890 304108 193900 304164
rect 193956 304108 578620 304164
rect 578676 304108 578686 304164
rect 197698 303660 197708 303716
rect 197764 303660 243628 303716
rect 243684 303660 243694 303716
rect 141138 303548 141148 303604
rect 141204 303548 188412 303604
rect 188468 303548 188478 303604
rect 198930 303548 198940 303604
rect 198996 303548 246988 303604
rect 247044 303548 247054 303604
rect 334338 303548 334348 303604
rect 334404 303548 377468 303604
rect 377524 303548 377534 303604
rect 397170 303548 397180 303604
rect 397236 303548 478828 303604
rect 478884 303548 478894 303604
rect 9426 303436 9436 303492
rect 9492 303436 26908 303492
rect 26964 303436 26974 303492
rect 137778 303436 137788 303492
rect 137844 303436 188524 303492
rect 188580 303436 188590 303492
rect 197586 303436 197596 303492
rect 197652 303436 250348 303492
rect 250404 303436 250414 303492
rect 315858 303436 315868 303492
rect 315924 303436 379260 303492
rect 379316 303436 379326 303492
rect 397282 303436 397292 303492
rect 397348 303436 485548 303492
rect 485604 303436 485614 303492
rect 9650 303324 9660 303380
rect 9716 303324 80668 303380
rect 80724 303324 80734 303380
rect 134418 303324 134428 303380
rect 134484 303324 188636 303380
rect 188692 303324 322588 303380
rect 322644 303324 377244 303380
rect 377300 303324 377310 303380
rect 397618 303324 397628 303380
rect 397684 303324 490588 303380
rect 490644 303324 490654 303380
rect 547698 303324 547708 303380
rect 547764 303324 580188 303380
rect 580244 303324 580254 303380
rect 6402 303212 6412 303268
rect 6468 303212 92428 303268
rect 92484 303212 92494 303268
rect 126018 303212 126028 303268
rect 126084 303212 190876 303268
rect 190932 303212 190942 303268
rect 194562 303212 194572 303268
rect 194628 303212 372988 303268
rect 373044 303212 373054 303268
rect 400418 303212 400428 303268
rect 400484 303212 493948 303268
rect 494004 303212 494014 303268
rect 512418 303212 512428 303268
rect 512484 303212 580300 303268
rect 580356 303212 580366 303268
rect 188402 302540 188412 302596
rect 188468 302540 376348 302596
rect 376404 302540 377356 302596
rect 377412 302540 377422 302596
rect 188514 302428 188524 302484
rect 188580 302428 378028 302484
rect 378084 302428 378812 302484
rect 378868 302428 378878 302484
rect 198706 302204 198716 302260
rect 198772 302204 258748 302260
rect 258804 302204 258814 302260
rect 192658 302092 192668 302148
rect 192724 302092 277228 302148
rect 277284 302092 277294 302148
rect 179778 301980 179788 302036
rect 179844 301980 190092 302036
rect 190148 301980 369628 302036
rect 369684 301980 378924 302036
rect 378980 301980 378990 302036
rect 190978 301868 190988 301924
rect 191044 301868 378252 301924
rect 378308 301868 378318 301924
rect 7410 301756 7420 301812
rect 7476 301756 20188 301812
rect 20244 301756 20254 301812
rect 191426 301756 191436 301812
rect 191492 301756 379820 301812
rect 379876 301756 379886 301812
rect 9090 301644 9100 301700
rect 9156 301644 23548 301700
rect 23604 301644 23614 301700
rect 191202 301644 191212 301700
rect 191268 301644 383068 301700
rect 383124 301644 383134 301700
rect 554418 301644 554428 301700
rect 554484 301644 578732 301700
rect 578788 301644 578798 301700
rect -960 301364 480 301560
rect 6290 301532 6300 301588
rect 6356 301532 35308 301588
rect 35364 301532 35374 301588
rect 194338 301532 194348 301588
rect 194404 301532 587132 301588
rect 587188 301532 587198 301588
rect -960 301336 4844 301364
rect 392 301308 4844 301336
rect 4900 301308 4910 301364
rect 378242 300860 378252 300916
rect 378308 300860 378700 300916
rect 378756 300860 378766 300916
rect 197698 300748 197708 300804
rect 197764 300748 397628 300804
rect 397684 300748 397694 300804
rect 591560 295876 593000 296072
rect 589810 295820 589820 295876
rect 589876 295848 593000 295876
rect 589876 295820 591640 295848
rect -960 290500 480 290696
rect -960 290472 4620 290500
rect 392 290444 4620 290472
rect 4676 290444 4686 290500
rect 591560 284760 593000 284984
rect -960 279608 480 279832
rect 591560 273672 593000 273896
rect -960 268884 480 268968
rect -960 268828 2492 268884
rect 2548 268828 2558 268884
rect -960 268744 480 268828
rect 591560 262584 593000 262808
rect -960 257880 480 258104
rect 591560 251496 593000 251720
rect -960 247044 480 247240
rect -960 247016 9212 247044
rect 392 246988 9212 247016
rect 9268 246988 9278 247044
rect 591560 240408 593000 240632
rect -960 236152 480 236376
rect 591560 229320 593000 229544
rect -960 225316 480 225512
rect -960 225288 532 225316
rect 392 225260 532 225288
rect 476 225204 532 225260
rect 18 225148 28 225204
rect 84 225148 532 225204
rect 591560 218232 593000 218456
rect -960 214424 480 214648
rect 591560 207144 593000 207368
rect -960 203588 480 203784
rect -960 203560 9324 203588
rect 392 203532 9324 203560
rect 9380 203532 9390 203588
rect 591560 196056 593000 196280
rect -960 192696 480 192920
rect 591560 184968 593000 185192
rect -960 181860 480 182056
rect -960 181832 2604 181860
rect 392 181804 2604 181832
rect 2660 181804 2670 181860
rect 198146 177996 198156 178052
rect 198212 177996 198716 178052
rect 198772 177996 198782 178052
rect 591560 173880 593000 174104
rect -960 170968 480 171192
rect 196466 169036 196476 169092
rect 196532 169036 199388 169092
rect 199444 169036 199454 169092
rect 195906 168588 195916 168644
rect 195972 168588 198044 168644
rect 198100 168588 198110 168644
rect 197250 168028 197260 168084
rect 197316 168028 197372 168084
rect 197428 168028 197438 168084
rect 591560 162792 593000 163016
rect 189634 161308 189644 161364
rect 189700 161308 198268 161364
rect 198324 161308 198334 161364
rect 378018 160860 378028 160916
rect 378084 160860 378364 160916
rect 378420 160860 378430 160916
rect -960 160132 480 160328
rect 188066 160188 188076 160244
rect 188132 160188 301308 160244
rect 301364 160188 301374 160244
rect -960 160104 6076 160132
rect 392 160076 6076 160104
rect 6132 160076 6142 160132
rect 198146 160076 198156 160132
rect 198212 160076 218204 160132
rect 218260 160076 218270 160132
rect 269378 160076 269388 160132
rect 269444 160076 274652 160132
rect 274708 160076 274718 160132
rect 297490 160076 297500 160132
rect 297556 160076 304444 160132
rect 304500 160076 304510 160132
rect 97458 159964 97468 160020
rect 97524 159964 226828 160020
rect 226884 159964 226894 160020
rect 346098 159964 346108 160020
rect 346164 159964 378140 160020
rect 378196 159964 378206 160020
rect 199266 159852 199276 159908
rect 199332 159852 240380 159908
rect 240436 159852 240446 159908
rect 330642 159852 330652 159908
rect 330708 159852 378028 159908
rect 378084 159852 378094 159908
rect 123666 159740 123676 159796
rect 123732 159740 191436 159796
rect 191492 159740 191502 159796
rect 197474 159740 197484 159796
rect 197540 159740 225148 159796
rect 225204 159740 225214 159796
rect 228498 159740 228508 159796
rect 228564 159740 286076 159796
rect 286132 159740 286142 159796
rect 300738 159740 300748 159796
rect 300804 159740 335580 159796
rect 335636 159740 377468 159796
rect 377524 159740 377534 159796
rect 5842 159628 5852 159684
rect 5908 159628 17052 159684
rect 17108 159628 17118 159684
rect 198146 159628 198156 159684
rect 198212 159628 198268 159684
rect 198324 159628 198334 159684
rect 198706 159628 198716 159684
rect 198772 159628 199164 159684
rect 199220 159628 202580 159684
rect 225250 159628 225260 159684
rect 225316 159628 236572 159684
rect 236628 159628 236638 159684
rect 313394 159628 313404 159684
rect 313460 159628 330876 159684
rect 330932 159628 330942 159684
rect 331762 159628 331772 159684
rect 331828 159628 377356 159684
rect 377412 159628 377422 159684
rect 378130 159628 378140 159684
rect 378196 159628 378812 159684
rect 378868 159628 378878 159684
rect 397058 159628 397068 159684
rect 397124 159628 479388 159684
rect 479444 159628 479454 159684
rect 202524 159572 202580 159628
rect 6514 159516 6524 159572
rect 6580 159516 77980 159572
rect 78036 159516 78876 159572
rect 78932 159516 78942 159572
rect 112242 159516 112252 159572
rect 112308 159516 188076 159572
rect 188132 159516 188142 159572
rect 194114 159516 194124 159572
rect 194180 159516 202300 159572
rect 202356 159516 202366 159572
rect 202524 159516 217532 159572
rect 217588 159516 217598 159572
rect 218194 159516 218204 159572
rect 218260 159516 259420 159572
rect 259476 159516 259486 159572
rect 346994 159516 347004 159572
rect 347060 159516 378700 159572
rect 378756 159516 378766 159572
rect 407138 159516 407148 159572
rect 407204 159516 589932 159572
rect 589988 159516 589998 159572
rect 7634 159404 7644 159460
rect 7700 159404 55132 159460
rect 55188 159404 56364 159460
rect 56420 159404 56430 159460
rect 199042 159404 199052 159460
rect 199108 159404 232764 159460
rect 232820 159404 232830 159460
rect 327954 159404 327964 159460
rect 328020 159404 346108 159460
rect 346164 159404 346174 159460
rect 397618 159404 397628 159460
rect 397684 159404 490812 159460
rect 490868 159404 490878 159460
rect 513202 159404 513212 159460
rect 513268 159404 580300 159460
rect 580356 159404 580366 159460
rect 9762 159292 9772 159348
rect 9828 159292 39900 159348
rect 39956 159292 39966 159348
rect 397282 159292 397292 159348
rect 397348 159292 487004 159348
rect 487060 159292 487070 159348
rect 551058 159292 551068 159348
rect 551124 159292 581308 159348
rect 581364 159292 581374 159348
rect 9650 159180 9660 159236
rect 9716 159180 32284 159236
rect 32340 159180 33292 159236
rect 33348 159180 33358 159236
rect 93202 159180 93212 159236
rect 93268 159180 194908 159236
rect 194964 159180 194974 159236
rect 263778 159180 263788 159236
rect 263844 159180 282268 159236
rect 282324 159180 282334 159236
rect 350802 159180 350812 159236
rect 350868 159180 378476 159236
rect 378532 159180 383068 159236
rect 383124 159180 383134 159236
rect 559458 159180 559468 159236
rect 559524 159180 581420 159236
rect 581476 159180 581486 159236
rect 81778 159068 81788 159124
rect 81844 159068 195916 159124
rect 195972 159068 195982 159124
rect 230290 159068 230300 159124
rect 230356 159068 308924 159124
rect 308980 159068 308990 159124
rect 330866 159068 330876 159124
rect 330932 159068 378028 159124
rect 378084 159068 378094 159124
rect 62290 158956 62300 159012
rect 62356 158956 195692 159012
rect 195748 158956 195758 159012
rect 199938 158956 199948 159012
rect 200004 158956 366044 159012
rect 366100 158956 366110 159012
rect 31938 158844 31948 158900
rect 32004 158844 197708 158900
rect 197764 158844 197774 158900
rect 197922 158844 197932 158900
rect 197988 158844 509852 158900
rect 509908 158844 509918 158900
rect 9538 158732 9548 158788
rect 9604 158732 55468 158788
rect 55524 158732 55534 158788
rect 166338 158732 166348 158788
rect 166404 158732 566972 158788
rect 567028 158732 567038 158788
rect 197362 158396 197372 158452
rect 197428 158396 199052 158452
rect 199108 158396 199118 158452
rect 398972 158396 399196 158452
rect 399252 158396 399262 158452
rect 194898 158284 194908 158340
rect 194964 158284 196476 158340
rect 196532 158284 206892 158340
rect 206948 158284 206958 158340
rect 398972 158228 399028 158396
rect 190866 158172 190876 158228
rect 190932 158172 206668 158228
rect 206724 158172 206734 158228
rect 213938 158172 213948 158228
rect 214004 158172 230188 158228
rect 230244 158172 230254 158228
rect 238802 158172 238812 158228
rect 238868 158172 263900 158228
rect 263956 158172 263966 158228
rect 285618 158172 285628 158228
rect 285684 158172 309148 158228
rect 309204 158172 309214 158228
rect 315410 158172 315420 158228
rect 315476 158172 343196 158228
rect 343252 158172 343262 158228
rect 378354 158172 378364 158228
rect 378420 158172 378700 158228
rect 378756 158172 378766 158228
rect 398962 158172 398972 158228
rect 399028 158172 399038 158228
rect 399410 158172 399420 158228
rect 399476 158172 399868 158228
rect 399924 158172 399934 158228
rect 190642 158060 190652 158116
rect 190708 158060 252028 158116
rect 252084 158060 252094 158116
rect 253810 158060 253820 158116
rect 253876 158060 269276 158116
rect 269332 158060 269342 158116
rect 283826 158060 283836 158116
rect 283892 158060 329756 158116
rect 329812 158060 329822 158116
rect 378018 158060 378028 158116
rect 378084 158060 379820 158116
rect 379876 158060 379886 158116
rect 198818 157948 198828 158004
rect 198884 157948 569604 158004
rect 569548 157892 569604 157948
rect 9090 157836 9100 157892
rect 9156 157836 24668 157892
rect 24724 157836 24734 157892
rect 169362 157836 169372 157892
rect 169428 157836 188860 157892
rect 188916 157836 188926 157892
rect 189970 157836 189980 157892
rect 190036 157836 305116 157892
rect 305172 157836 305182 157892
rect 309138 157836 309148 157892
rect 309204 157836 320348 157892
rect 320404 157836 377020 157892
rect 377076 157836 377086 157892
rect 398738 157836 398748 157892
rect 398804 157836 471772 157892
rect 471828 157836 471838 157892
rect 569548 157836 570780 157892
rect 570836 157836 579740 157892
rect 579796 157836 579806 157892
rect 7410 157724 7420 157780
rect 7476 157724 20860 157780
rect 20916 157724 22652 157780
rect 22708 157724 22718 157780
rect 188962 157724 188972 157780
rect 189028 157724 300748 157780
rect 300804 157724 300814 157780
rect 343186 157724 343196 157780
rect 343252 157724 379036 157780
rect 379092 157724 379102 157780
rect 399746 157724 399756 157780
rect 399812 157724 445228 157780
rect 445284 157724 445294 157780
rect 532690 157724 532700 157780
rect 532756 157724 579964 157780
rect 580020 157724 580030 157780
rect 6290 157612 6300 157668
rect 6356 157612 36092 157668
rect 36148 157612 36158 157668
rect 153682 157612 153692 157668
rect 153748 157612 190652 157668
rect 190708 157612 190718 157668
rect 199378 157612 199388 157668
rect 199444 157612 221340 157668
rect 221396 157612 221406 157668
rect 270834 157612 270844 157668
rect 270900 157612 283836 157668
rect 283892 157612 283902 157668
rect 305106 157612 305116 157668
rect 305172 157612 330652 157668
rect 330708 157612 330718 157668
rect 354610 157612 354620 157668
rect 354676 157612 378588 157668
rect 378644 157612 378654 157668
rect 398850 157612 398860 157668
rect 398916 157612 441308 157668
rect 441364 157612 441374 157668
rect 547698 157612 547708 157668
rect 547764 157612 580188 157668
rect 580244 157612 580254 157668
rect 9426 157500 9436 157556
rect 9492 157500 28476 157556
rect 28532 157500 28542 157556
rect 162082 157500 162092 157556
rect 162148 157500 191212 157556
rect 191268 157500 191278 157556
rect 301298 157500 301308 157556
rect 301364 157500 320012 157556
rect 320068 157500 320078 157556
rect 358418 157500 358428 157556
rect 358484 157500 379148 157556
rect 379204 157500 379214 157556
rect 397506 157500 397516 157556
rect 397572 157500 422268 157556
rect 422324 157500 422334 157556
rect 555538 157500 555548 157556
rect 555604 157500 578732 157556
rect 578788 157500 578798 157556
rect 7970 157388 7980 157444
rect 8036 157388 63084 157444
rect 63140 157388 63150 157444
rect 165554 157388 165564 157444
rect 165620 157388 190764 157444
rect 190820 157388 190830 157444
rect 293682 157388 293692 157444
rect 293748 157388 359548 157444
rect 359604 157388 359614 157444
rect 362226 157388 362236 157444
rect 362292 157388 379708 157444
rect 379764 157388 379774 157444
rect 397954 157388 397964 157444
rect 398020 157388 414652 157444
rect 414708 157388 414718 157444
rect 563602 157388 563612 157444
rect 563668 157388 584668 157444
rect 584724 157388 584734 157444
rect 3154 157276 3164 157332
rect 3220 157276 13244 157332
rect 13300 157276 13310 157332
rect 173842 157276 173852 157332
rect 173908 157276 188748 157332
rect 188804 157276 188814 157332
rect 198258 157276 198268 157332
rect 198324 157276 223804 157332
rect 223860 157276 223870 157332
rect 226818 157276 226828 157332
rect 226884 157276 356188 157332
rect 356244 157276 356254 157332
rect 377458 157276 377468 157332
rect 377524 157276 388892 157332
rect 388948 157276 388958 157332
rect 397842 157276 397852 157332
rect 397908 157276 410844 157332
rect 410900 157276 410910 157332
rect 506034 157276 506044 157332
rect 506100 157276 580076 157332
rect 580132 157276 580142 157332
rect 28466 157164 28476 157220
rect 28532 157164 46172 157220
rect 46228 157164 46238 157220
rect 56354 157164 56364 157220
rect 56420 157164 86492 157220
rect 86548 157164 86558 157220
rect 180562 157164 180572 157220
rect 180628 157164 190092 157220
rect 190148 157164 190158 157220
rect 197138 157164 197148 157220
rect 197204 157164 339388 157220
rect 339444 157164 339454 157220
rect 357970 157164 357980 157220
rect 358036 157164 399756 157220
rect 399812 157164 399822 157220
rect 39890 157052 39900 157108
rect 39956 157052 71372 157108
rect 71428 157052 71438 157108
rect 78866 157052 78876 157108
rect 78932 157052 86716 157108
rect 86772 157052 86782 157108
rect 90626 157052 90636 157108
rect 90692 157052 97020 157108
rect 97076 157052 97086 157108
rect 199602 157052 199612 157108
rect 199668 157052 540316 157108
rect 540372 157052 540382 157108
rect 8082 156940 8092 156996
rect 8148 156940 59724 156996
rect 59780 156940 59790 156996
rect 116722 156940 116732 156996
rect 116788 156940 189980 156996
rect 190036 156940 190046 156996
rect 369842 156940 369852 156996
rect 369908 156940 378924 156996
rect 378980 156940 378990 156996
rect 158722 156828 158732 156884
rect 158788 156828 190988 156884
rect 191044 156828 191054 156884
rect 211698 156828 211708 156884
rect 211764 156828 213724 156884
rect 213780 156828 213790 156884
rect 198818 156492 198828 156548
rect 198884 156492 207004 156548
rect 207060 156492 207070 156548
rect 33282 156380 33292 156436
rect 33348 156380 41132 156436
rect 41188 156380 41198 156436
rect 74162 156380 74172 156436
rect 74228 156380 78988 156436
rect 202514 156380 202524 156436
rect 202580 156380 270396 156436
rect 270452 156380 270462 156436
rect 332658 156380 332668 156436
rect 332724 156380 344484 156436
rect 348002 156380 348012 156436
rect 348068 156380 357868 156436
rect 357924 156380 357934 156436
rect 378242 156380 378252 156436
rect 378308 156380 379036 156436
rect 379092 156380 379102 156436
rect 78932 156324 78988 156380
rect 24658 156268 24668 156324
rect 24724 156268 27692 156324
rect 27748 156268 27758 156324
rect 36082 156268 36092 156324
rect 36148 156268 37772 156324
rect 37828 156268 37838 156324
rect 78932 156268 91532 156324
rect 91588 156268 91598 156324
rect 163762 156268 163772 156324
rect 163828 156268 165564 156324
rect 165620 156268 165630 156324
rect 167122 156268 167132 156324
rect 167188 156268 169372 156324
rect 169428 156268 169438 156324
rect 175522 156268 175532 156324
rect 175588 156268 176988 156324
rect 177044 156268 177054 156324
rect 199042 156268 199052 156324
rect 199108 156268 199388 156324
rect 199444 156268 199454 156324
rect 206770 156268 206780 156324
rect 206836 156268 213052 156324
rect 213108 156268 213118 156324
rect 215068 156268 294252 156324
rect 294308 156268 294318 156324
rect 215068 156212 215124 156268
rect 10434 156156 10444 156212
rect 10500 156156 69692 156212
rect 69748 156156 70364 156212
rect 70420 156156 70430 156212
rect 194002 156156 194012 156212
rect 194068 156156 206108 156212
rect 206164 156156 206174 156212
rect 206658 156156 206668 156212
rect 206724 156156 215124 156212
rect 344428 156212 344484 156380
rect 344642 156268 344652 156324
rect 344708 156268 376348 156324
rect 376404 156268 376414 156324
rect 377010 156268 377020 156324
rect 377076 156268 377356 156324
rect 377412 156268 377422 156324
rect 551030 156268 551068 156324
rect 551124 156268 551134 156324
rect 563574 156268 563612 156324
rect 563668 156268 563678 156324
rect 344428 156156 347900 156212
rect 347956 156156 347966 156212
rect 356178 156156 356188 156212
rect 356244 156156 521276 156212
rect 521332 156156 578284 156212
rect 578340 156156 578350 156212
rect 84802 156044 84812 156100
rect 84868 156044 173068 156100
rect 197922 156044 197932 156100
rect 197988 156044 209916 156100
rect 209972 156044 209982 156100
rect 282146 156044 282156 156100
rect 282212 156044 285628 156100
rect 285684 156044 285694 156100
rect 329746 156044 329756 156100
rect 329812 156044 343308 156100
rect 343364 156044 343374 156100
rect 357858 156044 357868 156100
rect 357924 156044 377244 156100
rect 377300 156044 377468 156100
rect 377524 156044 377534 156100
rect 379138 156044 379148 156100
rect 379204 156044 383068 156100
rect 383124 156044 383134 156100
rect 384692 156044 398636 156100
rect 398692 156044 455308 156100
rect 525186 156044 525196 156100
rect 525252 156044 578620 156100
rect 578676 156044 578686 156100
rect 173012 155988 173068 156044
rect 173012 155932 197260 155988
rect 197316 155932 199836 155988
rect 199892 155932 269388 155988
rect 269444 155932 269454 155988
rect 320002 155932 320012 155988
rect 320068 155932 343196 155988
rect 343252 155932 343262 155988
rect 196018 155820 196028 155876
rect 196084 155820 357980 155876
rect 358036 155820 358046 155876
rect 359538 155820 359548 155876
rect 359604 155820 378140 155876
rect 378196 155820 378206 155876
rect 384692 155764 384748 156044
rect 455252 155988 455308 156044
rect 399634 155932 399644 155988
rect 399700 155932 452732 155988
rect 452788 155932 452798 155988
rect 455252 155932 467964 155988
rect 468020 155932 468030 155988
rect 528322 155932 528332 155988
rect 528388 155932 578396 155988
rect 578452 155932 578462 155988
rect 399410 155820 399420 155876
rect 399476 155820 448924 155876
rect 448980 155820 448990 155876
rect 544114 155820 544124 155876
rect 544180 155820 578508 155876
rect 578564 155820 578574 155876
rect 195794 155708 195804 155764
rect 195860 155708 384748 155764
rect 31892 155596 48748 155652
rect 48804 155596 93212 155652
rect 93268 155596 93278 155652
rect 117618 155596 117628 155652
rect 117684 155596 397404 155652
rect 397460 155596 429884 155652
rect 429940 155596 429950 155652
rect 31892 155428 31948 155596
rect 52882 155484 52892 155540
rect 52948 155484 112252 155540
rect 112308 155484 112318 155540
rect 114258 155484 114268 155540
rect 114324 155484 397628 155540
rect 397684 155484 418460 155540
rect 418516 155484 418526 155540
rect 6402 155372 6412 155428
rect 6468 155372 31948 155428
rect 82338 155372 82348 155428
rect 82404 155372 555548 155428
rect 555604 155372 555614 155428
rect 528294 155148 528332 155204
rect 528388 155148 528398 155204
rect 459442 154812 459452 154868
rect 459508 154812 460348 154868
rect 460404 154812 460414 154868
rect 481282 154812 481292 154868
rect 481348 154812 483196 154868
rect 483252 154812 483262 154868
rect 493042 154812 493052 154868
rect 493108 154812 494620 154868
rect 494676 154812 494686 154868
rect 220052 154700 231868 154756
rect 220052 154644 220108 154700
rect 231812 154644 231868 154700
rect 198146 154588 198156 154644
rect 198212 154588 220108 154644
rect 221676 154588 228676 154644
rect 231812 154588 260764 154644
rect 260820 154588 260830 154644
rect 262098 154588 262108 154644
rect 262164 154588 282212 154644
rect 9762 154476 9772 154532
rect 9828 154476 66332 154532
rect 66388 154476 66398 154532
rect 100930 154476 100940 154532
rect 100996 154476 191156 154532
rect 197250 154476 197260 154532
rect 197316 154476 197596 154532
rect 197652 154476 197662 154532
rect 206994 154476 207004 154532
rect 207060 154476 209356 154532
rect 209412 154476 209422 154532
rect 9874 154364 9884 154420
rect 9940 154364 51212 154420
rect 51268 154364 51278 154420
rect 131282 154364 131292 154420
rect 131348 154364 189644 154420
rect 189700 154364 189710 154420
rect 191100 154308 191156 154476
rect 195794 154364 195804 154420
rect 195860 154364 196252 154420
rect 196308 154364 206780 154420
rect 206836 154364 206846 154420
rect 221676 154308 221732 154588
rect 9986 154252 9996 154308
rect 10052 154252 47516 154308
rect 47572 154252 47852 154308
rect 47908 154252 47918 154308
rect 191100 154252 191884 154308
rect 191940 154252 198044 154308
rect 198100 154252 198110 154308
rect 209906 154252 209916 154308
rect 209972 154252 221732 154308
rect 228620 154308 228676 154588
rect 282156 154532 282212 154588
rect 287308 154588 319116 154644
rect 319172 154588 319182 154644
rect 342178 154588 342188 154644
rect 342244 154588 355348 154644
rect 287308 154532 287364 154588
rect 282156 154476 287364 154532
rect 355292 154532 355348 154588
rect 355292 154476 400316 154532
rect 400372 154476 400652 154532
rect 400708 154476 400718 154532
rect 230178 154364 230188 154420
rect 230244 154364 289884 154420
rect 289940 154364 289950 154420
rect 294242 154364 294252 154420
rect 294308 154364 316540 154420
rect 316596 154364 378700 154420
rect 378756 154364 379260 154420
rect 379316 154364 379326 154420
rect 379698 154364 379708 154420
rect 379764 154364 386428 154420
rect 386484 154364 386494 154420
rect 399074 154364 399084 154420
rect 399140 154364 464156 154420
rect 464212 154364 464222 154420
rect 518242 154364 518252 154420
rect 518308 154364 579852 154420
rect 579908 154364 579918 154420
rect 228620 154252 253708 154308
rect 253764 154252 253774 154308
rect 269266 154252 269276 154308
rect 269332 154252 282156 154308
rect 282212 154252 282222 154308
rect 304434 154252 304444 154308
rect 304500 154252 344652 154308
rect 344708 154252 344718 154308
rect 399522 154252 399532 154308
rect 399588 154252 456540 154308
rect 456596 154252 456606 154308
rect 8194 154140 8204 154196
rect 8260 154140 43708 154196
rect 43764 154140 44492 154196
rect 44548 154140 44558 154196
rect 203298 154140 203308 154196
rect 203364 154140 230300 154196
rect 230356 154140 230366 154196
rect 231812 154140 238700 154196
rect 238756 154140 238766 154196
rect 319106 154140 319116 154196
rect 319172 154140 342188 154196
rect 342244 154140 342254 154196
rect 343186 154140 343196 154196
rect 343252 154140 377132 154196
rect 377188 154140 377198 154196
rect 399186 154140 399196 154196
rect 399252 154140 437500 154196
rect 437556 154140 437566 154196
rect 231812 154084 231868 154140
rect 213042 154028 213052 154084
rect 213108 154028 231868 154084
rect 238578 154028 238588 154084
rect 238644 154028 251804 154084
rect 251860 154028 251870 154084
rect 270386 154028 270396 154084
rect 270452 154028 547708 154084
rect 547764 154028 547774 154084
rect 110002 153916 110012 153972
rect 110068 153916 131292 153972
rect 131348 153916 131358 153972
rect 168018 153916 168028 153972
rect 168084 153916 184604 153972
rect 184660 153916 184670 153972
rect 205650 153916 205660 153972
rect 205716 153916 211708 153972
rect 211764 153916 211774 153972
rect 215058 153916 215068 153972
rect 215124 153916 263788 153972
rect 263844 153916 263854 153972
rect 343298 153916 343308 153972
rect 343364 153916 378812 153972
rect 378868 153916 378878 153972
rect 107426 153804 107436 153860
rect 107492 153804 127484 153860
rect 127540 153804 127550 153860
rect 127698 153804 127708 153860
rect 127764 153804 262108 153860
rect 262164 153804 262174 153860
rect 278450 153804 278460 153860
rect 278516 153804 283388 153860
rect 283444 153804 283454 153860
rect 359538 153804 359548 153860
rect 359604 153804 399644 153860
rect 399700 153804 399710 153860
rect 99138 153692 99148 153748
rect 99204 153692 193900 153748
rect 193956 153692 193966 153748
rect 197026 153692 197036 153748
rect 197092 153692 506044 153748
rect 506100 153692 506110 153748
rect 519026 153692 519036 153748
rect 519092 153692 578060 153748
rect 578116 153692 578126 153748
rect 195682 153580 195692 153636
rect 195748 153580 197820 153636
rect 197876 153580 228956 153636
rect 229012 153580 229022 153636
rect 196242 153356 196252 153412
rect 196308 153356 317212 153412
rect 317268 153356 317278 153412
rect 84018 153244 84028 153300
rect 84084 153244 362796 153300
rect 362852 153244 362862 153300
rect 199154 153132 199164 153188
rect 199220 153132 215124 153188
rect 197250 153020 197260 153076
rect 197316 153020 201180 153076
rect 201236 153020 201246 153076
rect 193218 152908 193228 152964
rect 193284 152908 204988 152964
rect 205044 152908 205054 152964
rect 215068 152852 215124 153132
rect 7746 152796 7756 152852
rect 7812 152796 74172 152852
rect 74228 152796 74238 152852
rect 198034 152796 198044 152852
rect 198100 152796 205660 152852
rect 205716 152796 205726 152852
rect 215068 152796 247996 152852
rect 248052 152796 248062 152852
rect 253698 152796 253708 152852
rect 253764 152796 263228 152852
rect 263284 152796 263294 152852
rect 263890 152796 263900 152852
rect 263956 152796 532700 152852
rect 532756 152796 532766 152852
rect 201170 152684 201180 152740
rect 201236 152684 223356 152740
rect 223412 152684 223422 152740
rect 223794 152684 223804 152740
rect 223860 152684 253820 152740
rect 253876 152684 253886 152740
rect 260754 152684 260764 152740
rect 260820 152684 359548 152740
rect 359604 152684 359614 152740
rect 362786 152684 362796 152740
rect 362852 152684 559468 152740
rect 559524 152684 559534 152740
rect 189410 152572 189420 152628
rect 189476 152572 215068 152628
rect 215124 152572 215134 152628
rect 216738 152572 216748 152628
rect 216804 152572 244188 152628
rect 244244 152572 244254 152628
rect 253698 152572 253708 152628
rect 253764 152572 267036 152628
rect 267092 152572 267102 152628
rect 324146 152572 324156 152628
rect 324212 152572 332668 152628
rect 332724 152572 332734 152628
rect 378914 152572 378924 152628
rect 378980 152572 379708 152628
rect 379764 152572 379774 152628
rect 408212 152572 433692 152628
rect 433748 152572 433758 152628
rect 503122 152572 503132 152628
rect 503188 152572 578172 152628
rect 578228 152572 578238 152628
rect 160402 152460 160412 152516
rect 160468 152460 197036 152516
rect 197092 152460 199724 152516
rect 199780 152460 255612 152516
rect 255668 152460 255678 152516
rect 283378 152460 283388 152516
rect 283444 152460 363356 152516
rect 363412 152460 363422 152516
rect 126018 152348 126028 152404
rect 126084 152348 198156 152404
rect 198212 152348 198222 152404
rect 198370 152348 198380 152404
rect 198436 152348 373660 152404
rect 373716 152348 373726 152404
rect 100818 152236 100828 152292
rect 100884 152236 193228 152292
rect 193284 152236 193294 152292
rect 196578 152236 196588 152292
rect 196644 152236 397964 152292
rect 398020 152236 398030 152292
rect 408212 152180 408268 152572
rect 119298 152124 119308 152180
rect 119364 152124 397740 152180
rect 397796 152124 408268 152180
rect 62962 152012 62972 152068
rect 63028 152012 100940 152068
rect 100996 152012 101006 152068
rect 110898 152012 110908 152068
rect 110964 152012 397852 152068
rect 397908 152012 397918 152068
rect 204978 151900 204988 151956
rect 205044 151900 225484 151956
rect 225540 151900 225550 151956
rect 591560 151704 593000 151928
rect 197698 151340 197708 151396
rect 197764 151340 208348 151396
rect 208292 151284 208348 151340
rect 199378 151228 199388 151284
rect 199444 151228 199948 151284
rect 200004 151228 200014 151284
rect 208292 151228 214228 151284
rect 214172 151172 214228 151228
rect 191426 151116 191436 151172
rect 191492 151116 192668 151172
rect 192724 151116 192734 151172
rect 195458 151116 195468 151172
rect 195524 151116 196364 151172
rect 196420 151116 209916 151172
rect 209972 151116 209982 151172
rect 214172 151116 216748 151172
rect 216804 151116 216814 151172
rect 223346 151116 223356 151172
rect 223412 151116 238588 151172
rect 238644 151116 238654 151172
rect 252018 151116 252028 151172
rect 252084 151116 315420 151172
rect 315476 151116 315486 151172
rect 317202 151116 317212 151172
rect 317268 151116 400204 151172
rect 400260 151116 475580 151172
rect 475636 151116 475646 151172
rect 496402 151116 496412 151172
rect 496468 151116 498428 151172
rect 498484 151116 579628 151172
rect 579684 151116 579694 151172
rect 197810 151004 197820 151060
rect 197876 151004 202524 151060
rect 202580 151004 202590 151060
rect 208292 151004 213948 151060
rect 214004 151004 214014 151060
rect 215058 151004 215068 151060
rect 215124 151004 228508 151060
rect 228564 151004 228574 151060
rect 238690 151004 238700 151060
rect 238756 151004 253708 151060
rect 253764 151004 253774 151060
rect 398066 151004 398076 151060
rect 398132 151004 426076 151060
rect 426132 151004 426142 151060
rect 208292 150948 208348 151004
rect 198034 150892 198044 150948
rect 198100 150892 208348 150948
rect 209346 150892 209356 150948
rect 209412 150892 225260 150948
rect 225316 150892 225326 150948
rect 225474 150892 225484 150948
rect 225540 150892 238812 150948
rect 238868 150892 238878 150948
rect 206882 150780 206892 150836
rect 206948 150780 214956 150836
rect 215012 150780 215022 150836
rect 53778 150556 53788 150612
rect 53844 150556 203308 150612
rect 203364 150556 203374 150612
rect 363346 150556 363356 150612
rect 363412 150556 378924 150612
rect 378980 150556 378990 150612
rect 78978 150444 78988 150500
rect 79044 150444 544124 150500
rect 544180 150444 544190 150500
rect 9650 150332 9660 150388
rect 9716 150332 43820 150388
rect 43876 150332 81788 150388
rect 81844 150332 81854 150388
rect 156258 150332 156268 150388
rect 156324 150332 199388 150388
rect 199444 150332 199454 150388
rect 140242 149660 140252 149716
rect 140308 149660 195692 149716
rect 195748 149660 195758 149716
rect 89058 149548 89068 149604
rect 89124 149548 191436 149604
rect 191492 149548 191502 149604
rect -960 149240 480 149464
rect 134418 149436 134428 149492
rect 134484 149436 188636 149492
rect 188692 149436 188702 149492
rect 403218 149436 403228 149492
rect 403284 149436 589708 149492
rect 589764 149436 589774 149492
rect 400642 149324 400652 149380
rect 400708 149324 459452 149380
rect 459508 149324 459518 149380
rect 169698 148876 169708 148932
rect 169764 148876 198380 148932
rect 198436 148876 198446 148932
rect 31892 148764 45388 148820
rect 45444 148764 89068 148820
rect 89124 148764 89134 148820
rect 157938 148764 157948 148820
rect 158004 148764 188300 148820
rect 188356 148764 188366 148820
rect 31892 148708 31948 148764
rect 6626 148652 6636 148708
rect 6692 148652 31948 148708
rect 63858 148652 63868 148708
rect 63924 148652 197932 148708
rect 197988 148652 197998 148708
rect 192332 148204 194908 148260
rect 194964 148204 194974 148260
rect 109218 148092 109228 148148
rect 109284 148092 141036 148148
rect 141092 148092 141102 148148
rect 192332 148036 192388 148204
rect 136882 147980 136892 148036
rect 136948 147980 192388 148036
rect 194572 147980 196140 148036
rect 196196 147980 198716 148036
rect 198772 147980 198782 148036
rect 194572 147924 194628 147980
rect 135202 147868 135212 147924
rect 135268 147868 194628 147924
rect 194898 147868 194908 147924
rect 194964 147868 196364 147924
rect 196420 147868 197932 147924
rect 197988 147868 197998 147924
rect 146178 147756 146188 147812
rect 146244 147756 188972 147812
rect 189028 147756 189038 147812
rect 67172 147084 84812 147140
rect 84868 147084 84878 147140
rect 107538 147084 107548 147140
rect 107604 147084 134428 147140
rect 134484 147084 134494 147140
rect 67172 147028 67228 147084
rect 9874 146972 9884 147028
rect 9940 146972 65548 147028
rect 65604 146972 67228 147028
rect 73042 146972 73052 147028
rect 73108 146972 149548 147028
rect 149604 146972 149614 147028
rect 148642 146412 148652 146468
rect 148708 146412 196252 146468
rect 196308 146412 198044 146468
rect 198100 146412 198110 146468
rect 142034 146300 142044 146356
rect 142100 146300 197372 146356
rect 197428 146300 197438 146356
rect 136994 146188 137004 146244
rect 137060 146188 199052 146244
rect 199108 146188 199118 146244
rect 75618 145516 75628 145572
rect 75684 145516 190764 145572
rect 190820 145516 190830 145572
rect 68898 145404 68908 145460
rect 68964 145404 188188 145460
rect 188244 145404 188254 145460
rect 21858 145292 21868 145348
rect 21924 145292 198828 145348
rect 198884 145292 198894 145348
rect 150322 144620 150332 144676
rect 150388 144620 198268 144676
rect 198324 144620 199164 144676
rect 199220 144620 199230 144676
rect 143714 144508 143724 144564
rect 143780 144508 199388 144564
rect 199444 144508 199454 144564
rect 59602 143836 59612 143892
rect 59668 143836 119420 143892
rect 119476 143836 119486 143892
rect 87378 143724 87388 143780
rect 87444 143724 158732 143780
rect 158788 143724 158798 143780
rect 29362 143612 29372 143668
rect 29428 143612 180572 143668
rect 180628 143612 180638 143668
rect 143602 142940 143612 142996
rect 143668 142940 198156 142996
rect 198212 142940 198828 142996
rect 198884 142940 198894 142996
rect 138562 142828 138572 142884
rect 138628 142828 197484 142884
rect 197540 142828 197550 142884
rect 112578 142156 112588 142212
rect 112644 142156 196588 142212
rect 196644 142156 196654 142212
rect 70578 142044 70588 142100
rect 70644 142044 197484 142100
rect 197540 142044 197550 142100
rect 67218 141932 67228 141988
rect 67284 141932 197148 141988
rect 197204 141932 197214 141988
rect 591560 140616 593000 140840
rect 50418 140252 50428 140308
rect 50484 140252 116732 140308
rect 116788 140252 116798 140308
rect 159618 140252 159628 140308
rect 159684 140252 189196 140308
rect 189252 140252 189262 140308
rect 107314 139356 107324 139412
rect 107380 139356 107660 139412
rect 107716 139356 107726 139412
rect 125972 139356 137788 139412
rect 137844 139356 188524 139412
rect 188580 139356 188590 139412
rect 104962 139020 104972 139076
rect 105028 139020 122668 139076
rect 122724 139020 122734 139076
rect 125972 138964 126028 139356
rect 107650 138908 107660 138964
rect 107716 138908 126028 138964
rect 122658 138796 122668 138852
rect 122724 138796 196028 138852
rect 196084 138796 196094 138852
rect 77298 138684 77308 138740
rect 77364 138684 199388 138740
rect 199444 138684 199454 138740
rect -960 138376 480 138600
rect 26898 138572 26908 138628
rect 26964 138572 196252 138628
rect 196308 138572 196318 138628
rect 517346 138572 517356 138628
rect 517412 138572 535948 138628
rect 536004 138572 536014 138628
rect 47058 137788 47068 137844
rect 47124 137788 107324 137844
rect 107380 137788 107390 137844
rect 141026 137676 141036 137732
rect 141092 137676 188412 137732
rect 188468 137676 188478 137732
rect 131058 137004 131068 137060
rect 131124 137004 195804 137060
rect 195860 137004 195870 137060
rect 47842 136892 47852 136948
rect 47908 136892 141932 136948
rect 141988 136892 141998 136948
rect 141922 136444 141932 136500
rect 141988 136444 143612 136500
rect 143668 136444 143678 136500
rect 71362 135996 71372 136052
rect 71428 135996 139468 136052
rect 139524 135996 140252 136052
rect 140308 135996 140318 136052
rect 27682 135212 27692 135268
rect 27748 135212 135324 135268
rect 135380 135212 135390 135268
rect 66322 133644 66332 133700
rect 66388 133644 148876 133700
rect 148932 133644 148942 133700
rect 36978 133532 36988 133588
rect 37044 133532 197036 133588
rect 197092 133532 197102 133588
rect 37762 132636 37772 132692
rect 37828 132636 137788 132692
rect 137844 132636 138572 132692
rect 138628 132636 138638 132692
rect 59714 131852 59724 131908
rect 59780 131852 145292 131908
rect 145348 131852 145358 131908
rect 101042 131180 101052 131236
rect 101108 131180 197484 131236
rect 197540 131180 197550 131236
rect 96002 131068 96012 131124
rect 96068 131068 199276 131124
rect 199332 131068 199342 131124
rect 69682 130956 69692 131012
rect 69748 130956 149772 131012
rect 149828 130956 150332 131012
rect 150388 130956 150398 131012
rect 86706 130172 86716 130228
rect 86772 130172 153804 130228
rect 153860 130172 153870 130228
rect 591560 129528 593000 129752
rect 27458 129388 27468 129444
rect 27524 129388 188972 129444
rect 189028 129388 189038 129444
rect 44482 129276 44492 129332
rect 44548 129276 141148 129332
rect 141204 129276 142044 129332
rect 142100 129276 142110 129332
rect 173012 129276 198268 129332
rect 198324 129276 199052 129332
rect 199108 129276 199118 129332
rect 173012 129220 173068 129276
rect 104178 129164 104188 129220
rect 104244 129164 105532 129220
rect 105588 129164 173068 129220
rect 63074 128492 63084 128548
rect 63140 128492 147868 128548
rect 147924 128492 147934 128548
rect 171378 128492 171388 128548
rect 171444 128492 191548 128548
rect 191604 128492 191614 128548
rect -960 127540 480 127736
rect 28802 127708 28812 127764
rect 28868 127708 194012 127764
rect 194068 127708 194078 127764
rect 46162 127596 46172 127652
rect 46228 127596 135212 127652
rect 135268 127596 135278 127652
rect -960 127512 532 127540
rect 392 127484 532 127512
rect 476 127428 532 127484
rect 364 127372 532 127428
rect 364 126084 420 127372
rect 47170 126924 47180 126980
rect 47236 126924 105532 126980
rect 105588 126924 105598 126980
rect 94098 126812 94108 126868
rect 94164 126812 173852 126868
rect 173908 126812 173918 126868
rect 120978 126252 120988 126308
rect 121044 126252 193004 126308
rect 193060 126252 193070 126308
rect 85698 126140 85708 126196
rect 85764 126140 192668 126196
rect 192724 126140 192734 126196
rect 364 126028 11788 126084
rect 11844 126028 11854 126084
rect 34178 126028 34188 126084
rect 34244 126028 197484 126084
rect 197540 126028 197550 126084
rect 89058 125916 89068 125972
rect 89124 125916 90636 125972
rect 90692 125916 189756 125972
rect 189812 125916 189822 125972
rect 90066 125244 90076 125300
rect 90132 125244 162092 125300
rect 162148 125244 162158 125300
rect 91410 125132 91420 125188
rect 91476 125132 163772 125188
rect 163828 125132 163838 125188
rect 173012 124572 194516 124628
rect 173012 124516 173068 124572
rect 153794 124460 153804 124516
rect 153860 124460 173068 124516
rect 188860 124460 192892 124516
rect 192948 124460 192958 124516
rect 188860 124404 188916 124460
rect 194460 124404 194516 124572
rect 122322 124348 122332 124404
rect 122388 124348 188916 124404
rect 189746 124348 189756 124404
rect 189812 124348 190652 124404
rect 190708 124348 190718 124404
rect 194450 124348 194460 124404
rect 194516 124348 195804 124404
rect 195860 124348 195870 124404
rect 51202 124236 51212 124292
rect 51268 124236 143836 124292
rect 143892 124236 143902 124292
rect 107426 124124 107436 124180
rect 107492 124124 190876 124180
rect 190932 124124 190942 124180
rect 44370 123564 44380 123620
rect 44436 123564 89068 123620
rect 89124 123564 89134 123620
rect 91522 123564 91532 123620
rect 91588 123564 151900 123620
rect 151956 123564 151966 123620
rect 89170 123452 89180 123508
rect 89236 123452 153692 123508
rect 153748 123452 153758 123508
rect 155922 123452 155932 123508
rect 155988 123452 175532 123508
rect 175588 123452 175598 123508
rect 145282 122780 145292 122836
rect 145348 122780 146524 122836
rect 146580 122780 199164 122836
rect 199220 122780 199230 122836
rect 104850 122668 104860 122724
rect 104916 122668 107436 122724
rect 107492 122668 107502 122724
rect 125010 122668 125020 122724
rect 125076 122668 195804 122724
rect 195860 122668 195870 122724
rect 41122 122556 41132 122612
rect 41188 122556 137116 122612
rect 137172 122556 137182 122612
rect 194898 122556 194908 122612
rect 194964 122556 197260 122612
rect 197316 122556 197326 122612
rect 107314 121884 107324 121940
rect 107380 121884 191660 121940
rect 191716 121884 191726 121940
rect 57810 121772 57820 121828
rect 57876 121772 194684 121828
rect 194740 121772 194750 121828
rect 173012 121324 194908 121380
rect 194964 121324 196028 121380
rect 196084 121324 196094 121380
rect 173012 121268 173068 121324
rect 147858 121212 147868 121268
rect 147924 121212 173068 121268
rect 191314 121212 191324 121268
rect 191380 121212 191660 121268
rect 191716 121212 191726 121268
rect 33618 121100 33628 121156
rect 33684 121100 194684 121156
rect 194740 121100 194750 121156
rect 30930 120988 30940 121044
rect 30996 120988 199388 121044
rect 199444 120988 199454 121044
rect 47058 120652 47068 120708
rect 47124 120652 47740 120708
rect 47796 120652 47806 120708
rect 100818 120652 100828 120708
rect 100884 120652 101500 120708
rect 101556 120652 101566 120708
rect 86482 120316 86492 120372
rect 86548 120316 145180 120372
rect 145236 120316 145246 120372
rect 92754 120204 92764 120260
rect 92820 120204 167132 120260
rect 167188 120204 167198 120260
rect 22642 120092 22652 120148
rect 22708 120092 133084 120148
rect 133140 120092 133150 120148
rect 194786 119980 194796 120036
rect 194852 119980 195468 120036
rect 195524 119980 195534 120036
rect 151890 119644 151900 119700
rect 151956 119644 194796 119700
rect 194852 119644 194862 119700
rect 145170 119532 145180 119588
rect 145236 119532 197708 119588
rect 197764 119532 197774 119588
rect 116946 119420 116956 119476
rect 117012 119420 197932 119476
rect 197988 119420 197998 119476
rect 25554 119308 25564 119364
rect 25620 119308 193116 119364
rect 193172 119308 193182 119364
rect 24210 119196 24220 119252
rect 24276 119196 29372 119252
rect 29428 119196 29438 119252
rect 41682 119196 41692 119252
rect 41748 119196 45388 119252
rect 45444 119196 45454 119252
rect 67218 119196 67228 119252
rect 67284 119196 73052 119252
rect 73108 119196 73118 119252
rect 103506 119196 103516 119252
rect 103572 119196 104972 119252
rect 105028 119196 105038 119252
rect 134418 119196 134428 119252
rect 134484 119196 135324 119252
rect 135380 119196 148652 119252
rect 148708 119196 148718 119252
rect 148866 119196 148876 119252
rect 148932 119196 160412 119252
rect 160468 119196 160478 119252
rect 106194 119084 106204 119140
rect 106260 119084 110012 119140
rect 110068 119084 110078 119140
rect 133074 119084 133084 119140
rect 133140 119084 136892 119140
rect 136948 119084 136958 119140
rect 49746 118972 49756 119028
rect 49812 118972 52892 119028
rect 52948 118972 52958 119028
rect 178770 118748 178780 118804
rect 178836 118748 195692 118804
rect 195748 118748 195758 118804
rect 43026 118636 43036 118692
rect 43092 118636 48748 118692
rect 48804 118636 48814 118692
rect 53778 118636 53788 118692
rect 53844 118636 59612 118692
rect 59668 118636 59678 118692
rect 173394 118636 173404 118692
rect 173460 118636 194572 118692
rect 194628 118636 194638 118692
rect 45714 118524 45724 118580
rect 45780 118524 62972 118580
rect 63028 118524 63038 118580
rect 165330 118524 165340 118580
rect 165396 118524 189084 118580
rect 189140 118524 189150 118580
rect 40338 118412 40348 118468
rect 40404 118412 65548 118468
rect 65604 118412 65614 118468
rect 80658 118412 80668 118468
rect 80724 118412 197820 118468
rect 197876 118412 197886 118468
rect 591560 118440 593000 118664
rect 87378 118300 87388 118356
rect 87444 118300 89180 118356
rect 89236 118300 89246 118356
rect 38994 118076 39004 118132
rect 39060 118076 43820 118132
rect 43876 118076 43886 118132
rect 154578 118076 154588 118132
rect 154644 118076 194124 118132
rect 194180 118076 194190 118132
rect 127698 117964 127708 118020
rect 127764 117964 189308 118020
rect 189364 117964 189374 118020
rect 95442 117852 95452 117908
rect 95508 117852 176876 117908
rect 176932 117852 176942 117908
rect 115602 117740 115612 117796
rect 115668 117740 199052 117796
rect 199108 117740 199118 117796
rect 52434 117628 52444 117684
rect 52500 117628 193900 117684
rect 193956 117628 193966 117684
rect -960 116676 480 116872
rect 176866 116732 176876 116788
rect 176932 116732 194572 116788
rect 194628 116732 194638 116788
rect -960 116648 10892 116676
rect 392 116620 10892 116648
rect 10948 116620 10958 116676
rect 168018 116396 168028 116452
rect 168084 116396 195468 116452
rect 195524 116396 195534 116452
rect 130386 116284 130396 116340
rect 130452 116284 195916 116340
rect 195972 116284 195982 116340
rect 82002 116172 82012 116228
rect 82068 116172 197820 116228
rect 197876 116172 197886 116228
rect 66546 116060 66556 116116
rect 66612 116060 196252 116116
rect 196308 116060 196318 116116
rect 36866 115948 36876 116004
rect 36932 115948 195692 116004
rect 195748 115948 195758 116004
rect 19506 114380 19516 114436
rect 19572 114380 21672 114436
rect 19282 113036 19292 113092
rect 19348 113036 21672 113092
rect 20066 111692 20076 111748
rect 20132 111692 21672 111748
rect 19954 110348 19964 110404
rect 20020 110348 21672 110404
rect 19842 109004 19852 109060
rect 19908 109004 21672 109060
rect 19394 107660 19404 107716
rect 19460 107660 21672 107716
rect 591560 107352 593000 107576
rect 20178 106316 20188 106372
rect 20244 106316 21672 106372
rect -960 105784 480 106008
rect 20402 104972 20412 105028
rect 20468 104972 21672 105028
rect 198034 104076 198044 104132
rect 198100 104076 198268 104132
rect 198324 104076 198334 104132
rect 395602 104076 395612 104132
rect 395668 104076 396396 104132
rect 396452 104076 481292 104132
rect 481348 104076 481358 104132
rect 20290 103628 20300 103684
rect 20356 103628 21672 103684
rect 400642 102396 400652 102452
rect 400708 102396 493052 102452
rect 493108 102396 493118 102452
rect 16258 102284 16268 102340
rect 16324 102284 21672 102340
rect 517346 101500 517356 101556
rect 517412 101500 520072 101556
rect 19954 100940 19964 100996
rect 20020 100940 21672 100996
rect 516562 100828 516572 100884
rect 516628 100828 517356 100884
rect 517412 100828 517422 100884
rect 19506 99596 19516 99652
rect 19572 99596 21672 99652
rect 19730 98252 19740 98308
rect 19796 98252 21672 98308
rect 19618 96908 19628 96964
rect 19684 96908 21672 96964
rect 591560 96264 593000 96488
rect 19170 95564 19180 95620
rect 19236 95564 21672 95620
rect -960 94948 480 95144
rect -960 94920 532 94948
rect 392 94892 532 94920
rect 476 94836 532 94892
rect 364 94780 532 94836
rect 364 94164 420 94780
rect 19730 94220 19740 94276
rect 19796 94220 21672 94276
rect 364 94108 19404 94164
rect 19460 94108 19470 94164
rect 16146 92876 16156 92932
rect 16212 92876 21672 92932
rect 20066 91532 20076 91588
rect 20132 91532 21672 91588
rect 19618 90188 19628 90244
rect 19684 90188 21672 90244
rect 19170 88844 19180 88900
rect 19236 88844 21672 88900
rect 16034 87500 16044 87556
rect 16100 87500 21672 87556
rect 22194 86156 22204 86212
rect 22260 86156 22270 86212
rect 591560 85176 593000 85400
rect 519026 84924 519036 84980
rect 519092 84924 520072 84980
rect 18386 84812 18396 84868
rect 18452 84812 21672 84868
rect -960 84056 480 84280
rect 569884 84196 569940 84952
rect 569884 84140 572908 84196
rect 572852 84084 572908 84140
rect 572852 84028 589820 84084
rect 589876 84028 589886 84084
rect 20290 83468 20300 83524
rect 20356 83468 21672 83524
rect 22306 82124 22316 82180
rect 22372 82124 22382 82180
rect 20178 80780 20188 80836
rect 20244 80780 21672 80836
rect 21644 79044 21700 79464
rect 4946 78988 4956 79044
rect 5012 78988 21700 79044
rect 21644 77364 21700 78120
rect 11666 77308 11676 77364
rect 11732 77308 21700 77364
rect 21644 75684 21700 76776
rect 3266 75628 3276 75684
rect 3332 75628 21700 75684
rect 21644 74452 21700 75432
rect 9986 74396 9996 74452
rect 10052 74396 21700 74452
rect 8372 74060 21672 74116
rect 591560 74088 593000 74312
rect 8372 74004 8428 74060
rect 6514 73948 6524 74004
rect 6580 73948 8428 74004
rect 19618 73612 19628 73668
rect 19684 73612 22092 73668
rect 22148 73612 22158 73668
rect 19954 73500 19964 73556
rect 20020 73500 21980 73556
rect 22036 73500 22046 73556
rect -960 73220 480 73416
rect 20066 73388 20076 73444
rect 20132 73388 22092 73444
rect 22148 73388 22158 73444
rect -960 73192 532 73220
rect 392 73164 532 73192
rect 476 73108 532 73164
rect 364 73052 532 73108
rect 364 72324 420 73052
rect 19842 72492 19852 72548
rect 19908 72492 20972 72548
rect 21028 72492 21038 72548
rect 21644 72436 21700 72744
rect 6626 72380 6636 72436
rect 6692 72380 21700 72436
rect 364 72268 21868 72324
rect 21924 72268 21934 72324
rect 18162 71372 18172 71428
rect 18228 71372 21672 71428
rect 8372 71148 21028 71204
rect 8372 70868 8428 71148
rect 4386 70812 4396 70868
rect 4452 70812 8428 70868
rect 15092 70924 18116 70980
rect 18274 70924 18284 70980
rect 18340 70924 19516 70980
rect 19572 70924 19582 70980
rect 15092 70756 15148 70924
rect 18060 70868 18116 70924
rect 20972 70868 21028 71148
rect 18060 70812 19572 70868
rect 20972 70812 31948 70868
rect 19516 70756 19572 70812
rect 31892 70756 31948 70812
rect 4834 70700 4844 70756
rect 4900 70700 15148 70756
rect 18162 70700 18172 70756
rect 18228 70700 19292 70756
rect 19348 70700 19358 70756
rect 19516 70700 21812 70756
rect 22082 70700 22092 70756
rect 22148 70700 23324 70756
rect 23380 70700 23390 70756
rect 31892 70700 47404 70756
rect 47460 70700 47470 70756
rect 11554 70588 11564 70644
rect 11620 70588 18172 70644
rect 18228 70588 18238 70644
rect 21756 70532 21812 70700
rect 21970 70588 21980 70644
rect 22036 70588 22876 70644
rect 22932 70588 22942 70644
rect 21756 70476 21980 70532
rect 22036 70476 22046 70532
rect 22194 70476 22204 70532
rect 22260 70476 23100 70532
rect 23156 70476 23166 70532
rect 20178 70140 20188 70196
rect 20244 70140 64092 70196
rect 64148 70140 64158 70196
rect 20402 70028 20412 70084
rect 20468 70028 64540 70084
rect 64596 70028 64606 70084
rect 19170 69916 19180 69972
rect 19236 69916 64876 69972
rect 64932 69916 64942 69972
rect 20066 69804 20076 69860
rect 20132 69804 64204 69860
rect 64260 69804 64270 69860
rect 19730 69692 19740 69748
rect 19796 69692 63980 69748
rect 64036 69692 64046 69748
rect 21858 69356 21868 69412
rect 21924 69356 33292 69412
rect 33348 69356 33358 69412
rect 19394 69132 19404 69188
rect 19460 69132 30940 69188
rect 30996 69132 31006 69188
rect 31154 69132 31164 69188
rect 31220 69132 40348 69188
rect 40404 69132 40414 69188
rect 77970 69132 77980 69188
rect 78036 69132 190876 69188
rect 190932 69132 190942 69188
rect 10098 69020 10108 69076
rect 10164 69020 35644 69076
rect 35700 69020 35710 69076
rect 75618 69020 75628 69076
rect 75684 69020 192332 69076
rect 192388 69020 192398 69076
rect 4722 68908 4732 68964
rect 4788 68908 45052 68964
rect 45108 68908 45118 68964
rect 66210 68908 66220 68964
rect 66276 68908 190652 68964
rect 190708 68908 190718 68964
rect 21970 68796 21980 68852
rect 22036 68796 31164 68852
rect 31220 68796 31230 68852
rect 68562 68796 68572 68852
rect 68628 68796 197372 68852
rect 197428 68796 197438 68852
rect 80322 68684 80332 68740
rect 80388 68684 197596 68740
rect 197652 68684 197662 68740
rect 20290 68572 20300 68628
rect 20356 68572 31948 68628
rect 36978 68572 36988 68628
rect 37044 68572 37324 68628
rect 37380 68572 37390 68628
rect 41990 68572 42028 68628
rect 42084 68572 42094 68628
rect 48738 68572 48748 68628
rect 48804 68572 49084 68628
rect 49140 68572 49150 68628
rect 52070 68572 52108 68628
rect 52164 68572 52174 68628
rect 53750 68572 53788 68628
rect 53844 68572 53854 68628
rect 55458 68572 55468 68628
rect 55524 68572 56140 68628
rect 56196 68572 56206 68628
rect 58604 68572 64316 68628
rect 64372 68572 64382 68628
rect 89730 68572 89740 68628
rect 89796 68572 192556 68628
rect 192612 68572 192622 68628
rect 31892 68516 31948 68572
rect 58604 68516 58660 68572
rect 19506 68460 19516 68516
rect 19572 68460 28868 68516
rect 31892 68460 58660 68516
rect 58790 68460 58828 68516
rect 58884 68460 58894 68516
rect 60722 68460 60732 68516
rect 60788 68460 60844 68516
rect 60900 68460 60910 68516
rect 28812 68404 28868 68460
rect 25526 68348 25564 68404
rect 25620 68348 25630 68404
rect 28550 68348 28588 68404
rect 28644 68348 28654 68404
rect 28812 68348 61348 68404
rect 61292 68264 61348 68348
rect 520044 67284 520100 68376
rect 388882 67228 388892 67284
rect 388948 67228 520100 67284
rect 63858 67116 63868 67172
rect 63924 67116 189868 67172
rect 189924 67116 189934 67172
rect 73266 67004 73276 67060
rect 73332 67004 192444 67060
rect 192500 67004 192510 67060
rect 10882 66892 10892 66948
rect 10948 66892 12068 66948
rect 87378 66892 87388 66948
rect 87444 66892 194236 66948
rect 194292 66892 194302 66948
rect 12012 66584 12068 66892
rect 61516 66164 61572 66808
rect 85026 66780 85036 66836
rect 85092 66780 188972 66836
rect 189028 66780 189038 66836
rect 61506 66108 61516 66164
rect 61572 66108 61582 66164
rect 146178 65884 146188 65940
rect 146244 65884 147980 65940
rect 148036 65884 148046 65940
rect 96786 65548 96796 65604
rect 96852 65548 98252 65604
rect 98308 65548 98318 65604
rect 110898 65548 110908 65604
rect 110964 65548 113372 65604
rect 113428 65548 113438 65604
rect 115602 65548 115612 65604
rect 115668 65548 116732 65604
rect 116788 65548 116798 65604
rect 162642 65548 162652 65604
rect 162708 65548 163772 65604
rect 163828 65548 163838 65604
rect 70914 65436 70924 65492
rect 70980 65436 194012 65492
rect 194068 65436 194078 65492
rect 61516 64708 61572 65352
rect 164994 64764 165004 64820
rect 165060 64764 180572 64820
rect 180628 64764 180638 64820
rect 61506 64652 61516 64708
rect 61572 64652 61582 64708
rect 147970 64652 147980 64708
rect 148036 64652 154588 64708
rect 154644 64652 154654 64708
rect 155586 64652 155596 64708
rect 155652 64652 171500 64708
rect 171556 64652 171566 64708
rect 61880 63868 64764 63924
rect 64820 63868 64830 63924
rect 82674 63756 82684 63812
rect 82740 63756 194348 63812
rect 194404 63756 194414 63812
rect 113250 62972 113260 63028
rect 113316 62972 162092 63028
rect 162148 62972 162158 63028
rect 172050 62972 172060 63028
rect 172116 62972 191548 63028
rect 191604 62972 191614 63028
rect 591560 63000 593000 63224
rect 392 62552 10108 62580
rect -960 62524 10108 62552
rect 10164 62524 10174 62580
rect -960 62328 480 62524
rect 61880 62412 64652 62468
rect 64708 62412 64718 62468
rect 129714 61292 129724 61348
rect 129780 61292 190764 61348
rect 190820 61292 190830 61348
rect 61880 60956 65100 61012
rect 65156 60956 65166 61012
rect 11778 60508 11788 60564
rect 11844 60508 12068 60564
rect 12012 60424 12068 60508
rect 61880 59500 64092 59556
rect 64148 59500 64158 59556
rect 61880 58044 64428 58100
rect 64484 58044 64494 58100
rect 61880 56588 64316 56644
rect 64372 56588 64382 56644
rect 61880 55132 64988 55188
rect 65044 55132 65054 55188
rect 9314 54796 9324 54852
rect 9380 54796 12068 54852
rect 12012 54264 12068 54796
rect 61880 53676 64540 53732
rect 64596 53676 64606 53732
rect 61880 52220 64316 52276
rect 64372 52220 64382 52276
rect 591560 51912 593000 52136
rect -960 51464 480 51688
rect 61880 50764 63980 50820
rect 64036 50764 64046 50820
rect 61880 49308 64540 49364
rect 64596 49308 64606 49364
rect 12012 47124 12068 48104
rect 61880 47852 64428 47908
rect 64484 47852 64494 47908
rect 18 47068 28 47124
rect 84 47068 12068 47124
rect 61880 46396 64316 46452
rect 64372 46396 64382 46452
rect 61516 44324 61572 44968
rect 61506 44268 61516 44324
rect 61572 44268 61582 44324
rect 61880 43484 64204 43540
rect 64260 43484 64270 43540
rect 61880 42028 63868 42084
rect 63924 42028 63934 42084
rect -960 40628 480 40824
rect -960 40600 10892 40628
rect 392 40572 10892 40600
rect 10948 40572 10958 40628
rect 12012 40516 12068 41944
rect 591560 40824 593000 41048
rect 61880 40572 64876 40628
rect 64932 40572 64942 40628
rect 6066 40460 6076 40516
rect 6132 40460 12068 40516
rect 61880 39116 62188 39172
rect 62244 39116 62254 39172
rect 61516 37044 61572 37688
rect 61506 36988 61516 37044
rect 61572 36988 61582 37044
rect 12012 35364 12068 35784
rect 61852 35588 61908 36232
rect 61852 35532 61964 35588
rect 62020 35532 62030 35588
rect 2594 35308 2604 35364
rect 2660 35308 12068 35364
rect 61730 34748 61740 34804
rect 61796 34748 61806 34804
rect 61880 33292 64092 33348
rect 64148 33292 64158 33348
rect 61880 31836 62300 31892
rect 62356 31836 62366 31892
rect 61880 30380 63868 30436
rect 63924 30380 63934 30436
rect 9202 30156 9212 30212
rect 9268 30156 12068 30212
rect -960 29764 480 29960
rect -960 29736 11004 29764
rect 392 29708 11004 29736
rect 11060 29708 11070 29764
rect 12012 29624 12068 30156
rect 591560 29736 593000 29960
rect 61880 28924 64204 28980
rect 64260 28924 64270 28980
rect 107538 27692 107548 27748
rect 107604 27692 157052 27748
rect 157108 27692 157118 27748
rect 61880 27468 63980 27524
rect 64036 27468 64046 27524
rect 61926 27132 61964 27188
rect 62020 27132 62030 27188
rect 152898 26796 152908 26852
rect 152964 26796 163996 26852
rect 164052 26796 164062 26852
rect 61880 26012 63980 26068
rect 64036 26012 64046 26068
rect 163762 26012 163772 26068
rect 163828 26012 178108 26068
rect 178164 26012 178174 26068
rect 61628 23940 61684 24584
rect 100818 24332 100828 24388
rect 100884 24332 152908 24388
rect 152964 24332 152974 24388
rect 61618 23884 61628 23940
rect 61684 23884 61694 23940
rect 12012 21924 12068 23464
rect 61516 22484 61572 23128
rect 147858 22876 147868 22932
rect 147924 22876 158060 22932
rect 158116 22876 158126 22932
rect 102498 22652 102508 22708
rect 102564 22652 145292 22708
rect 145348 22652 145358 22708
rect 157938 22652 157948 22708
rect 158004 22652 171388 22708
rect 171444 22652 171454 22708
rect 61506 22428 61516 22484
rect 61572 22428 61582 22484
rect 2482 21868 2492 21924
rect 2548 21868 12068 21924
rect 61842 21644 61852 21700
rect 61908 21644 61918 21700
rect 4946 21420 4956 21476
rect 5012 21420 63868 21476
rect 63924 21420 63934 21476
rect 6514 21308 6524 21364
rect 6580 21308 61628 21364
rect 61684 21308 61694 21364
rect 9986 21196 9996 21252
rect 10052 21196 63980 21252
rect 64036 21196 64046 21252
rect 8306 21084 8316 21140
rect 8372 21084 60732 21140
rect 60788 21084 60798 21140
rect 99138 21084 99148 21140
rect 99204 21084 148652 21140
rect 148708 21084 148718 21140
rect 22642 20972 22652 21028
rect 22708 20972 60844 21028
rect 60900 20972 60910 21028
rect 119298 20972 119308 21028
rect 119364 20972 179788 21028
rect 179844 20972 179854 21028
rect 60610 20860 60620 20916
rect 60676 20860 61628 20916
rect 61684 20860 61694 20916
rect 11554 20188 11564 20244
rect 11620 20188 61852 20244
rect 61908 20188 61918 20244
rect 10994 20076 11004 20132
rect 11060 20076 25564 20132
rect 25620 20076 25630 20132
rect 6626 19964 6636 20020
rect 6692 19964 61516 20020
rect 61572 19964 61582 20020
rect 11666 19852 11676 19908
rect 11732 19852 64204 19908
rect 64260 19852 64270 19908
rect 7522 19740 7532 19796
rect 7588 19740 53788 19796
rect 53844 19740 53854 19796
rect 20290 19628 20300 19684
rect 20356 19628 60620 19684
rect 60676 19628 60686 19684
rect 23314 19516 23324 19572
rect 23380 19516 60620 19572
rect 60676 19516 60686 19572
rect 3266 19404 3276 19460
rect 3332 19404 63980 19460
rect 64036 19404 64046 19460
rect -960 18872 480 19096
rect 591560 18648 593000 18872
rect 14914 18508 14924 18564
rect 14980 18508 175532 18564
rect 175588 18508 175598 18564
rect 9986 18396 9996 18452
rect 10052 18396 58828 18452
rect 58884 18396 58894 18452
rect 19730 18284 19740 18340
rect 19796 18284 64316 18340
rect 64372 18284 64382 18340
rect 23090 18172 23100 18228
rect 23156 18172 64540 18228
rect 64596 18172 64606 18228
rect 22754 18060 22764 18116
rect 22820 18060 64092 18116
rect 64148 18060 64158 18116
rect 4610 17948 4620 18004
rect 4676 17948 42028 18004
rect 42084 17948 42094 18004
rect 53330 17612 53340 17668
rect 53396 17612 199276 17668
rect 199332 17612 199342 17668
rect 20402 17500 20412 17556
rect 20468 17500 23436 17556
rect 23492 17500 23502 17556
rect 42354 16828 42364 16884
rect 42420 16828 44716 16884
rect 44772 16828 44782 16884
rect 7634 16716 7644 16772
rect 7700 16716 55468 16772
rect 55524 16716 55534 16772
rect 19170 16604 19180 16660
rect 19236 16604 64428 16660
rect 64484 16604 64494 16660
rect 7858 16492 7868 16548
rect 7924 16492 52108 16548
rect 52164 16492 52174 16548
rect 19618 16380 19628 16436
rect 19684 16380 63868 16436
rect 63924 16380 63934 16436
rect 20178 16268 20188 16324
rect 20244 16268 62300 16324
rect 62356 16268 62366 16324
rect 10882 16156 10892 16212
rect 10948 16156 36988 16212
rect 37044 16156 37054 16212
rect 23426 15036 23436 15092
rect 23492 15036 131068 15092
rect 131124 15036 131628 15092
rect 131684 15036 131694 15092
rect 16258 14924 16268 14980
rect 16324 14924 64988 14980
rect 65044 14924 65054 14980
rect 16146 14812 16156 14868
rect 16212 14812 60732 14868
rect 60788 14812 60798 14868
rect 19954 14700 19964 14756
rect 20020 14700 64540 14756
rect 64596 14700 64606 14756
rect 18386 14588 18396 14644
rect 18452 14588 60508 14644
rect 60564 14588 60574 14644
rect 149538 14588 149548 14644
rect 149604 14588 160412 14644
rect 160468 14588 160478 14644
rect 22866 14476 22876 14532
rect 22932 14476 64764 14532
rect 64820 14476 64830 14532
rect 90738 14364 90748 14420
rect 90804 14364 140028 14420
rect 140084 14364 140094 14420
rect 131618 14252 131628 14308
rect 131684 14252 196588 14308
rect 196644 14252 196654 14308
rect 44706 13356 44716 13412
rect 44772 13356 173068 13412
rect 173124 13356 174636 13412
rect 174692 13356 174702 13412
rect 196130 13356 196140 13412
rect 196196 13356 198492 13412
rect 198548 13356 198558 13412
rect 18274 13244 18284 13300
rect 18340 13244 64316 13300
rect 64372 13244 64382 13300
rect 194450 13244 194460 13300
rect 194516 13244 198828 13300
rect 198884 13244 198894 13300
rect 19394 13132 19404 13188
rect 19460 13132 65100 13188
rect 65156 13132 65166 13188
rect 20962 13020 20972 13076
rect 21028 13020 64652 13076
rect 64708 13020 64718 13076
rect 18162 12908 18172 12964
rect 18228 12908 60396 12964
rect 60452 12908 60462 12964
rect 4162 12796 4172 12852
rect 4228 12796 48748 12852
rect 48804 12796 48814 12852
rect 159618 12796 159628 12852
rect 159684 12796 174748 12852
rect 174804 12796 174814 12852
rect 174626 12684 174636 12740
rect 174692 12684 194908 12740
rect 194964 12684 194974 12740
rect 58818 12572 58828 12628
rect 58884 12572 198604 12628
rect 198660 12572 198670 12628
rect 530898 12572 530908 12628
rect 530964 12572 567868 12628
rect 567924 12572 567934 12628
rect 169698 11116 169708 11172
rect 169764 11116 188860 11172
rect 188916 11116 188926 11172
rect 124338 11004 124348 11060
rect 124404 11004 170268 11060
rect 170324 11004 170334 11060
rect 47842 10892 47852 10948
rect 47908 10892 198940 10948
rect 198996 10892 199006 10948
rect 196018 10444 196028 10500
rect 196084 10444 203196 10500
rect 203252 10444 203262 10500
rect 196242 10332 196252 10388
rect 196308 10332 200172 10388
rect 200228 10332 200238 10388
rect 188962 10220 188972 10276
rect 189028 10220 198268 10276
rect 198324 10220 198334 10276
rect 16034 9996 16044 10052
rect 16100 9996 62188 10052
rect 62244 9996 62254 10052
rect 199266 9996 199276 10052
rect 199332 9996 518252 10052
rect 518308 9996 518318 10052
rect 194562 9884 194572 9940
rect 194628 9884 513212 9940
rect 513268 9884 513278 9940
rect 195794 9772 195804 9828
rect 195860 9772 399420 9828
rect 399476 9772 399486 9828
rect 177202 9660 177212 9716
rect 177268 9660 335580 9716
rect 335636 9660 335646 9716
rect 199490 9548 199500 9604
rect 199556 9548 205100 9604
rect 205156 9548 205166 9604
rect 116722 9324 116732 9380
rect 116788 9324 174300 9380
rect 174356 9324 174366 9380
rect 126018 9212 126028 9268
rect 126084 9212 191100 9268
rect 191156 9212 191166 9268
rect 197922 9212 197932 9268
rect 197988 9212 347788 9268
rect 347844 9212 347854 9268
rect 196242 8652 196252 8708
rect 196308 8652 213724 8708
rect 213780 8652 213790 8708
rect 350802 8652 350812 8708
rect 350868 8652 378476 8708
rect 378532 8652 378542 8708
rect 198482 8540 198492 8596
rect 198548 8540 217532 8596
rect 217588 8540 217598 8596
rect 320338 8540 320348 8596
rect 320404 8540 377356 8596
rect 377412 8540 377422 8596
rect 142818 8428 142828 8484
rect 142884 8428 151900 8484
rect 151956 8428 151966 8484
rect 198146 8428 198156 8484
rect 198212 8428 236572 8484
rect 236628 8428 236638 8484
rect 335570 8428 335580 8484
rect 335636 8428 516572 8484
rect 516628 8428 516638 8484
rect 4498 8316 4508 8372
rect 4564 8316 202300 8372
rect 202356 8316 202366 8372
rect 369842 8316 369852 8372
rect 369908 8316 379708 8372
rect 379764 8316 379774 8372
rect -960 8036 480 8232
rect 4274 8204 4284 8260
rect 4340 8204 206108 8260
rect 206164 8204 206174 8260
rect 327954 8204 327964 8260
rect 328020 8204 378140 8260
rect 378196 8204 378206 8260
rect 362226 8092 362236 8148
rect 362292 8092 386428 8148
rect 386484 8092 386494 8148
rect -960 8008 532 8036
rect 392 7980 532 8008
rect 136098 7980 136108 8036
rect 136164 7980 141820 8036
rect 141876 7980 141886 8036
rect 358418 7980 358428 8036
rect 358484 7980 383068 8036
rect 383124 7980 383134 8036
rect 476 7924 532 7980
rect 364 7868 532 7924
rect 134418 7868 134428 7924
rect 134484 7868 138460 7924
rect 138516 7868 138526 7924
rect 193890 7868 193900 7924
rect 193956 7868 308924 7924
rect 308980 7868 308990 7924
rect 346994 7868 347004 7924
rect 347060 7868 378364 7924
rect 378420 7868 378430 7924
rect 364 6804 420 7868
rect 199154 7756 199164 7812
rect 199220 7756 247996 7812
rect 248052 7756 248062 7812
rect 354610 7756 354620 7812
rect 354676 7756 378588 7812
rect 378644 7756 378654 7812
rect 105858 7644 105868 7700
rect 105924 7644 134428 7700
rect 134484 7644 134494 7700
rect 166338 7644 166348 7700
rect 166404 7644 182364 7700
rect 182420 7644 182430 7700
rect 117618 7532 117628 7588
rect 117684 7532 177660 7588
rect 177716 7532 177726 7588
rect 196354 7532 196364 7588
rect 196420 7532 209916 7588
rect 209972 7532 209982 7588
rect 591560 7560 593000 7784
rect 137778 7420 137788 7476
rect 137844 7420 145180 7476
rect 145236 7420 145246 7476
rect 200162 7420 200172 7476
rect 200228 7420 339388 7476
rect 339444 7420 339454 7476
rect 197474 7308 197484 7364
rect 197540 7308 496412 7364
rect 496468 7308 496478 7364
rect 195458 7196 195468 7252
rect 195524 7196 373660 7252
rect 373716 7196 373726 7252
rect 194114 7084 194124 7140
rect 194180 7084 366044 7140
rect 366100 7084 366110 7140
rect 203186 6860 203196 6916
rect 203252 6860 206780 6916
rect 206836 6860 206846 6916
rect 364 6748 28588 6804
rect 28644 6748 28654 6804
rect 141138 6748 141148 6804
rect 141204 6748 148540 6804
rect 148596 6748 148606 6804
rect 199378 6748 199388 6804
rect 199444 6748 199948 6804
rect 200004 6748 200014 6804
rect 206658 6748 206668 6804
rect 206724 6748 356188 6804
rect 356244 6748 356254 6804
rect 195682 6636 195692 6692
rect 195748 6636 503132 6692
rect 503188 6636 503198 6692
rect 192994 6524 193004 6580
rect 193060 6524 399308 6580
rect 399364 6524 399374 6580
rect 195906 6412 195916 6468
rect 195972 6412 270844 6468
rect 270900 6412 378812 6468
rect 378868 6412 378878 6468
rect 199154 6300 199164 6356
rect 199220 6300 259420 6356
rect 259476 6300 259486 6356
rect 297378 6300 297388 6356
rect 297444 6300 376348 6356
rect 376404 6300 376414 6356
rect 197362 6188 197372 6244
rect 197428 6188 232764 6244
rect 232820 6188 232830 6244
rect 312722 6188 312732 6244
rect 312788 6188 378028 6244
rect 378084 6188 378094 6244
rect 94098 6076 94108 6132
rect 94164 6076 144060 6132
rect 144116 6076 144126 6132
rect 197586 6076 197596 6132
rect 197652 6076 225148 6132
rect 225204 6076 225214 6132
rect 316530 6076 316540 6132
rect 316596 6076 378700 6132
rect 378756 6076 378766 6132
rect 122658 5964 122668 6020
rect 122724 5964 181468 6020
rect 181524 5964 181534 6020
rect 199714 5964 199724 6020
rect 199780 5964 230188 6020
rect 230244 5964 230254 6020
rect 343186 5964 343196 6020
rect 343252 5964 378252 6020
rect 378308 5964 378318 6020
rect 30258 5852 30268 5908
rect 30324 5852 204540 5908
rect 204596 5852 204606 5908
rect 205090 5852 205100 5908
rect 205156 5852 223356 5908
rect 223412 5852 223422 5908
rect 352594 5852 352604 5908
rect 352660 5852 556108 5908
rect 556164 5852 556174 5908
rect 189298 5740 189308 5796
rect 189364 5740 206668 5796
rect 206724 5740 206734 5796
rect 230290 5180 230300 5236
rect 230356 5180 314972 5236
rect 315028 5180 315038 5236
rect 224914 5068 224924 5124
rect 224980 5068 341628 5124
rect 341684 5068 341694 5124
rect 148642 4956 148652 5012
rect 148708 4956 150780 5012
rect 150836 4956 150846 5012
rect 160402 4956 160412 5012
rect 160468 4956 161980 5012
rect 162036 4956 162046 5012
rect 223346 4956 223356 5012
rect 223412 4956 230300 5012
rect 230356 4956 230366 5012
rect 157042 4844 157052 4900
rect 157108 4844 164220 4900
rect 164276 4844 164286 4900
rect 199826 4844 199836 4900
rect 199892 4844 274652 4900
rect 274708 4844 274718 4900
rect 277218 4844 277228 4900
rect 277284 4844 278460 4900
rect 278516 4844 378924 4900
rect 378980 4844 378990 4900
rect 145282 4732 145292 4788
rect 145348 4732 157500 4788
rect 157556 4732 157566 4788
rect 162082 4732 162092 4788
rect 162148 4732 170940 4788
rect 170996 4732 171006 4788
rect 194786 4732 194796 4788
rect 194852 4732 263228 4788
rect 263284 4732 263294 4788
rect 301298 4732 301308 4788
rect 301364 4732 377244 4788
rect 377300 4732 377310 4788
rect 134418 4620 134428 4676
rect 134484 4620 160860 4676
rect 160916 4620 160926 4676
rect 199938 4620 199948 4676
rect 200004 4620 205940 4676
rect 206770 4620 206780 4676
rect 206836 4620 251804 4676
rect 251860 4620 251870 4676
rect 305106 4620 305116 4676
rect 305172 4620 378028 4676
rect 378084 4620 378094 4676
rect 205884 4564 205940 4620
rect 98242 4508 98252 4564
rect 98308 4508 147420 4564
rect 147476 4508 147486 4564
rect 149492 4508 167580 4564
rect 167636 4508 167646 4564
rect 198594 4508 198604 4564
rect 198660 4508 205660 4564
rect 205716 4508 205726 4564
rect 205884 4508 240380 4564
rect 240436 4508 240446 4564
rect 324146 4508 324156 4564
rect 324212 4508 377468 4564
rect 377524 4508 377534 4564
rect 149492 4452 149548 4508
rect 113362 4396 113372 4452
rect 113428 4396 149548 4452
rect 163986 4396 163996 4452
rect 164052 4396 165340 4452
rect 165396 4396 165406 4452
rect 170258 4396 170268 4452
rect 170324 4396 187740 4452
rect 187796 4396 187806 4452
rect 195682 4396 195692 4452
rect 195748 4396 228956 4452
rect 229012 4396 229022 4452
rect 230178 4396 230188 4452
rect 230244 4396 255612 4452
rect 255668 4396 255678 4452
rect 331762 4396 331772 4452
rect 331828 4396 377580 4452
rect 377636 4396 377646 4452
rect 35298 4284 35308 4340
rect 35364 4284 198940 4340
rect 198996 4284 199006 4340
rect 199266 4284 199276 4340
rect 199332 4284 202300 4340
rect 202356 4284 202366 4340
rect 25218 4172 25228 4228
rect 25284 4172 198884 4228
rect 204978 4172 204988 4228
rect 205044 4172 528332 4228
rect 528388 4172 528398 4228
rect 198828 4116 198884 4172
rect 168914 4060 168924 4116
rect 168980 4060 171500 4116
rect 171556 4060 171566 4116
rect 180562 4060 180572 4116
rect 180628 4060 182140 4116
rect 182196 4060 182206 4116
rect 182354 4060 182364 4116
rect 182420 4060 185500 4116
rect 185556 4060 185566 4116
rect 190754 4060 190764 4116
rect 190820 4060 194460 4116
rect 194516 4060 194526 4116
rect 196578 4060 196588 4116
rect 196644 4060 197820 4116
rect 197876 4060 197886 4116
rect 198828 4060 201180 4116
rect 201236 4060 201246 4116
rect 195906 3948 195916 4004
rect 195972 3948 399084 4004
rect 399140 3948 399150 4004
rect 199042 3836 199052 3892
rect 199108 3836 221340 3892
rect 221396 3836 221406 3892
rect 198930 3724 198940 3780
rect 198996 3724 207900 3780
rect 207956 3724 207966 3780
rect 181458 3500 181468 3556
rect 181524 3500 184380 3556
rect 184436 3500 184446 3556
rect 226828 3388 330204 3444
rect 330260 3388 330270 3444
rect 226828 3332 226884 3388
rect 199042 3276 199052 3332
rect 199108 3276 226884 3332
rect 197474 3164 197484 3220
rect 197540 3164 204988 3220
rect 205044 3164 205054 3220
rect 205202 3164 205212 3220
rect 205268 3164 551068 3220
rect 551124 3164 551134 3220
rect 191314 3052 191324 3108
rect 191380 3052 297276 3108
rect 297332 3052 297342 3108
rect 314962 3052 314972 3108
rect 315028 3052 397180 3108
rect 397236 3052 397246 3108
rect 190642 2940 190652 2996
rect 190708 2940 286076 2996
rect 286132 2940 286142 2996
rect 293682 2940 293692 2996
rect 293748 2940 378140 2996
rect 378196 2940 378206 2996
rect 191426 2828 191436 2884
rect 191492 2828 277228 2884
rect 277284 2828 277294 2884
rect 330194 2828 330204 2884
rect 330260 2828 397516 2884
rect 397572 2828 397582 2884
rect 196466 2716 196476 2772
rect 196532 2716 282268 2772
rect 282324 2716 282334 2772
rect 347778 2716 347788 2772
rect 347844 2716 397740 2772
rect 397796 2716 397806 2772
rect 197922 2604 197932 2660
rect 197988 2604 205212 2660
rect 205268 2604 205278 2660
rect 205538 2604 205548 2660
rect 205604 2604 267036 2660
rect 267092 2604 267102 2660
rect 356178 2604 356188 2660
rect 356244 2604 399532 2660
rect 399588 2604 399598 2660
rect 180450 2492 180460 2548
rect 180516 2492 196588 2548
rect 198818 2492 198828 2548
rect 198884 2492 205324 2548
rect 205380 2492 205390 2548
rect 205660 2492 574588 2548
rect 574644 2492 574654 2548
rect 196532 2324 196588 2492
rect 205660 2324 205716 2492
rect 196532 2268 205716 2324
rect 198258 1596 198268 1652
rect 198324 1596 224924 1652
rect 224980 1596 224990 1652
rect 192882 1484 192892 1540
rect 192948 1484 398972 1540
rect 399028 1484 399038 1540
rect 193106 1372 193116 1428
rect 193172 1372 398860 1428
rect 398916 1372 398926 1428
rect 194674 1260 194684 1316
rect 194740 1260 400652 1316
rect 400708 1260 400718 1316
rect 194002 1148 194012 1204
rect 194068 1148 395612 1204
rect 395668 1148 395678 1204
rect 198034 1036 198044 1092
rect 198100 1036 293692 1092
rect 293748 1036 293758 1092
rect 341618 1036 341628 1092
rect 341684 1036 397068 1092
rect 397124 1036 397134 1092
rect 198034 924 198044 980
rect 198100 924 289884 980
rect 289940 924 289950 980
rect 197698 812 197708 868
rect 197764 812 244188 868
rect 244244 812 244254 868
rect 192658 700 192668 756
rect 192724 700 563612 756
rect 563668 700 563678 756
<< via3 >>
rect 9996 587916 10052 587972
rect 190652 587468 190708 587524
rect 197372 587244 197428 587300
rect 194012 587132 194068 587188
rect 7644 551180 7700 551236
rect 190876 539308 190932 539364
rect 197596 493948 197652 494004
rect 197484 316876 197540 316932
rect 9884 316764 9940 316820
rect 189196 316764 189252 316820
rect 189420 316652 189476 316708
rect 190764 316652 190820 316708
rect 198156 315084 198212 315140
rect 9772 313404 9828 313460
rect 199612 313292 199668 313348
rect 198044 310044 198100 310100
rect 376348 309932 376404 309988
rect 189084 308252 189140 308308
rect 188972 306572 189028 306628
rect 198156 305788 198212 305844
rect 189420 305228 189476 305284
rect 199052 305116 199108 305172
rect 195692 304892 195748 304948
rect 9660 303324 9716 303380
rect 397628 303324 397684 303380
rect 197708 300748 197764 300804
rect 397628 300748 397684 300804
rect 199388 169036 199444 169092
rect 198044 168588 198100 168644
rect 197260 168028 197316 168084
rect 378028 160860 378084 160916
rect 378028 159852 378084 159908
rect 198268 159628 198324 159684
rect 397628 159404 397684 159460
rect 197708 158844 197764 158900
rect 197932 158844 197988 158900
rect 198828 157948 198884 158004
rect 199612 157052 199668 157108
rect 211708 156828 211764 156884
rect 376348 156268 376404 156324
rect 551068 156268 551124 156324
rect 563612 156268 563668 156324
rect 197260 155932 197316 155988
rect 199836 155932 199892 155988
rect 378140 155820 378196 155876
rect 195804 155708 195860 155764
rect 528332 155148 528388 155204
rect 198156 154588 198212 154644
rect 9772 154476 9828 154532
rect 198044 154252 198100 154308
rect 205660 153916 205716 153972
rect 211708 153916 211764 153972
rect 197036 153692 197092 153748
rect 196252 153356 196308 153412
rect 205660 152796 205716 152852
rect 189420 152572 189476 152628
rect 199724 152460 199780 152516
rect 198156 152348 198212 152404
rect 198044 150892 198100 150948
rect 9660 150332 9716 150388
rect 197932 148652 197988 148708
rect 9884 146972 9940 147028
rect 190764 145516 190820 145572
rect 198828 145292 198884 145348
rect 198268 144620 198324 144676
rect 199164 144620 199220 144676
rect 197484 142044 197540 142100
rect 189196 140252 189252 140308
rect 199388 138684 199444 138740
rect 196252 138572 196308 138628
rect 195804 137004 195860 137060
rect 197036 133532 197092 133588
rect 199276 131068 199332 131124
rect 198268 129276 198324 129332
rect 199052 129276 199108 129332
rect 197484 126028 197540 126084
rect 189756 125916 189812 125972
rect 189756 124348 189812 124404
rect 199388 120988 199444 121044
rect 195692 118748 195748 118804
rect 189084 118524 189140 118580
rect 199052 117740 199108 117796
rect 195916 116284 195972 116340
rect 196252 116060 196308 116116
rect 195692 115948 195748 116004
rect 19516 114380 19572 114436
rect 19404 107660 19460 107716
rect 198268 104076 198324 104132
rect 16268 102284 16324 102340
rect 19964 100940 20020 100996
rect 19180 95564 19236 95620
rect 19740 94220 19796 94276
rect 16156 92876 16212 92932
rect 20076 91532 20132 91588
rect 19628 90188 19684 90244
rect 16044 87500 16100 87556
rect 22204 86156 22260 86212
rect 18396 84812 18452 84868
rect 20300 83468 20356 83524
rect 22316 82124 22372 82180
rect 20188 80780 20244 80836
rect 22092 73612 22148 73668
rect 21980 73500 22036 73556
rect 22092 73388 22148 73444
rect 20972 72492 21028 72548
rect 18284 70924 18340 70980
rect 18172 70700 18228 70756
rect 22092 70700 22148 70756
rect 23324 70700 23380 70756
rect 21980 70588 22036 70644
rect 22876 70588 22932 70644
rect 22204 70476 22260 70532
rect 23100 70476 23156 70532
rect 20076 69804 20132 69860
rect 190876 69132 190932 69188
rect 190652 68908 190708 68964
rect 197372 68796 197428 68852
rect 197596 68684 197652 68740
rect 36988 68572 37044 68628
rect 42028 68572 42084 68628
rect 48748 68572 48804 68628
rect 52108 68572 52164 68628
rect 53788 68572 53844 68628
rect 55468 68572 55524 68628
rect 19516 68460 19572 68516
rect 58828 68460 58884 68516
rect 60732 68460 60788 68516
rect 25564 68348 25620 68404
rect 28588 68348 28644 68404
rect 188972 66780 189028 66836
rect 194012 65436 194068 65492
rect 64540 53676 64596 53732
rect 64316 46396 64372 46452
rect 61964 35532 62020 35588
rect 61740 34748 61796 34804
rect 64092 33292 64148 33348
rect 63868 30380 63924 30436
rect 64204 28924 64260 28980
rect 63980 27468 64036 27524
rect 61964 27132 62020 27188
rect 61628 23884 61684 23940
rect 61852 21644 61908 21700
rect 63868 21420 63924 21476
rect 61628 21308 61684 21364
rect 60732 21084 60788 21140
rect 22652 20972 22708 21028
rect 60620 20860 60676 20916
rect 61628 20860 61684 20916
rect 61852 20188 61908 20244
rect 25564 20076 25620 20132
rect 64204 19852 64260 19908
rect 53788 19740 53844 19796
rect 20300 19628 20356 19684
rect 60620 19628 60676 19684
rect 23324 19516 23380 19572
rect 63980 19404 64036 19460
rect 9996 18396 10052 18452
rect 58828 18396 58884 18452
rect 19740 18284 19796 18340
rect 64316 18284 64372 18340
rect 23100 18172 23156 18228
rect 22764 18060 22820 18116
rect 64092 18060 64148 18116
rect 42028 17948 42084 18004
rect 7644 16716 7700 16772
rect 55468 16716 55524 16772
rect 19180 16604 19236 16660
rect 52108 16492 52164 16548
rect 19628 16380 19684 16436
rect 20188 16268 20244 16324
rect 36988 16156 37044 16212
rect 16268 14924 16324 14980
rect 16156 14812 16212 14868
rect 19964 14700 20020 14756
rect 64540 14700 64596 14756
rect 18396 14588 18452 14644
rect 22876 14476 22932 14532
rect 18284 13244 18340 13300
rect 19404 13132 19460 13188
rect 20972 13020 21028 13076
rect 18172 12908 18228 12964
rect 48748 12796 48804 12852
rect 196252 10332 196308 10388
rect 16044 9996 16100 10052
rect 199276 9996 199332 10052
rect 199500 9548 199556 9604
rect 197484 7308 197540 7364
rect 28588 6748 28644 6804
rect 195692 6636 195748 6692
rect 199164 6300 199220 6356
rect 376348 6300 376404 6356
rect 199724 5964 199780 6020
rect 199836 4844 199892 4900
rect 378028 4620 378084 4676
rect 198940 4284 198996 4340
rect 528332 4172 528388 4228
rect 195916 3948 195972 4004
rect 198940 3724 198996 3780
rect 199052 3276 199108 3332
rect 551068 3164 551124 3220
rect 378140 2940 378196 2996
rect 198044 924 198100 980
rect 563612 700 563668 756
<< metal4 >>
rect -1916 598172 -1296 598268
rect -1916 598116 -1820 598172
rect -1764 598116 -1696 598172
rect -1640 598116 -1572 598172
rect -1516 598116 -1448 598172
rect -1392 598116 -1296 598172
rect -1916 598048 -1296 598116
rect -1916 597992 -1820 598048
rect -1764 597992 -1696 598048
rect -1640 597992 -1572 598048
rect -1516 597992 -1448 598048
rect -1392 597992 -1296 598048
rect -1916 597924 -1296 597992
rect -1916 597868 -1820 597924
rect -1764 597868 -1696 597924
rect -1640 597868 -1572 597924
rect -1516 597868 -1448 597924
rect -1392 597868 -1296 597924
rect -1916 597800 -1296 597868
rect -1916 597744 -1820 597800
rect -1764 597744 -1696 597800
rect -1640 597744 -1572 597800
rect -1516 597744 -1448 597800
rect -1392 597744 -1296 597800
rect -1916 586350 -1296 597744
rect -1916 586294 -1820 586350
rect -1764 586294 -1696 586350
rect -1640 586294 -1572 586350
rect -1516 586294 -1448 586350
rect -1392 586294 -1296 586350
rect -1916 586226 -1296 586294
rect -1916 586170 -1820 586226
rect -1764 586170 -1696 586226
rect -1640 586170 -1572 586226
rect -1516 586170 -1448 586226
rect -1392 586170 -1296 586226
rect -1916 586102 -1296 586170
rect -1916 586046 -1820 586102
rect -1764 586046 -1696 586102
rect -1640 586046 -1572 586102
rect -1516 586046 -1448 586102
rect -1392 586046 -1296 586102
rect -1916 585978 -1296 586046
rect -1916 585922 -1820 585978
rect -1764 585922 -1696 585978
rect -1640 585922 -1572 585978
rect -1516 585922 -1448 585978
rect -1392 585922 -1296 585978
rect -1916 568350 -1296 585922
rect -1916 568294 -1820 568350
rect -1764 568294 -1696 568350
rect -1640 568294 -1572 568350
rect -1516 568294 -1448 568350
rect -1392 568294 -1296 568350
rect -1916 568226 -1296 568294
rect -1916 568170 -1820 568226
rect -1764 568170 -1696 568226
rect -1640 568170 -1572 568226
rect -1516 568170 -1448 568226
rect -1392 568170 -1296 568226
rect -1916 568102 -1296 568170
rect -1916 568046 -1820 568102
rect -1764 568046 -1696 568102
rect -1640 568046 -1572 568102
rect -1516 568046 -1448 568102
rect -1392 568046 -1296 568102
rect -1916 567978 -1296 568046
rect -1916 567922 -1820 567978
rect -1764 567922 -1696 567978
rect -1640 567922 -1572 567978
rect -1516 567922 -1448 567978
rect -1392 567922 -1296 567978
rect -1916 550350 -1296 567922
rect -1916 550294 -1820 550350
rect -1764 550294 -1696 550350
rect -1640 550294 -1572 550350
rect -1516 550294 -1448 550350
rect -1392 550294 -1296 550350
rect -1916 550226 -1296 550294
rect -1916 550170 -1820 550226
rect -1764 550170 -1696 550226
rect -1640 550170 -1572 550226
rect -1516 550170 -1448 550226
rect -1392 550170 -1296 550226
rect -1916 550102 -1296 550170
rect -1916 550046 -1820 550102
rect -1764 550046 -1696 550102
rect -1640 550046 -1572 550102
rect -1516 550046 -1448 550102
rect -1392 550046 -1296 550102
rect -1916 549978 -1296 550046
rect -1916 549922 -1820 549978
rect -1764 549922 -1696 549978
rect -1640 549922 -1572 549978
rect -1516 549922 -1448 549978
rect -1392 549922 -1296 549978
rect -1916 532350 -1296 549922
rect -1916 532294 -1820 532350
rect -1764 532294 -1696 532350
rect -1640 532294 -1572 532350
rect -1516 532294 -1448 532350
rect -1392 532294 -1296 532350
rect -1916 532226 -1296 532294
rect -1916 532170 -1820 532226
rect -1764 532170 -1696 532226
rect -1640 532170 -1572 532226
rect -1516 532170 -1448 532226
rect -1392 532170 -1296 532226
rect -1916 532102 -1296 532170
rect -1916 532046 -1820 532102
rect -1764 532046 -1696 532102
rect -1640 532046 -1572 532102
rect -1516 532046 -1448 532102
rect -1392 532046 -1296 532102
rect -1916 531978 -1296 532046
rect -1916 531922 -1820 531978
rect -1764 531922 -1696 531978
rect -1640 531922 -1572 531978
rect -1516 531922 -1448 531978
rect -1392 531922 -1296 531978
rect -1916 514350 -1296 531922
rect -1916 514294 -1820 514350
rect -1764 514294 -1696 514350
rect -1640 514294 -1572 514350
rect -1516 514294 -1448 514350
rect -1392 514294 -1296 514350
rect -1916 514226 -1296 514294
rect -1916 514170 -1820 514226
rect -1764 514170 -1696 514226
rect -1640 514170 -1572 514226
rect -1516 514170 -1448 514226
rect -1392 514170 -1296 514226
rect -1916 514102 -1296 514170
rect -1916 514046 -1820 514102
rect -1764 514046 -1696 514102
rect -1640 514046 -1572 514102
rect -1516 514046 -1448 514102
rect -1392 514046 -1296 514102
rect -1916 513978 -1296 514046
rect -1916 513922 -1820 513978
rect -1764 513922 -1696 513978
rect -1640 513922 -1572 513978
rect -1516 513922 -1448 513978
rect -1392 513922 -1296 513978
rect -1916 496350 -1296 513922
rect -1916 496294 -1820 496350
rect -1764 496294 -1696 496350
rect -1640 496294 -1572 496350
rect -1516 496294 -1448 496350
rect -1392 496294 -1296 496350
rect -1916 496226 -1296 496294
rect -1916 496170 -1820 496226
rect -1764 496170 -1696 496226
rect -1640 496170 -1572 496226
rect -1516 496170 -1448 496226
rect -1392 496170 -1296 496226
rect -1916 496102 -1296 496170
rect -1916 496046 -1820 496102
rect -1764 496046 -1696 496102
rect -1640 496046 -1572 496102
rect -1516 496046 -1448 496102
rect -1392 496046 -1296 496102
rect -1916 495978 -1296 496046
rect -1916 495922 -1820 495978
rect -1764 495922 -1696 495978
rect -1640 495922 -1572 495978
rect -1516 495922 -1448 495978
rect -1392 495922 -1296 495978
rect -1916 478350 -1296 495922
rect -1916 478294 -1820 478350
rect -1764 478294 -1696 478350
rect -1640 478294 -1572 478350
rect -1516 478294 -1448 478350
rect -1392 478294 -1296 478350
rect -1916 478226 -1296 478294
rect -1916 478170 -1820 478226
rect -1764 478170 -1696 478226
rect -1640 478170 -1572 478226
rect -1516 478170 -1448 478226
rect -1392 478170 -1296 478226
rect -1916 478102 -1296 478170
rect -1916 478046 -1820 478102
rect -1764 478046 -1696 478102
rect -1640 478046 -1572 478102
rect -1516 478046 -1448 478102
rect -1392 478046 -1296 478102
rect -1916 477978 -1296 478046
rect -1916 477922 -1820 477978
rect -1764 477922 -1696 477978
rect -1640 477922 -1572 477978
rect -1516 477922 -1448 477978
rect -1392 477922 -1296 477978
rect -1916 460350 -1296 477922
rect -1916 460294 -1820 460350
rect -1764 460294 -1696 460350
rect -1640 460294 -1572 460350
rect -1516 460294 -1448 460350
rect -1392 460294 -1296 460350
rect -1916 460226 -1296 460294
rect -1916 460170 -1820 460226
rect -1764 460170 -1696 460226
rect -1640 460170 -1572 460226
rect -1516 460170 -1448 460226
rect -1392 460170 -1296 460226
rect -1916 460102 -1296 460170
rect -1916 460046 -1820 460102
rect -1764 460046 -1696 460102
rect -1640 460046 -1572 460102
rect -1516 460046 -1448 460102
rect -1392 460046 -1296 460102
rect -1916 459978 -1296 460046
rect -1916 459922 -1820 459978
rect -1764 459922 -1696 459978
rect -1640 459922 -1572 459978
rect -1516 459922 -1448 459978
rect -1392 459922 -1296 459978
rect -1916 442350 -1296 459922
rect -1916 442294 -1820 442350
rect -1764 442294 -1696 442350
rect -1640 442294 -1572 442350
rect -1516 442294 -1448 442350
rect -1392 442294 -1296 442350
rect -1916 442226 -1296 442294
rect -1916 442170 -1820 442226
rect -1764 442170 -1696 442226
rect -1640 442170 -1572 442226
rect -1516 442170 -1448 442226
rect -1392 442170 -1296 442226
rect -1916 442102 -1296 442170
rect -1916 442046 -1820 442102
rect -1764 442046 -1696 442102
rect -1640 442046 -1572 442102
rect -1516 442046 -1448 442102
rect -1392 442046 -1296 442102
rect -1916 441978 -1296 442046
rect -1916 441922 -1820 441978
rect -1764 441922 -1696 441978
rect -1640 441922 -1572 441978
rect -1516 441922 -1448 441978
rect -1392 441922 -1296 441978
rect -1916 424350 -1296 441922
rect -1916 424294 -1820 424350
rect -1764 424294 -1696 424350
rect -1640 424294 -1572 424350
rect -1516 424294 -1448 424350
rect -1392 424294 -1296 424350
rect -1916 424226 -1296 424294
rect -1916 424170 -1820 424226
rect -1764 424170 -1696 424226
rect -1640 424170 -1572 424226
rect -1516 424170 -1448 424226
rect -1392 424170 -1296 424226
rect -1916 424102 -1296 424170
rect -1916 424046 -1820 424102
rect -1764 424046 -1696 424102
rect -1640 424046 -1572 424102
rect -1516 424046 -1448 424102
rect -1392 424046 -1296 424102
rect -1916 423978 -1296 424046
rect -1916 423922 -1820 423978
rect -1764 423922 -1696 423978
rect -1640 423922 -1572 423978
rect -1516 423922 -1448 423978
rect -1392 423922 -1296 423978
rect -1916 406350 -1296 423922
rect -1916 406294 -1820 406350
rect -1764 406294 -1696 406350
rect -1640 406294 -1572 406350
rect -1516 406294 -1448 406350
rect -1392 406294 -1296 406350
rect -1916 406226 -1296 406294
rect -1916 406170 -1820 406226
rect -1764 406170 -1696 406226
rect -1640 406170 -1572 406226
rect -1516 406170 -1448 406226
rect -1392 406170 -1296 406226
rect -1916 406102 -1296 406170
rect -1916 406046 -1820 406102
rect -1764 406046 -1696 406102
rect -1640 406046 -1572 406102
rect -1516 406046 -1448 406102
rect -1392 406046 -1296 406102
rect -1916 405978 -1296 406046
rect -1916 405922 -1820 405978
rect -1764 405922 -1696 405978
rect -1640 405922 -1572 405978
rect -1516 405922 -1448 405978
rect -1392 405922 -1296 405978
rect -1916 388350 -1296 405922
rect -1916 388294 -1820 388350
rect -1764 388294 -1696 388350
rect -1640 388294 -1572 388350
rect -1516 388294 -1448 388350
rect -1392 388294 -1296 388350
rect -1916 388226 -1296 388294
rect -1916 388170 -1820 388226
rect -1764 388170 -1696 388226
rect -1640 388170 -1572 388226
rect -1516 388170 -1448 388226
rect -1392 388170 -1296 388226
rect -1916 388102 -1296 388170
rect -1916 388046 -1820 388102
rect -1764 388046 -1696 388102
rect -1640 388046 -1572 388102
rect -1516 388046 -1448 388102
rect -1392 388046 -1296 388102
rect -1916 387978 -1296 388046
rect -1916 387922 -1820 387978
rect -1764 387922 -1696 387978
rect -1640 387922 -1572 387978
rect -1516 387922 -1448 387978
rect -1392 387922 -1296 387978
rect -1916 370350 -1296 387922
rect -1916 370294 -1820 370350
rect -1764 370294 -1696 370350
rect -1640 370294 -1572 370350
rect -1516 370294 -1448 370350
rect -1392 370294 -1296 370350
rect -1916 370226 -1296 370294
rect -1916 370170 -1820 370226
rect -1764 370170 -1696 370226
rect -1640 370170 -1572 370226
rect -1516 370170 -1448 370226
rect -1392 370170 -1296 370226
rect -1916 370102 -1296 370170
rect -1916 370046 -1820 370102
rect -1764 370046 -1696 370102
rect -1640 370046 -1572 370102
rect -1516 370046 -1448 370102
rect -1392 370046 -1296 370102
rect -1916 369978 -1296 370046
rect -1916 369922 -1820 369978
rect -1764 369922 -1696 369978
rect -1640 369922 -1572 369978
rect -1516 369922 -1448 369978
rect -1392 369922 -1296 369978
rect -1916 352350 -1296 369922
rect -1916 352294 -1820 352350
rect -1764 352294 -1696 352350
rect -1640 352294 -1572 352350
rect -1516 352294 -1448 352350
rect -1392 352294 -1296 352350
rect -1916 352226 -1296 352294
rect -1916 352170 -1820 352226
rect -1764 352170 -1696 352226
rect -1640 352170 -1572 352226
rect -1516 352170 -1448 352226
rect -1392 352170 -1296 352226
rect -1916 352102 -1296 352170
rect -1916 352046 -1820 352102
rect -1764 352046 -1696 352102
rect -1640 352046 -1572 352102
rect -1516 352046 -1448 352102
rect -1392 352046 -1296 352102
rect -1916 351978 -1296 352046
rect -1916 351922 -1820 351978
rect -1764 351922 -1696 351978
rect -1640 351922 -1572 351978
rect -1516 351922 -1448 351978
rect -1392 351922 -1296 351978
rect -1916 334350 -1296 351922
rect -1916 334294 -1820 334350
rect -1764 334294 -1696 334350
rect -1640 334294 -1572 334350
rect -1516 334294 -1448 334350
rect -1392 334294 -1296 334350
rect -1916 334226 -1296 334294
rect -1916 334170 -1820 334226
rect -1764 334170 -1696 334226
rect -1640 334170 -1572 334226
rect -1516 334170 -1448 334226
rect -1392 334170 -1296 334226
rect -1916 334102 -1296 334170
rect -1916 334046 -1820 334102
rect -1764 334046 -1696 334102
rect -1640 334046 -1572 334102
rect -1516 334046 -1448 334102
rect -1392 334046 -1296 334102
rect -1916 333978 -1296 334046
rect -1916 333922 -1820 333978
rect -1764 333922 -1696 333978
rect -1640 333922 -1572 333978
rect -1516 333922 -1448 333978
rect -1392 333922 -1296 333978
rect -1916 316350 -1296 333922
rect -1916 316294 -1820 316350
rect -1764 316294 -1696 316350
rect -1640 316294 -1572 316350
rect -1516 316294 -1448 316350
rect -1392 316294 -1296 316350
rect -1916 316226 -1296 316294
rect -1916 316170 -1820 316226
rect -1764 316170 -1696 316226
rect -1640 316170 -1572 316226
rect -1516 316170 -1448 316226
rect -1392 316170 -1296 316226
rect -1916 316102 -1296 316170
rect -1916 316046 -1820 316102
rect -1764 316046 -1696 316102
rect -1640 316046 -1572 316102
rect -1516 316046 -1448 316102
rect -1392 316046 -1296 316102
rect -1916 315978 -1296 316046
rect -1916 315922 -1820 315978
rect -1764 315922 -1696 315978
rect -1640 315922 -1572 315978
rect -1516 315922 -1448 315978
rect -1392 315922 -1296 315978
rect -1916 298350 -1296 315922
rect -1916 298294 -1820 298350
rect -1764 298294 -1696 298350
rect -1640 298294 -1572 298350
rect -1516 298294 -1448 298350
rect -1392 298294 -1296 298350
rect -1916 298226 -1296 298294
rect -1916 298170 -1820 298226
rect -1764 298170 -1696 298226
rect -1640 298170 -1572 298226
rect -1516 298170 -1448 298226
rect -1392 298170 -1296 298226
rect -1916 298102 -1296 298170
rect -1916 298046 -1820 298102
rect -1764 298046 -1696 298102
rect -1640 298046 -1572 298102
rect -1516 298046 -1448 298102
rect -1392 298046 -1296 298102
rect -1916 297978 -1296 298046
rect -1916 297922 -1820 297978
rect -1764 297922 -1696 297978
rect -1640 297922 -1572 297978
rect -1516 297922 -1448 297978
rect -1392 297922 -1296 297978
rect -1916 280350 -1296 297922
rect -1916 280294 -1820 280350
rect -1764 280294 -1696 280350
rect -1640 280294 -1572 280350
rect -1516 280294 -1448 280350
rect -1392 280294 -1296 280350
rect -1916 280226 -1296 280294
rect -1916 280170 -1820 280226
rect -1764 280170 -1696 280226
rect -1640 280170 -1572 280226
rect -1516 280170 -1448 280226
rect -1392 280170 -1296 280226
rect -1916 280102 -1296 280170
rect -1916 280046 -1820 280102
rect -1764 280046 -1696 280102
rect -1640 280046 -1572 280102
rect -1516 280046 -1448 280102
rect -1392 280046 -1296 280102
rect -1916 279978 -1296 280046
rect -1916 279922 -1820 279978
rect -1764 279922 -1696 279978
rect -1640 279922 -1572 279978
rect -1516 279922 -1448 279978
rect -1392 279922 -1296 279978
rect -1916 262350 -1296 279922
rect -1916 262294 -1820 262350
rect -1764 262294 -1696 262350
rect -1640 262294 -1572 262350
rect -1516 262294 -1448 262350
rect -1392 262294 -1296 262350
rect -1916 262226 -1296 262294
rect -1916 262170 -1820 262226
rect -1764 262170 -1696 262226
rect -1640 262170 -1572 262226
rect -1516 262170 -1448 262226
rect -1392 262170 -1296 262226
rect -1916 262102 -1296 262170
rect -1916 262046 -1820 262102
rect -1764 262046 -1696 262102
rect -1640 262046 -1572 262102
rect -1516 262046 -1448 262102
rect -1392 262046 -1296 262102
rect -1916 261978 -1296 262046
rect -1916 261922 -1820 261978
rect -1764 261922 -1696 261978
rect -1640 261922 -1572 261978
rect -1516 261922 -1448 261978
rect -1392 261922 -1296 261978
rect -1916 244350 -1296 261922
rect -1916 244294 -1820 244350
rect -1764 244294 -1696 244350
rect -1640 244294 -1572 244350
rect -1516 244294 -1448 244350
rect -1392 244294 -1296 244350
rect -1916 244226 -1296 244294
rect -1916 244170 -1820 244226
rect -1764 244170 -1696 244226
rect -1640 244170 -1572 244226
rect -1516 244170 -1448 244226
rect -1392 244170 -1296 244226
rect -1916 244102 -1296 244170
rect -1916 244046 -1820 244102
rect -1764 244046 -1696 244102
rect -1640 244046 -1572 244102
rect -1516 244046 -1448 244102
rect -1392 244046 -1296 244102
rect -1916 243978 -1296 244046
rect -1916 243922 -1820 243978
rect -1764 243922 -1696 243978
rect -1640 243922 -1572 243978
rect -1516 243922 -1448 243978
rect -1392 243922 -1296 243978
rect -1916 226350 -1296 243922
rect -1916 226294 -1820 226350
rect -1764 226294 -1696 226350
rect -1640 226294 -1572 226350
rect -1516 226294 -1448 226350
rect -1392 226294 -1296 226350
rect -1916 226226 -1296 226294
rect -1916 226170 -1820 226226
rect -1764 226170 -1696 226226
rect -1640 226170 -1572 226226
rect -1516 226170 -1448 226226
rect -1392 226170 -1296 226226
rect -1916 226102 -1296 226170
rect -1916 226046 -1820 226102
rect -1764 226046 -1696 226102
rect -1640 226046 -1572 226102
rect -1516 226046 -1448 226102
rect -1392 226046 -1296 226102
rect -1916 225978 -1296 226046
rect -1916 225922 -1820 225978
rect -1764 225922 -1696 225978
rect -1640 225922 -1572 225978
rect -1516 225922 -1448 225978
rect -1392 225922 -1296 225978
rect -1916 208350 -1296 225922
rect -1916 208294 -1820 208350
rect -1764 208294 -1696 208350
rect -1640 208294 -1572 208350
rect -1516 208294 -1448 208350
rect -1392 208294 -1296 208350
rect -1916 208226 -1296 208294
rect -1916 208170 -1820 208226
rect -1764 208170 -1696 208226
rect -1640 208170 -1572 208226
rect -1516 208170 -1448 208226
rect -1392 208170 -1296 208226
rect -1916 208102 -1296 208170
rect -1916 208046 -1820 208102
rect -1764 208046 -1696 208102
rect -1640 208046 -1572 208102
rect -1516 208046 -1448 208102
rect -1392 208046 -1296 208102
rect -1916 207978 -1296 208046
rect -1916 207922 -1820 207978
rect -1764 207922 -1696 207978
rect -1640 207922 -1572 207978
rect -1516 207922 -1448 207978
rect -1392 207922 -1296 207978
rect -1916 190350 -1296 207922
rect -1916 190294 -1820 190350
rect -1764 190294 -1696 190350
rect -1640 190294 -1572 190350
rect -1516 190294 -1448 190350
rect -1392 190294 -1296 190350
rect -1916 190226 -1296 190294
rect -1916 190170 -1820 190226
rect -1764 190170 -1696 190226
rect -1640 190170 -1572 190226
rect -1516 190170 -1448 190226
rect -1392 190170 -1296 190226
rect -1916 190102 -1296 190170
rect -1916 190046 -1820 190102
rect -1764 190046 -1696 190102
rect -1640 190046 -1572 190102
rect -1516 190046 -1448 190102
rect -1392 190046 -1296 190102
rect -1916 189978 -1296 190046
rect -1916 189922 -1820 189978
rect -1764 189922 -1696 189978
rect -1640 189922 -1572 189978
rect -1516 189922 -1448 189978
rect -1392 189922 -1296 189978
rect -1916 172350 -1296 189922
rect -1916 172294 -1820 172350
rect -1764 172294 -1696 172350
rect -1640 172294 -1572 172350
rect -1516 172294 -1448 172350
rect -1392 172294 -1296 172350
rect -1916 172226 -1296 172294
rect -1916 172170 -1820 172226
rect -1764 172170 -1696 172226
rect -1640 172170 -1572 172226
rect -1516 172170 -1448 172226
rect -1392 172170 -1296 172226
rect -1916 172102 -1296 172170
rect -1916 172046 -1820 172102
rect -1764 172046 -1696 172102
rect -1640 172046 -1572 172102
rect -1516 172046 -1448 172102
rect -1392 172046 -1296 172102
rect -1916 171978 -1296 172046
rect -1916 171922 -1820 171978
rect -1764 171922 -1696 171978
rect -1640 171922 -1572 171978
rect -1516 171922 -1448 171978
rect -1392 171922 -1296 171978
rect -1916 154350 -1296 171922
rect -1916 154294 -1820 154350
rect -1764 154294 -1696 154350
rect -1640 154294 -1572 154350
rect -1516 154294 -1448 154350
rect -1392 154294 -1296 154350
rect -1916 154226 -1296 154294
rect -1916 154170 -1820 154226
rect -1764 154170 -1696 154226
rect -1640 154170 -1572 154226
rect -1516 154170 -1448 154226
rect -1392 154170 -1296 154226
rect -1916 154102 -1296 154170
rect -1916 154046 -1820 154102
rect -1764 154046 -1696 154102
rect -1640 154046 -1572 154102
rect -1516 154046 -1448 154102
rect -1392 154046 -1296 154102
rect -1916 153978 -1296 154046
rect -1916 153922 -1820 153978
rect -1764 153922 -1696 153978
rect -1640 153922 -1572 153978
rect -1516 153922 -1448 153978
rect -1392 153922 -1296 153978
rect -1916 136350 -1296 153922
rect -1916 136294 -1820 136350
rect -1764 136294 -1696 136350
rect -1640 136294 -1572 136350
rect -1516 136294 -1448 136350
rect -1392 136294 -1296 136350
rect -1916 136226 -1296 136294
rect -1916 136170 -1820 136226
rect -1764 136170 -1696 136226
rect -1640 136170 -1572 136226
rect -1516 136170 -1448 136226
rect -1392 136170 -1296 136226
rect -1916 136102 -1296 136170
rect -1916 136046 -1820 136102
rect -1764 136046 -1696 136102
rect -1640 136046 -1572 136102
rect -1516 136046 -1448 136102
rect -1392 136046 -1296 136102
rect -1916 135978 -1296 136046
rect -1916 135922 -1820 135978
rect -1764 135922 -1696 135978
rect -1640 135922 -1572 135978
rect -1516 135922 -1448 135978
rect -1392 135922 -1296 135978
rect -1916 118350 -1296 135922
rect -1916 118294 -1820 118350
rect -1764 118294 -1696 118350
rect -1640 118294 -1572 118350
rect -1516 118294 -1448 118350
rect -1392 118294 -1296 118350
rect -1916 118226 -1296 118294
rect -1916 118170 -1820 118226
rect -1764 118170 -1696 118226
rect -1640 118170 -1572 118226
rect -1516 118170 -1448 118226
rect -1392 118170 -1296 118226
rect -1916 118102 -1296 118170
rect -1916 118046 -1820 118102
rect -1764 118046 -1696 118102
rect -1640 118046 -1572 118102
rect -1516 118046 -1448 118102
rect -1392 118046 -1296 118102
rect -1916 117978 -1296 118046
rect -1916 117922 -1820 117978
rect -1764 117922 -1696 117978
rect -1640 117922 -1572 117978
rect -1516 117922 -1448 117978
rect -1392 117922 -1296 117978
rect -1916 100350 -1296 117922
rect -1916 100294 -1820 100350
rect -1764 100294 -1696 100350
rect -1640 100294 -1572 100350
rect -1516 100294 -1448 100350
rect -1392 100294 -1296 100350
rect -1916 100226 -1296 100294
rect -1916 100170 -1820 100226
rect -1764 100170 -1696 100226
rect -1640 100170 -1572 100226
rect -1516 100170 -1448 100226
rect -1392 100170 -1296 100226
rect -1916 100102 -1296 100170
rect -1916 100046 -1820 100102
rect -1764 100046 -1696 100102
rect -1640 100046 -1572 100102
rect -1516 100046 -1448 100102
rect -1392 100046 -1296 100102
rect -1916 99978 -1296 100046
rect -1916 99922 -1820 99978
rect -1764 99922 -1696 99978
rect -1640 99922 -1572 99978
rect -1516 99922 -1448 99978
rect -1392 99922 -1296 99978
rect -1916 82350 -1296 99922
rect -1916 82294 -1820 82350
rect -1764 82294 -1696 82350
rect -1640 82294 -1572 82350
rect -1516 82294 -1448 82350
rect -1392 82294 -1296 82350
rect -1916 82226 -1296 82294
rect -1916 82170 -1820 82226
rect -1764 82170 -1696 82226
rect -1640 82170 -1572 82226
rect -1516 82170 -1448 82226
rect -1392 82170 -1296 82226
rect -1916 82102 -1296 82170
rect -1916 82046 -1820 82102
rect -1764 82046 -1696 82102
rect -1640 82046 -1572 82102
rect -1516 82046 -1448 82102
rect -1392 82046 -1296 82102
rect -1916 81978 -1296 82046
rect -1916 81922 -1820 81978
rect -1764 81922 -1696 81978
rect -1640 81922 -1572 81978
rect -1516 81922 -1448 81978
rect -1392 81922 -1296 81978
rect -1916 64350 -1296 81922
rect -1916 64294 -1820 64350
rect -1764 64294 -1696 64350
rect -1640 64294 -1572 64350
rect -1516 64294 -1448 64350
rect -1392 64294 -1296 64350
rect -1916 64226 -1296 64294
rect -1916 64170 -1820 64226
rect -1764 64170 -1696 64226
rect -1640 64170 -1572 64226
rect -1516 64170 -1448 64226
rect -1392 64170 -1296 64226
rect -1916 64102 -1296 64170
rect -1916 64046 -1820 64102
rect -1764 64046 -1696 64102
rect -1640 64046 -1572 64102
rect -1516 64046 -1448 64102
rect -1392 64046 -1296 64102
rect -1916 63978 -1296 64046
rect -1916 63922 -1820 63978
rect -1764 63922 -1696 63978
rect -1640 63922 -1572 63978
rect -1516 63922 -1448 63978
rect -1392 63922 -1296 63978
rect -1916 46350 -1296 63922
rect -1916 46294 -1820 46350
rect -1764 46294 -1696 46350
rect -1640 46294 -1572 46350
rect -1516 46294 -1448 46350
rect -1392 46294 -1296 46350
rect -1916 46226 -1296 46294
rect -1916 46170 -1820 46226
rect -1764 46170 -1696 46226
rect -1640 46170 -1572 46226
rect -1516 46170 -1448 46226
rect -1392 46170 -1296 46226
rect -1916 46102 -1296 46170
rect -1916 46046 -1820 46102
rect -1764 46046 -1696 46102
rect -1640 46046 -1572 46102
rect -1516 46046 -1448 46102
rect -1392 46046 -1296 46102
rect -1916 45978 -1296 46046
rect -1916 45922 -1820 45978
rect -1764 45922 -1696 45978
rect -1640 45922 -1572 45978
rect -1516 45922 -1448 45978
rect -1392 45922 -1296 45978
rect -1916 28350 -1296 45922
rect -1916 28294 -1820 28350
rect -1764 28294 -1696 28350
rect -1640 28294 -1572 28350
rect -1516 28294 -1448 28350
rect -1392 28294 -1296 28350
rect -1916 28226 -1296 28294
rect -1916 28170 -1820 28226
rect -1764 28170 -1696 28226
rect -1640 28170 -1572 28226
rect -1516 28170 -1448 28226
rect -1392 28170 -1296 28226
rect -1916 28102 -1296 28170
rect -1916 28046 -1820 28102
rect -1764 28046 -1696 28102
rect -1640 28046 -1572 28102
rect -1516 28046 -1448 28102
rect -1392 28046 -1296 28102
rect -1916 27978 -1296 28046
rect -1916 27922 -1820 27978
rect -1764 27922 -1696 27978
rect -1640 27922 -1572 27978
rect -1516 27922 -1448 27978
rect -1392 27922 -1296 27978
rect -1916 10350 -1296 27922
rect -1916 10294 -1820 10350
rect -1764 10294 -1696 10350
rect -1640 10294 -1572 10350
rect -1516 10294 -1448 10350
rect -1392 10294 -1296 10350
rect -1916 10226 -1296 10294
rect -1916 10170 -1820 10226
rect -1764 10170 -1696 10226
rect -1640 10170 -1572 10226
rect -1516 10170 -1448 10226
rect -1392 10170 -1296 10226
rect -1916 10102 -1296 10170
rect -1916 10046 -1820 10102
rect -1764 10046 -1696 10102
rect -1640 10046 -1572 10102
rect -1516 10046 -1448 10102
rect -1392 10046 -1296 10102
rect -1916 9978 -1296 10046
rect -1916 9922 -1820 9978
rect -1764 9922 -1696 9978
rect -1640 9922 -1572 9978
rect -1516 9922 -1448 9978
rect -1392 9922 -1296 9978
rect -1916 -1120 -1296 9922
rect -956 597212 -336 597308
rect -956 597156 -860 597212
rect -804 597156 -736 597212
rect -680 597156 -612 597212
rect -556 597156 -488 597212
rect -432 597156 -336 597212
rect -956 597088 -336 597156
rect -956 597032 -860 597088
rect -804 597032 -736 597088
rect -680 597032 -612 597088
rect -556 597032 -488 597088
rect -432 597032 -336 597088
rect -956 596964 -336 597032
rect -956 596908 -860 596964
rect -804 596908 -736 596964
rect -680 596908 -612 596964
rect -556 596908 -488 596964
rect -432 596908 -336 596964
rect -956 596840 -336 596908
rect -956 596784 -860 596840
rect -804 596784 -736 596840
rect -680 596784 -612 596840
rect -556 596784 -488 596840
rect -432 596784 -336 596840
rect -956 580350 -336 596784
rect -956 580294 -860 580350
rect -804 580294 -736 580350
rect -680 580294 -612 580350
rect -556 580294 -488 580350
rect -432 580294 -336 580350
rect -956 580226 -336 580294
rect -956 580170 -860 580226
rect -804 580170 -736 580226
rect -680 580170 -612 580226
rect -556 580170 -488 580226
rect -432 580170 -336 580226
rect -956 580102 -336 580170
rect -956 580046 -860 580102
rect -804 580046 -736 580102
rect -680 580046 -612 580102
rect -556 580046 -488 580102
rect -432 580046 -336 580102
rect -956 579978 -336 580046
rect -956 579922 -860 579978
rect -804 579922 -736 579978
rect -680 579922 -612 579978
rect -556 579922 -488 579978
rect -432 579922 -336 579978
rect -956 562350 -336 579922
rect -956 562294 -860 562350
rect -804 562294 -736 562350
rect -680 562294 -612 562350
rect -556 562294 -488 562350
rect -432 562294 -336 562350
rect -956 562226 -336 562294
rect -956 562170 -860 562226
rect -804 562170 -736 562226
rect -680 562170 -612 562226
rect -556 562170 -488 562226
rect -432 562170 -336 562226
rect -956 562102 -336 562170
rect -956 562046 -860 562102
rect -804 562046 -736 562102
rect -680 562046 -612 562102
rect -556 562046 -488 562102
rect -432 562046 -336 562102
rect -956 561978 -336 562046
rect -956 561922 -860 561978
rect -804 561922 -736 561978
rect -680 561922 -612 561978
rect -556 561922 -488 561978
rect -432 561922 -336 561978
rect -956 544350 -336 561922
rect -956 544294 -860 544350
rect -804 544294 -736 544350
rect -680 544294 -612 544350
rect -556 544294 -488 544350
rect -432 544294 -336 544350
rect -956 544226 -336 544294
rect -956 544170 -860 544226
rect -804 544170 -736 544226
rect -680 544170 -612 544226
rect -556 544170 -488 544226
rect -432 544170 -336 544226
rect -956 544102 -336 544170
rect -956 544046 -860 544102
rect -804 544046 -736 544102
rect -680 544046 -612 544102
rect -556 544046 -488 544102
rect -432 544046 -336 544102
rect -956 543978 -336 544046
rect -956 543922 -860 543978
rect -804 543922 -736 543978
rect -680 543922 -612 543978
rect -556 543922 -488 543978
rect -432 543922 -336 543978
rect -956 526350 -336 543922
rect -956 526294 -860 526350
rect -804 526294 -736 526350
rect -680 526294 -612 526350
rect -556 526294 -488 526350
rect -432 526294 -336 526350
rect -956 526226 -336 526294
rect -956 526170 -860 526226
rect -804 526170 -736 526226
rect -680 526170 -612 526226
rect -556 526170 -488 526226
rect -432 526170 -336 526226
rect -956 526102 -336 526170
rect -956 526046 -860 526102
rect -804 526046 -736 526102
rect -680 526046 -612 526102
rect -556 526046 -488 526102
rect -432 526046 -336 526102
rect -956 525978 -336 526046
rect -956 525922 -860 525978
rect -804 525922 -736 525978
rect -680 525922 -612 525978
rect -556 525922 -488 525978
rect -432 525922 -336 525978
rect -956 508350 -336 525922
rect -956 508294 -860 508350
rect -804 508294 -736 508350
rect -680 508294 -612 508350
rect -556 508294 -488 508350
rect -432 508294 -336 508350
rect -956 508226 -336 508294
rect -956 508170 -860 508226
rect -804 508170 -736 508226
rect -680 508170 -612 508226
rect -556 508170 -488 508226
rect -432 508170 -336 508226
rect -956 508102 -336 508170
rect -956 508046 -860 508102
rect -804 508046 -736 508102
rect -680 508046 -612 508102
rect -556 508046 -488 508102
rect -432 508046 -336 508102
rect -956 507978 -336 508046
rect -956 507922 -860 507978
rect -804 507922 -736 507978
rect -680 507922 -612 507978
rect -556 507922 -488 507978
rect -432 507922 -336 507978
rect -956 490350 -336 507922
rect -956 490294 -860 490350
rect -804 490294 -736 490350
rect -680 490294 -612 490350
rect -556 490294 -488 490350
rect -432 490294 -336 490350
rect -956 490226 -336 490294
rect -956 490170 -860 490226
rect -804 490170 -736 490226
rect -680 490170 -612 490226
rect -556 490170 -488 490226
rect -432 490170 -336 490226
rect -956 490102 -336 490170
rect -956 490046 -860 490102
rect -804 490046 -736 490102
rect -680 490046 -612 490102
rect -556 490046 -488 490102
rect -432 490046 -336 490102
rect -956 489978 -336 490046
rect -956 489922 -860 489978
rect -804 489922 -736 489978
rect -680 489922 -612 489978
rect -556 489922 -488 489978
rect -432 489922 -336 489978
rect -956 472350 -336 489922
rect -956 472294 -860 472350
rect -804 472294 -736 472350
rect -680 472294 -612 472350
rect -556 472294 -488 472350
rect -432 472294 -336 472350
rect -956 472226 -336 472294
rect -956 472170 -860 472226
rect -804 472170 -736 472226
rect -680 472170 -612 472226
rect -556 472170 -488 472226
rect -432 472170 -336 472226
rect -956 472102 -336 472170
rect -956 472046 -860 472102
rect -804 472046 -736 472102
rect -680 472046 -612 472102
rect -556 472046 -488 472102
rect -432 472046 -336 472102
rect -956 471978 -336 472046
rect -956 471922 -860 471978
rect -804 471922 -736 471978
rect -680 471922 -612 471978
rect -556 471922 -488 471978
rect -432 471922 -336 471978
rect -956 454350 -336 471922
rect -956 454294 -860 454350
rect -804 454294 -736 454350
rect -680 454294 -612 454350
rect -556 454294 -488 454350
rect -432 454294 -336 454350
rect -956 454226 -336 454294
rect -956 454170 -860 454226
rect -804 454170 -736 454226
rect -680 454170 -612 454226
rect -556 454170 -488 454226
rect -432 454170 -336 454226
rect -956 454102 -336 454170
rect -956 454046 -860 454102
rect -804 454046 -736 454102
rect -680 454046 -612 454102
rect -556 454046 -488 454102
rect -432 454046 -336 454102
rect -956 453978 -336 454046
rect -956 453922 -860 453978
rect -804 453922 -736 453978
rect -680 453922 -612 453978
rect -556 453922 -488 453978
rect -432 453922 -336 453978
rect -956 436350 -336 453922
rect -956 436294 -860 436350
rect -804 436294 -736 436350
rect -680 436294 -612 436350
rect -556 436294 -488 436350
rect -432 436294 -336 436350
rect -956 436226 -336 436294
rect -956 436170 -860 436226
rect -804 436170 -736 436226
rect -680 436170 -612 436226
rect -556 436170 -488 436226
rect -432 436170 -336 436226
rect -956 436102 -336 436170
rect -956 436046 -860 436102
rect -804 436046 -736 436102
rect -680 436046 -612 436102
rect -556 436046 -488 436102
rect -432 436046 -336 436102
rect -956 435978 -336 436046
rect -956 435922 -860 435978
rect -804 435922 -736 435978
rect -680 435922 -612 435978
rect -556 435922 -488 435978
rect -432 435922 -336 435978
rect -956 418350 -336 435922
rect -956 418294 -860 418350
rect -804 418294 -736 418350
rect -680 418294 -612 418350
rect -556 418294 -488 418350
rect -432 418294 -336 418350
rect -956 418226 -336 418294
rect -956 418170 -860 418226
rect -804 418170 -736 418226
rect -680 418170 -612 418226
rect -556 418170 -488 418226
rect -432 418170 -336 418226
rect -956 418102 -336 418170
rect -956 418046 -860 418102
rect -804 418046 -736 418102
rect -680 418046 -612 418102
rect -556 418046 -488 418102
rect -432 418046 -336 418102
rect -956 417978 -336 418046
rect -956 417922 -860 417978
rect -804 417922 -736 417978
rect -680 417922 -612 417978
rect -556 417922 -488 417978
rect -432 417922 -336 417978
rect -956 400350 -336 417922
rect -956 400294 -860 400350
rect -804 400294 -736 400350
rect -680 400294 -612 400350
rect -556 400294 -488 400350
rect -432 400294 -336 400350
rect -956 400226 -336 400294
rect -956 400170 -860 400226
rect -804 400170 -736 400226
rect -680 400170 -612 400226
rect -556 400170 -488 400226
rect -432 400170 -336 400226
rect -956 400102 -336 400170
rect -956 400046 -860 400102
rect -804 400046 -736 400102
rect -680 400046 -612 400102
rect -556 400046 -488 400102
rect -432 400046 -336 400102
rect -956 399978 -336 400046
rect -956 399922 -860 399978
rect -804 399922 -736 399978
rect -680 399922 -612 399978
rect -556 399922 -488 399978
rect -432 399922 -336 399978
rect -956 382350 -336 399922
rect -956 382294 -860 382350
rect -804 382294 -736 382350
rect -680 382294 -612 382350
rect -556 382294 -488 382350
rect -432 382294 -336 382350
rect -956 382226 -336 382294
rect -956 382170 -860 382226
rect -804 382170 -736 382226
rect -680 382170 -612 382226
rect -556 382170 -488 382226
rect -432 382170 -336 382226
rect -956 382102 -336 382170
rect -956 382046 -860 382102
rect -804 382046 -736 382102
rect -680 382046 -612 382102
rect -556 382046 -488 382102
rect -432 382046 -336 382102
rect -956 381978 -336 382046
rect -956 381922 -860 381978
rect -804 381922 -736 381978
rect -680 381922 -612 381978
rect -556 381922 -488 381978
rect -432 381922 -336 381978
rect -956 364350 -336 381922
rect -956 364294 -860 364350
rect -804 364294 -736 364350
rect -680 364294 -612 364350
rect -556 364294 -488 364350
rect -432 364294 -336 364350
rect -956 364226 -336 364294
rect -956 364170 -860 364226
rect -804 364170 -736 364226
rect -680 364170 -612 364226
rect -556 364170 -488 364226
rect -432 364170 -336 364226
rect -956 364102 -336 364170
rect -956 364046 -860 364102
rect -804 364046 -736 364102
rect -680 364046 -612 364102
rect -556 364046 -488 364102
rect -432 364046 -336 364102
rect -956 363978 -336 364046
rect -956 363922 -860 363978
rect -804 363922 -736 363978
rect -680 363922 -612 363978
rect -556 363922 -488 363978
rect -432 363922 -336 363978
rect -956 346350 -336 363922
rect -956 346294 -860 346350
rect -804 346294 -736 346350
rect -680 346294 -612 346350
rect -556 346294 -488 346350
rect -432 346294 -336 346350
rect -956 346226 -336 346294
rect -956 346170 -860 346226
rect -804 346170 -736 346226
rect -680 346170 -612 346226
rect -556 346170 -488 346226
rect -432 346170 -336 346226
rect -956 346102 -336 346170
rect -956 346046 -860 346102
rect -804 346046 -736 346102
rect -680 346046 -612 346102
rect -556 346046 -488 346102
rect -432 346046 -336 346102
rect -956 345978 -336 346046
rect -956 345922 -860 345978
rect -804 345922 -736 345978
rect -680 345922 -612 345978
rect -556 345922 -488 345978
rect -432 345922 -336 345978
rect -956 328350 -336 345922
rect -956 328294 -860 328350
rect -804 328294 -736 328350
rect -680 328294 -612 328350
rect -556 328294 -488 328350
rect -432 328294 -336 328350
rect -956 328226 -336 328294
rect -956 328170 -860 328226
rect -804 328170 -736 328226
rect -680 328170 -612 328226
rect -556 328170 -488 328226
rect -432 328170 -336 328226
rect -956 328102 -336 328170
rect -956 328046 -860 328102
rect -804 328046 -736 328102
rect -680 328046 -612 328102
rect -556 328046 -488 328102
rect -432 328046 -336 328102
rect -956 327978 -336 328046
rect -956 327922 -860 327978
rect -804 327922 -736 327978
rect -680 327922 -612 327978
rect -556 327922 -488 327978
rect -432 327922 -336 327978
rect -956 310350 -336 327922
rect -956 310294 -860 310350
rect -804 310294 -736 310350
rect -680 310294 -612 310350
rect -556 310294 -488 310350
rect -432 310294 -336 310350
rect -956 310226 -336 310294
rect -956 310170 -860 310226
rect -804 310170 -736 310226
rect -680 310170 -612 310226
rect -556 310170 -488 310226
rect -432 310170 -336 310226
rect -956 310102 -336 310170
rect -956 310046 -860 310102
rect -804 310046 -736 310102
rect -680 310046 -612 310102
rect -556 310046 -488 310102
rect -432 310046 -336 310102
rect -956 309978 -336 310046
rect -956 309922 -860 309978
rect -804 309922 -736 309978
rect -680 309922 -612 309978
rect -556 309922 -488 309978
rect -432 309922 -336 309978
rect -956 292350 -336 309922
rect -956 292294 -860 292350
rect -804 292294 -736 292350
rect -680 292294 -612 292350
rect -556 292294 -488 292350
rect -432 292294 -336 292350
rect -956 292226 -336 292294
rect -956 292170 -860 292226
rect -804 292170 -736 292226
rect -680 292170 -612 292226
rect -556 292170 -488 292226
rect -432 292170 -336 292226
rect -956 292102 -336 292170
rect -956 292046 -860 292102
rect -804 292046 -736 292102
rect -680 292046 -612 292102
rect -556 292046 -488 292102
rect -432 292046 -336 292102
rect -956 291978 -336 292046
rect -956 291922 -860 291978
rect -804 291922 -736 291978
rect -680 291922 -612 291978
rect -556 291922 -488 291978
rect -432 291922 -336 291978
rect -956 274350 -336 291922
rect -956 274294 -860 274350
rect -804 274294 -736 274350
rect -680 274294 -612 274350
rect -556 274294 -488 274350
rect -432 274294 -336 274350
rect -956 274226 -336 274294
rect -956 274170 -860 274226
rect -804 274170 -736 274226
rect -680 274170 -612 274226
rect -556 274170 -488 274226
rect -432 274170 -336 274226
rect -956 274102 -336 274170
rect -956 274046 -860 274102
rect -804 274046 -736 274102
rect -680 274046 -612 274102
rect -556 274046 -488 274102
rect -432 274046 -336 274102
rect -956 273978 -336 274046
rect -956 273922 -860 273978
rect -804 273922 -736 273978
rect -680 273922 -612 273978
rect -556 273922 -488 273978
rect -432 273922 -336 273978
rect -956 256350 -336 273922
rect -956 256294 -860 256350
rect -804 256294 -736 256350
rect -680 256294 -612 256350
rect -556 256294 -488 256350
rect -432 256294 -336 256350
rect -956 256226 -336 256294
rect -956 256170 -860 256226
rect -804 256170 -736 256226
rect -680 256170 -612 256226
rect -556 256170 -488 256226
rect -432 256170 -336 256226
rect -956 256102 -336 256170
rect -956 256046 -860 256102
rect -804 256046 -736 256102
rect -680 256046 -612 256102
rect -556 256046 -488 256102
rect -432 256046 -336 256102
rect -956 255978 -336 256046
rect -956 255922 -860 255978
rect -804 255922 -736 255978
rect -680 255922 -612 255978
rect -556 255922 -488 255978
rect -432 255922 -336 255978
rect -956 238350 -336 255922
rect -956 238294 -860 238350
rect -804 238294 -736 238350
rect -680 238294 -612 238350
rect -556 238294 -488 238350
rect -432 238294 -336 238350
rect -956 238226 -336 238294
rect -956 238170 -860 238226
rect -804 238170 -736 238226
rect -680 238170 -612 238226
rect -556 238170 -488 238226
rect -432 238170 -336 238226
rect -956 238102 -336 238170
rect -956 238046 -860 238102
rect -804 238046 -736 238102
rect -680 238046 -612 238102
rect -556 238046 -488 238102
rect -432 238046 -336 238102
rect -956 237978 -336 238046
rect -956 237922 -860 237978
rect -804 237922 -736 237978
rect -680 237922 -612 237978
rect -556 237922 -488 237978
rect -432 237922 -336 237978
rect -956 220350 -336 237922
rect -956 220294 -860 220350
rect -804 220294 -736 220350
rect -680 220294 -612 220350
rect -556 220294 -488 220350
rect -432 220294 -336 220350
rect -956 220226 -336 220294
rect -956 220170 -860 220226
rect -804 220170 -736 220226
rect -680 220170 -612 220226
rect -556 220170 -488 220226
rect -432 220170 -336 220226
rect -956 220102 -336 220170
rect -956 220046 -860 220102
rect -804 220046 -736 220102
rect -680 220046 -612 220102
rect -556 220046 -488 220102
rect -432 220046 -336 220102
rect -956 219978 -336 220046
rect -956 219922 -860 219978
rect -804 219922 -736 219978
rect -680 219922 -612 219978
rect -556 219922 -488 219978
rect -432 219922 -336 219978
rect -956 202350 -336 219922
rect -956 202294 -860 202350
rect -804 202294 -736 202350
rect -680 202294 -612 202350
rect -556 202294 -488 202350
rect -432 202294 -336 202350
rect -956 202226 -336 202294
rect -956 202170 -860 202226
rect -804 202170 -736 202226
rect -680 202170 -612 202226
rect -556 202170 -488 202226
rect -432 202170 -336 202226
rect -956 202102 -336 202170
rect -956 202046 -860 202102
rect -804 202046 -736 202102
rect -680 202046 -612 202102
rect -556 202046 -488 202102
rect -432 202046 -336 202102
rect -956 201978 -336 202046
rect -956 201922 -860 201978
rect -804 201922 -736 201978
rect -680 201922 -612 201978
rect -556 201922 -488 201978
rect -432 201922 -336 201978
rect -956 184350 -336 201922
rect -956 184294 -860 184350
rect -804 184294 -736 184350
rect -680 184294 -612 184350
rect -556 184294 -488 184350
rect -432 184294 -336 184350
rect -956 184226 -336 184294
rect -956 184170 -860 184226
rect -804 184170 -736 184226
rect -680 184170 -612 184226
rect -556 184170 -488 184226
rect -432 184170 -336 184226
rect -956 184102 -336 184170
rect -956 184046 -860 184102
rect -804 184046 -736 184102
rect -680 184046 -612 184102
rect -556 184046 -488 184102
rect -432 184046 -336 184102
rect -956 183978 -336 184046
rect -956 183922 -860 183978
rect -804 183922 -736 183978
rect -680 183922 -612 183978
rect -556 183922 -488 183978
rect -432 183922 -336 183978
rect -956 166350 -336 183922
rect -956 166294 -860 166350
rect -804 166294 -736 166350
rect -680 166294 -612 166350
rect -556 166294 -488 166350
rect -432 166294 -336 166350
rect -956 166226 -336 166294
rect -956 166170 -860 166226
rect -804 166170 -736 166226
rect -680 166170 -612 166226
rect -556 166170 -488 166226
rect -432 166170 -336 166226
rect -956 166102 -336 166170
rect -956 166046 -860 166102
rect -804 166046 -736 166102
rect -680 166046 -612 166102
rect -556 166046 -488 166102
rect -432 166046 -336 166102
rect -956 165978 -336 166046
rect -956 165922 -860 165978
rect -804 165922 -736 165978
rect -680 165922 -612 165978
rect -556 165922 -488 165978
rect -432 165922 -336 165978
rect -956 148350 -336 165922
rect -956 148294 -860 148350
rect -804 148294 -736 148350
rect -680 148294 -612 148350
rect -556 148294 -488 148350
rect -432 148294 -336 148350
rect -956 148226 -336 148294
rect -956 148170 -860 148226
rect -804 148170 -736 148226
rect -680 148170 -612 148226
rect -556 148170 -488 148226
rect -432 148170 -336 148226
rect -956 148102 -336 148170
rect -956 148046 -860 148102
rect -804 148046 -736 148102
rect -680 148046 -612 148102
rect -556 148046 -488 148102
rect -432 148046 -336 148102
rect -956 147978 -336 148046
rect -956 147922 -860 147978
rect -804 147922 -736 147978
rect -680 147922 -612 147978
rect -556 147922 -488 147978
rect -432 147922 -336 147978
rect -956 130350 -336 147922
rect -956 130294 -860 130350
rect -804 130294 -736 130350
rect -680 130294 -612 130350
rect -556 130294 -488 130350
rect -432 130294 -336 130350
rect -956 130226 -336 130294
rect -956 130170 -860 130226
rect -804 130170 -736 130226
rect -680 130170 -612 130226
rect -556 130170 -488 130226
rect -432 130170 -336 130226
rect -956 130102 -336 130170
rect -956 130046 -860 130102
rect -804 130046 -736 130102
rect -680 130046 -612 130102
rect -556 130046 -488 130102
rect -432 130046 -336 130102
rect -956 129978 -336 130046
rect -956 129922 -860 129978
rect -804 129922 -736 129978
rect -680 129922 -612 129978
rect -556 129922 -488 129978
rect -432 129922 -336 129978
rect -956 112350 -336 129922
rect -956 112294 -860 112350
rect -804 112294 -736 112350
rect -680 112294 -612 112350
rect -556 112294 -488 112350
rect -432 112294 -336 112350
rect -956 112226 -336 112294
rect -956 112170 -860 112226
rect -804 112170 -736 112226
rect -680 112170 -612 112226
rect -556 112170 -488 112226
rect -432 112170 -336 112226
rect -956 112102 -336 112170
rect -956 112046 -860 112102
rect -804 112046 -736 112102
rect -680 112046 -612 112102
rect -556 112046 -488 112102
rect -432 112046 -336 112102
rect -956 111978 -336 112046
rect -956 111922 -860 111978
rect -804 111922 -736 111978
rect -680 111922 -612 111978
rect -556 111922 -488 111978
rect -432 111922 -336 111978
rect -956 94350 -336 111922
rect -956 94294 -860 94350
rect -804 94294 -736 94350
rect -680 94294 -612 94350
rect -556 94294 -488 94350
rect -432 94294 -336 94350
rect -956 94226 -336 94294
rect -956 94170 -860 94226
rect -804 94170 -736 94226
rect -680 94170 -612 94226
rect -556 94170 -488 94226
rect -432 94170 -336 94226
rect -956 94102 -336 94170
rect -956 94046 -860 94102
rect -804 94046 -736 94102
rect -680 94046 -612 94102
rect -556 94046 -488 94102
rect -432 94046 -336 94102
rect -956 93978 -336 94046
rect -956 93922 -860 93978
rect -804 93922 -736 93978
rect -680 93922 -612 93978
rect -556 93922 -488 93978
rect -432 93922 -336 93978
rect -956 76350 -336 93922
rect -956 76294 -860 76350
rect -804 76294 -736 76350
rect -680 76294 -612 76350
rect -556 76294 -488 76350
rect -432 76294 -336 76350
rect -956 76226 -336 76294
rect -956 76170 -860 76226
rect -804 76170 -736 76226
rect -680 76170 -612 76226
rect -556 76170 -488 76226
rect -432 76170 -336 76226
rect -956 76102 -336 76170
rect -956 76046 -860 76102
rect -804 76046 -736 76102
rect -680 76046 -612 76102
rect -556 76046 -488 76102
rect -432 76046 -336 76102
rect -956 75978 -336 76046
rect -956 75922 -860 75978
rect -804 75922 -736 75978
rect -680 75922 -612 75978
rect -556 75922 -488 75978
rect -432 75922 -336 75978
rect -956 58350 -336 75922
rect -956 58294 -860 58350
rect -804 58294 -736 58350
rect -680 58294 -612 58350
rect -556 58294 -488 58350
rect -432 58294 -336 58350
rect -956 58226 -336 58294
rect -956 58170 -860 58226
rect -804 58170 -736 58226
rect -680 58170 -612 58226
rect -556 58170 -488 58226
rect -432 58170 -336 58226
rect -956 58102 -336 58170
rect -956 58046 -860 58102
rect -804 58046 -736 58102
rect -680 58046 -612 58102
rect -556 58046 -488 58102
rect -432 58046 -336 58102
rect -956 57978 -336 58046
rect -956 57922 -860 57978
rect -804 57922 -736 57978
rect -680 57922 -612 57978
rect -556 57922 -488 57978
rect -432 57922 -336 57978
rect -956 40350 -336 57922
rect -956 40294 -860 40350
rect -804 40294 -736 40350
rect -680 40294 -612 40350
rect -556 40294 -488 40350
rect -432 40294 -336 40350
rect -956 40226 -336 40294
rect -956 40170 -860 40226
rect -804 40170 -736 40226
rect -680 40170 -612 40226
rect -556 40170 -488 40226
rect -432 40170 -336 40226
rect -956 40102 -336 40170
rect -956 40046 -860 40102
rect -804 40046 -736 40102
rect -680 40046 -612 40102
rect -556 40046 -488 40102
rect -432 40046 -336 40102
rect -956 39978 -336 40046
rect -956 39922 -860 39978
rect -804 39922 -736 39978
rect -680 39922 -612 39978
rect -556 39922 -488 39978
rect -432 39922 -336 39978
rect -956 22350 -336 39922
rect -956 22294 -860 22350
rect -804 22294 -736 22350
rect -680 22294 -612 22350
rect -556 22294 -488 22350
rect -432 22294 -336 22350
rect -956 22226 -336 22294
rect -956 22170 -860 22226
rect -804 22170 -736 22226
rect -680 22170 -612 22226
rect -556 22170 -488 22226
rect -432 22170 -336 22226
rect -956 22102 -336 22170
rect -956 22046 -860 22102
rect -804 22046 -736 22102
rect -680 22046 -612 22102
rect -556 22046 -488 22102
rect -432 22046 -336 22102
rect -956 21978 -336 22046
rect -956 21922 -860 21978
rect -804 21922 -736 21978
rect -680 21922 -612 21978
rect -556 21922 -488 21978
rect -432 21922 -336 21978
rect -956 4350 -336 21922
rect -956 4294 -860 4350
rect -804 4294 -736 4350
rect -680 4294 -612 4350
rect -556 4294 -488 4350
rect -432 4294 -336 4350
rect -956 4226 -336 4294
rect -956 4170 -860 4226
rect -804 4170 -736 4226
rect -680 4170 -612 4226
rect -556 4170 -488 4226
rect -432 4170 -336 4226
rect -956 4102 -336 4170
rect -956 4046 -860 4102
rect -804 4046 -736 4102
rect -680 4046 -612 4102
rect -556 4046 -488 4102
rect -432 4046 -336 4102
rect -956 3978 -336 4046
rect -956 3922 -860 3978
rect -804 3922 -736 3978
rect -680 3922 -612 3978
rect -556 3922 -488 3978
rect -432 3922 -336 3978
rect -956 -160 -336 3922
rect -956 -216 -860 -160
rect -804 -216 -736 -160
rect -680 -216 -612 -160
rect -556 -216 -488 -160
rect -432 -216 -336 -160
rect -956 -284 -336 -216
rect -956 -340 -860 -284
rect -804 -340 -736 -284
rect -680 -340 -612 -284
rect -556 -340 -488 -284
rect -432 -340 -336 -284
rect -956 -408 -336 -340
rect -956 -464 -860 -408
rect -804 -464 -736 -408
rect -680 -464 -612 -408
rect -556 -464 -488 -408
rect -432 -464 -336 -408
rect -956 -532 -336 -464
rect -956 -588 -860 -532
rect -804 -588 -736 -532
rect -680 -588 -612 -532
rect -556 -588 -488 -532
rect -432 -588 -336 -532
rect -956 -684 -336 -588
rect 3154 597212 3774 598268
rect 3154 597156 3250 597212
rect 3306 597156 3374 597212
rect 3430 597156 3498 597212
rect 3554 597156 3622 597212
rect 3678 597156 3774 597212
rect 3154 597088 3774 597156
rect 3154 597032 3250 597088
rect 3306 597032 3374 597088
rect 3430 597032 3498 597088
rect 3554 597032 3622 597088
rect 3678 597032 3774 597088
rect 3154 596964 3774 597032
rect 3154 596908 3250 596964
rect 3306 596908 3374 596964
rect 3430 596908 3498 596964
rect 3554 596908 3622 596964
rect 3678 596908 3774 596964
rect 3154 596840 3774 596908
rect 3154 596784 3250 596840
rect 3306 596784 3374 596840
rect 3430 596784 3498 596840
rect 3554 596784 3622 596840
rect 3678 596784 3774 596840
rect 3154 580350 3774 596784
rect 3154 580294 3250 580350
rect 3306 580294 3374 580350
rect 3430 580294 3498 580350
rect 3554 580294 3622 580350
rect 3678 580294 3774 580350
rect 3154 580226 3774 580294
rect 3154 580170 3250 580226
rect 3306 580170 3374 580226
rect 3430 580170 3498 580226
rect 3554 580170 3622 580226
rect 3678 580170 3774 580226
rect 3154 580102 3774 580170
rect 3154 580046 3250 580102
rect 3306 580046 3374 580102
rect 3430 580046 3498 580102
rect 3554 580046 3622 580102
rect 3678 580046 3774 580102
rect 3154 579978 3774 580046
rect 3154 579922 3250 579978
rect 3306 579922 3374 579978
rect 3430 579922 3498 579978
rect 3554 579922 3622 579978
rect 3678 579922 3774 579978
rect 3154 562350 3774 579922
rect 3154 562294 3250 562350
rect 3306 562294 3374 562350
rect 3430 562294 3498 562350
rect 3554 562294 3622 562350
rect 3678 562294 3774 562350
rect 3154 562226 3774 562294
rect 3154 562170 3250 562226
rect 3306 562170 3374 562226
rect 3430 562170 3498 562226
rect 3554 562170 3622 562226
rect 3678 562170 3774 562226
rect 3154 562102 3774 562170
rect 3154 562046 3250 562102
rect 3306 562046 3374 562102
rect 3430 562046 3498 562102
rect 3554 562046 3622 562102
rect 3678 562046 3774 562102
rect 3154 561978 3774 562046
rect 3154 561922 3250 561978
rect 3306 561922 3374 561978
rect 3430 561922 3498 561978
rect 3554 561922 3622 561978
rect 3678 561922 3774 561978
rect 3154 544350 3774 561922
rect 3154 544294 3250 544350
rect 3306 544294 3374 544350
rect 3430 544294 3498 544350
rect 3554 544294 3622 544350
rect 3678 544294 3774 544350
rect 3154 544226 3774 544294
rect 3154 544170 3250 544226
rect 3306 544170 3374 544226
rect 3430 544170 3498 544226
rect 3554 544170 3622 544226
rect 3678 544170 3774 544226
rect 3154 544102 3774 544170
rect 3154 544046 3250 544102
rect 3306 544046 3374 544102
rect 3430 544046 3498 544102
rect 3554 544046 3622 544102
rect 3678 544046 3774 544102
rect 3154 543978 3774 544046
rect 3154 543922 3250 543978
rect 3306 543922 3374 543978
rect 3430 543922 3498 543978
rect 3554 543922 3622 543978
rect 3678 543922 3774 543978
rect 3154 526350 3774 543922
rect 3154 526294 3250 526350
rect 3306 526294 3374 526350
rect 3430 526294 3498 526350
rect 3554 526294 3622 526350
rect 3678 526294 3774 526350
rect 3154 526226 3774 526294
rect 3154 526170 3250 526226
rect 3306 526170 3374 526226
rect 3430 526170 3498 526226
rect 3554 526170 3622 526226
rect 3678 526170 3774 526226
rect 3154 526102 3774 526170
rect 3154 526046 3250 526102
rect 3306 526046 3374 526102
rect 3430 526046 3498 526102
rect 3554 526046 3622 526102
rect 3678 526046 3774 526102
rect 3154 525978 3774 526046
rect 3154 525922 3250 525978
rect 3306 525922 3374 525978
rect 3430 525922 3498 525978
rect 3554 525922 3622 525978
rect 3678 525922 3774 525978
rect 3154 508350 3774 525922
rect 3154 508294 3250 508350
rect 3306 508294 3374 508350
rect 3430 508294 3498 508350
rect 3554 508294 3622 508350
rect 3678 508294 3774 508350
rect 3154 508226 3774 508294
rect 3154 508170 3250 508226
rect 3306 508170 3374 508226
rect 3430 508170 3498 508226
rect 3554 508170 3622 508226
rect 3678 508170 3774 508226
rect 3154 508102 3774 508170
rect 3154 508046 3250 508102
rect 3306 508046 3374 508102
rect 3430 508046 3498 508102
rect 3554 508046 3622 508102
rect 3678 508046 3774 508102
rect 3154 507978 3774 508046
rect 3154 507922 3250 507978
rect 3306 507922 3374 507978
rect 3430 507922 3498 507978
rect 3554 507922 3622 507978
rect 3678 507922 3774 507978
rect 3154 490350 3774 507922
rect 3154 490294 3250 490350
rect 3306 490294 3374 490350
rect 3430 490294 3498 490350
rect 3554 490294 3622 490350
rect 3678 490294 3774 490350
rect 3154 490226 3774 490294
rect 3154 490170 3250 490226
rect 3306 490170 3374 490226
rect 3430 490170 3498 490226
rect 3554 490170 3622 490226
rect 3678 490170 3774 490226
rect 3154 490102 3774 490170
rect 3154 490046 3250 490102
rect 3306 490046 3374 490102
rect 3430 490046 3498 490102
rect 3554 490046 3622 490102
rect 3678 490046 3774 490102
rect 3154 489978 3774 490046
rect 3154 489922 3250 489978
rect 3306 489922 3374 489978
rect 3430 489922 3498 489978
rect 3554 489922 3622 489978
rect 3678 489922 3774 489978
rect 3154 472350 3774 489922
rect 3154 472294 3250 472350
rect 3306 472294 3374 472350
rect 3430 472294 3498 472350
rect 3554 472294 3622 472350
rect 3678 472294 3774 472350
rect 3154 472226 3774 472294
rect 3154 472170 3250 472226
rect 3306 472170 3374 472226
rect 3430 472170 3498 472226
rect 3554 472170 3622 472226
rect 3678 472170 3774 472226
rect 3154 472102 3774 472170
rect 3154 472046 3250 472102
rect 3306 472046 3374 472102
rect 3430 472046 3498 472102
rect 3554 472046 3622 472102
rect 3678 472046 3774 472102
rect 3154 471978 3774 472046
rect 3154 471922 3250 471978
rect 3306 471922 3374 471978
rect 3430 471922 3498 471978
rect 3554 471922 3622 471978
rect 3678 471922 3774 471978
rect 3154 454350 3774 471922
rect 3154 454294 3250 454350
rect 3306 454294 3374 454350
rect 3430 454294 3498 454350
rect 3554 454294 3622 454350
rect 3678 454294 3774 454350
rect 3154 454226 3774 454294
rect 3154 454170 3250 454226
rect 3306 454170 3374 454226
rect 3430 454170 3498 454226
rect 3554 454170 3622 454226
rect 3678 454170 3774 454226
rect 3154 454102 3774 454170
rect 3154 454046 3250 454102
rect 3306 454046 3374 454102
rect 3430 454046 3498 454102
rect 3554 454046 3622 454102
rect 3678 454046 3774 454102
rect 3154 453978 3774 454046
rect 3154 453922 3250 453978
rect 3306 453922 3374 453978
rect 3430 453922 3498 453978
rect 3554 453922 3622 453978
rect 3678 453922 3774 453978
rect 3154 436350 3774 453922
rect 3154 436294 3250 436350
rect 3306 436294 3374 436350
rect 3430 436294 3498 436350
rect 3554 436294 3622 436350
rect 3678 436294 3774 436350
rect 3154 436226 3774 436294
rect 3154 436170 3250 436226
rect 3306 436170 3374 436226
rect 3430 436170 3498 436226
rect 3554 436170 3622 436226
rect 3678 436170 3774 436226
rect 3154 436102 3774 436170
rect 3154 436046 3250 436102
rect 3306 436046 3374 436102
rect 3430 436046 3498 436102
rect 3554 436046 3622 436102
rect 3678 436046 3774 436102
rect 3154 435978 3774 436046
rect 3154 435922 3250 435978
rect 3306 435922 3374 435978
rect 3430 435922 3498 435978
rect 3554 435922 3622 435978
rect 3678 435922 3774 435978
rect 3154 418350 3774 435922
rect 3154 418294 3250 418350
rect 3306 418294 3374 418350
rect 3430 418294 3498 418350
rect 3554 418294 3622 418350
rect 3678 418294 3774 418350
rect 3154 418226 3774 418294
rect 3154 418170 3250 418226
rect 3306 418170 3374 418226
rect 3430 418170 3498 418226
rect 3554 418170 3622 418226
rect 3678 418170 3774 418226
rect 3154 418102 3774 418170
rect 3154 418046 3250 418102
rect 3306 418046 3374 418102
rect 3430 418046 3498 418102
rect 3554 418046 3622 418102
rect 3678 418046 3774 418102
rect 3154 417978 3774 418046
rect 3154 417922 3250 417978
rect 3306 417922 3374 417978
rect 3430 417922 3498 417978
rect 3554 417922 3622 417978
rect 3678 417922 3774 417978
rect 3154 400350 3774 417922
rect 3154 400294 3250 400350
rect 3306 400294 3374 400350
rect 3430 400294 3498 400350
rect 3554 400294 3622 400350
rect 3678 400294 3774 400350
rect 3154 400226 3774 400294
rect 3154 400170 3250 400226
rect 3306 400170 3374 400226
rect 3430 400170 3498 400226
rect 3554 400170 3622 400226
rect 3678 400170 3774 400226
rect 3154 400102 3774 400170
rect 3154 400046 3250 400102
rect 3306 400046 3374 400102
rect 3430 400046 3498 400102
rect 3554 400046 3622 400102
rect 3678 400046 3774 400102
rect 3154 399978 3774 400046
rect 3154 399922 3250 399978
rect 3306 399922 3374 399978
rect 3430 399922 3498 399978
rect 3554 399922 3622 399978
rect 3678 399922 3774 399978
rect 3154 382350 3774 399922
rect 3154 382294 3250 382350
rect 3306 382294 3374 382350
rect 3430 382294 3498 382350
rect 3554 382294 3622 382350
rect 3678 382294 3774 382350
rect 3154 382226 3774 382294
rect 3154 382170 3250 382226
rect 3306 382170 3374 382226
rect 3430 382170 3498 382226
rect 3554 382170 3622 382226
rect 3678 382170 3774 382226
rect 3154 382102 3774 382170
rect 3154 382046 3250 382102
rect 3306 382046 3374 382102
rect 3430 382046 3498 382102
rect 3554 382046 3622 382102
rect 3678 382046 3774 382102
rect 3154 381978 3774 382046
rect 3154 381922 3250 381978
rect 3306 381922 3374 381978
rect 3430 381922 3498 381978
rect 3554 381922 3622 381978
rect 3678 381922 3774 381978
rect 3154 364350 3774 381922
rect 3154 364294 3250 364350
rect 3306 364294 3374 364350
rect 3430 364294 3498 364350
rect 3554 364294 3622 364350
rect 3678 364294 3774 364350
rect 3154 364226 3774 364294
rect 3154 364170 3250 364226
rect 3306 364170 3374 364226
rect 3430 364170 3498 364226
rect 3554 364170 3622 364226
rect 3678 364170 3774 364226
rect 3154 364102 3774 364170
rect 3154 364046 3250 364102
rect 3306 364046 3374 364102
rect 3430 364046 3498 364102
rect 3554 364046 3622 364102
rect 3678 364046 3774 364102
rect 3154 363978 3774 364046
rect 3154 363922 3250 363978
rect 3306 363922 3374 363978
rect 3430 363922 3498 363978
rect 3554 363922 3622 363978
rect 3678 363922 3774 363978
rect 3154 346350 3774 363922
rect 3154 346294 3250 346350
rect 3306 346294 3374 346350
rect 3430 346294 3498 346350
rect 3554 346294 3622 346350
rect 3678 346294 3774 346350
rect 3154 346226 3774 346294
rect 3154 346170 3250 346226
rect 3306 346170 3374 346226
rect 3430 346170 3498 346226
rect 3554 346170 3622 346226
rect 3678 346170 3774 346226
rect 3154 346102 3774 346170
rect 3154 346046 3250 346102
rect 3306 346046 3374 346102
rect 3430 346046 3498 346102
rect 3554 346046 3622 346102
rect 3678 346046 3774 346102
rect 3154 345978 3774 346046
rect 3154 345922 3250 345978
rect 3306 345922 3374 345978
rect 3430 345922 3498 345978
rect 3554 345922 3622 345978
rect 3678 345922 3774 345978
rect 3154 328350 3774 345922
rect 3154 328294 3250 328350
rect 3306 328294 3374 328350
rect 3430 328294 3498 328350
rect 3554 328294 3622 328350
rect 3678 328294 3774 328350
rect 3154 328226 3774 328294
rect 3154 328170 3250 328226
rect 3306 328170 3374 328226
rect 3430 328170 3498 328226
rect 3554 328170 3622 328226
rect 3678 328170 3774 328226
rect 3154 328102 3774 328170
rect 3154 328046 3250 328102
rect 3306 328046 3374 328102
rect 3430 328046 3498 328102
rect 3554 328046 3622 328102
rect 3678 328046 3774 328102
rect 3154 327978 3774 328046
rect 3154 327922 3250 327978
rect 3306 327922 3374 327978
rect 3430 327922 3498 327978
rect 3554 327922 3622 327978
rect 3678 327922 3774 327978
rect 3154 310350 3774 327922
rect 3154 310294 3250 310350
rect 3306 310294 3374 310350
rect 3430 310294 3498 310350
rect 3554 310294 3622 310350
rect 3678 310294 3774 310350
rect 3154 310226 3774 310294
rect 3154 310170 3250 310226
rect 3306 310170 3374 310226
rect 3430 310170 3498 310226
rect 3554 310170 3622 310226
rect 3678 310170 3774 310226
rect 3154 310102 3774 310170
rect 3154 310046 3250 310102
rect 3306 310046 3374 310102
rect 3430 310046 3498 310102
rect 3554 310046 3622 310102
rect 3678 310046 3774 310102
rect 3154 309978 3774 310046
rect 3154 309922 3250 309978
rect 3306 309922 3374 309978
rect 3430 309922 3498 309978
rect 3554 309922 3622 309978
rect 3678 309922 3774 309978
rect 3154 292350 3774 309922
rect 3154 292294 3250 292350
rect 3306 292294 3374 292350
rect 3430 292294 3498 292350
rect 3554 292294 3622 292350
rect 3678 292294 3774 292350
rect 3154 292226 3774 292294
rect 3154 292170 3250 292226
rect 3306 292170 3374 292226
rect 3430 292170 3498 292226
rect 3554 292170 3622 292226
rect 3678 292170 3774 292226
rect 3154 292102 3774 292170
rect 3154 292046 3250 292102
rect 3306 292046 3374 292102
rect 3430 292046 3498 292102
rect 3554 292046 3622 292102
rect 3678 292046 3774 292102
rect 3154 291978 3774 292046
rect 3154 291922 3250 291978
rect 3306 291922 3374 291978
rect 3430 291922 3498 291978
rect 3554 291922 3622 291978
rect 3678 291922 3774 291978
rect 3154 274350 3774 291922
rect 3154 274294 3250 274350
rect 3306 274294 3374 274350
rect 3430 274294 3498 274350
rect 3554 274294 3622 274350
rect 3678 274294 3774 274350
rect 3154 274226 3774 274294
rect 3154 274170 3250 274226
rect 3306 274170 3374 274226
rect 3430 274170 3498 274226
rect 3554 274170 3622 274226
rect 3678 274170 3774 274226
rect 3154 274102 3774 274170
rect 3154 274046 3250 274102
rect 3306 274046 3374 274102
rect 3430 274046 3498 274102
rect 3554 274046 3622 274102
rect 3678 274046 3774 274102
rect 3154 273978 3774 274046
rect 3154 273922 3250 273978
rect 3306 273922 3374 273978
rect 3430 273922 3498 273978
rect 3554 273922 3622 273978
rect 3678 273922 3774 273978
rect 3154 256350 3774 273922
rect 3154 256294 3250 256350
rect 3306 256294 3374 256350
rect 3430 256294 3498 256350
rect 3554 256294 3622 256350
rect 3678 256294 3774 256350
rect 3154 256226 3774 256294
rect 3154 256170 3250 256226
rect 3306 256170 3374 256226
rect 3430 256170 3498 256226
rect 3554 256170 3622 256226
rect 3678 256170 3774 256226
rect 3154 256102 3774 256170
rect 3154 256046 3250 256102
rect 3306 256046 3374 256102
rect 3430 256046 3498 256102
rect 3554 256046 3622 256102
rect 3678 256046 3774 256102
rect 3154 255978 3774 256046
rect 3154 255922 3250 255978
rect 3306 255922 3374 255978
rect 3430 255922 3498 255978
rect 3554 255922 3622 255978
rect 3678 255922 3774 255978
rect 3154 238350 3774 255922
rect 3154 238294 3250 238350
rect 3306 238294 3374 238350
rect 3430 238294 3498 238350
rect 3554 238294 3622 238350
rect 3678 238294 3774 238350
rect 3154 238226 3774 238294
rect 3154 238170 3250 238226
rect 3306 238170 3374 238226
rect 3430 238170 3498 238226
rect 3554 238170 3622 238226
rect 3678 238170 3774 238226
rect 3154 238102 3774 238170
rect 3154 238046 3250 238102
rect 3306 238046 3374 238102
rect 3430 238046 3498 238102
rect 3554 238046 3622 238102
rect 3678 238046 3774 238102
rect 3154 237978 3774 238046
rect 3154 237922 3250 237978
rect 3306 237922 3374 237978
rect 3430 237922 3498 237978
rect 3554 237922 3622 237978
rect 3678 237922 3774 237978
rect 3154 220350 3774 237922
rect 3154 220294 3250 220350
rect 3306 220294 3374 220350
rect 3430 220294 3498 220350
rect 3554 220294 3622 220350
rect 3678 220294 3774 220350
rect 3154 220226 3774 220294
rect 3154 220170 3250 220226
rect 3306 220170 3374 220226
rect 3430 220170 3498 220226
rect 3554 220170 3622 220226
rect 3678 220170 3774 220226
rect 3154 220102 3774 220170
rect 3154 220046 3250 220102
rect 3306 220046 3374 220102
rect 3430 220046 3498 220102
rect 3554 220046 3622 220102
rect 3678 220046 3774 220102
rect 3154 219978 3774 220046
rect 3154 219922 3250 219978
rect 3306 219922 3374 219978
rect 3430 219922 3498 219978
rect 3554 219922 3622 219978
rect 3678 219922 3774 219978
rect 3154 202350 3774 219922
rect 3154 202294 3250 202350
rect 3306 202294 3374 202350
rect 3430 202294 3498 202350
rect 3554 202294 3622 202350
rect 3678 202294 3774 202350
rect 3154 202226 3774 202294
rect 3154 202170 3250 202226
rect 3306 202170 3374 202226
rect 3430 202170 3498 202226
rect 3554 202170 3622 202226
rect 3678 202170 3774 202226
rect 3154 202102 3774 202170
rect 3154 202046 3250 202102
rect 3306 202046 3374 202102
rect 3430 202046 3498 202102
rect 3554 202046 3622 202102
rect 3678 202046 3774 202102
rect 3154 201978 3774 202046
rect 3154 201922 3250 201978
rect 3306 201922 3374 201978
rect 3430 201922 3498 201978
rect 3554 201922 3622 201978
rect 3678 201922 3774 201978
rect 3154 184350 3774 201922
rect 3154 184294 3250 184350
rect 3306 184294 3374 184350
rect 3430 184294 3498 184350
rect 3554 184294 3622 184350
rect 3678 184294 3774 184350
rect 3154 184226 3774 184294
rect 3154 184170 3250 184226
rect 3306 184170 3374 184226
rect 3430 184170 3498 184226
rect 3554 184170 3622 184226
rect 3678 184170 3774 184226
rect 3154 184102 3774 184170
rect 3154 184046 3250 184102
rect 3306 184046 3374 184102
rect 3430 184046 3498 184102
rect 3554 184046 3622 184102
rect 3678 184046 3774 184102
rect 3154 183978 3774 184046
rect 3154 183922 3250 183978
rect 3306 183922 3374 183978
rect 3430 183922 3498 183978
rect 3554 183922 3622 183978
rect 3678 183922 3774 183978
rect 3154 166350 3774 183922
rect 3154 166294 3250 166350
rect 3306 166294 3374 166350
rect 3430 166294 3498 166350
rect 3554 166294 3622 166350
rect 3678 166294 3774 166350
rect 3154 166226 3774 166294
rect 3154 166170 3250 166226
rect 3306 166170 3374 166226
rect 3430 166170 3498 166226
rect 3554 166170 3622 166226
rect 3678 166170 3774 166226
rect 3154 166102 3774 166170
rect 3154 166046 3250 166102
rect 3306 166046 3374 166102
rect 3430 166046 3498 166102
rect 3554 166046 3622 166102
rect 3678 166046 3774 166102
rect 3154 165978 3774 166046
rect 3154 165922 3250 165978
rect 3306 165922 3374 165978
rect 3430 165922 3498 165978
rect 3554 165922 3622 165978
rect 3678 165922 3774 165978
rect 3154 148350 3774 165922
rect 3154 148294 3250 148350
rect 3306 148294 3374 148350
rect 3430 148294 3498 148350
rect 3554 148294 3622 148350
rect 3678 148294 3774 148350
rect 3154 148226 3774 148294
rect 3154 148170 3250 148226
rect 3306 148170 3374 148226
rect 3430 148170 3498 148226
rect 3554 148170 3622 148226
rect 3678 148170 3774 148226
rect 3154 148102 3774 148170
rect 3154 148046 3250 148102
rect 3306 148046 3374 148102
rect 3430 148046 3498 148102
rect 3554 148046 3622 148102
rect 3678 148046 3774 148102
rect 3154 147978 3774 148046
rect 3154 147922 3250 147978
rect 3306 147922 3374 147978
rect 3430 147922 3498 147978
rect 3554 147922 3622 147978
rect 3678 147922 3774 147978
rect 3154 130350 3774 147922
rect 3154 130294 3250 130350
rect 3306 130294 3374 130350
rect 3430 130294 3498 130350
rect 3554 130294 3622 130350
rect 3678 130294 3774 130350
rect 3154 130226 3774 130294
rect 3154 130170 3250 130226
rect 3306 130170 3374 130226
rect 3430 130170 3498 130226
rect 3554 130170 3622 130226
rect 3678 130170 3774 130226
rect 3154 130102 3774 130170
rect 3154 130046 3250 130102
rect 3306 130046 3374 130102
rect 3430 130046 3498 130102
rect 3554 130046 3622 130102
rect 3678 130046 3774 130102
rect 3154 129978 3774 130046
rect 3154 129922 3250 129978
rect 3306 129922 3374 129978
rect 3430 129922 3498 129978
rect 3554 129922 3622 129978
rect 3678 129922 3774 129978
rect 3154 112350 3774 129922
rect 3154 112294 3250 112350
rect 3306 112294 3374 112350
rect 3430 112294 3498 112350
rect 3554 112294 3622 112350
rect 3678 112294 3774 112350
rect 3154 112226 3774 112294
rect 3154 112170 3250 112226
rect 3306 112170 3374 112226
rect 3430 112170 3498 112226
rect 3554 112170 3622 112226
rect 3678 112170 3774 112226
rect 3154 112102 3774 112170
rect 3154 112046 3250 112102
rect 3306 112046 3374 112102
rect 3430 112046 3498 112102
rect 3554 112046 3622 112102
rect 3678 112046 3774 112102
rect 3154 111978 3774 112046
rect 3154 111922 3250 111978
rect 3306 111922 3374 111978
rect 3430 111922 3498 111978
rect 3554 111922 3622 111978
rect 3678 111922 3774 111978
rect 3154 94350 3774 111922
rect 3154 94294 3250 94350
rect 3306 94294 3374 94350
rect 3430 94294 3498 94350
rect 3554 94294 3622 94350
rect 3678 94294 3774 94350
rect 3154 94226 3774 94294
rect 3154 94170 3250 94226
rect 3306 94170 3374 94226
rect 3430 94170 3498 94226
rect 3554 94170 3622 94226
rect 3678 94170 3774 94226
rect 3154 94102 3774 94170
rect 3154 94046 3250 94102
rect 3306 94046 3374 94102
rect 3430 94046 3498 94102
rect 3554 94046 3622 94102
rect 3678 94046 3774 94102
rect 3154 93978 3774 94046
rect 3154 93922 3250 93978
rect 3306 93922 3374 93978
rect 3430 93922 3498 93978
rect 3554 93922 3622 93978
rect 3678 93922 3774 93978
rect 3154 76350 3774 93922
rect 3154 76294 3250 76350
rect 3306 76294 3374 76350
rect 3430 76294 3498 76350
rect 3554 76294 3622 76350
rect 3678 76294 3774 76350
rect 3154 76226 3774 76294
rect 3154 76170 3250 76226
rect 3306 76170 3374 76226
rect 3430 76170 3498 76226
rect 3554 76170 3622 76226
rect 3678 76170 3774 76226
rect 3154 76102 3774 76170
rect 3154 76046 3250 76102
rect 3306 76046 3374 76102
rect 3430 76046 3498 76102
rect 3554 76046 3622 76102
rect 3678 76046 3774 76102
rect 3154 75978 3774 76046
rect 3154 75922 3250 75978
rect 3306 75922 3374 75978
rect 3430 75922 3498 75978
rect 3554 75922 3622 75978
rect 3678 75922 3774 75978
rect 3154 58350 3774 75922
rect 3154 58294 3250 58350
rect 3306 58294 3374 58350
rect 3430 58294 3498 58350
rect 3554 58294 3622 58350
rect 3678 58294 3774 58350
rect 3154 58226 3774 58294
rect 3154 58170 3250 58226
rect 3306 58170 3374 58226
rect 3430 58170 3498 58226
rect 3554 58170 3622 58226
rect 3678 58170 3774 58226
rect 3154 58102 3774 58170
rect 3154 58046 3250 58102
rect 3306 58046 3374 58102
rect 3430 58046 3498 58102
rect 3554 58046 3622 58102
rect 3678 58046 3774 58102
rect 3154 57978 3774 58046
rect 3154 57922 3250 57978
rect 3306 57922 3374 57978
rect 3430 57922 3498 57978
rect 3554 57922 3622 57978
rect 3678 57922 3774 57978
rect 3154 40350 3774 57922
rect 3154 40294 3250 40350
rect 3306 40294 3374 40350
rect 3430 40294 3498 40350
rect 3554 40294 3622 40350
rect 3678 40294 3774 40350
rect 3154 40226 3774 40294
rect 3154 40170 3250 40226
rect 3306 40170 3374 40226
rect 3430 40170 3498 40226
rect 3554 40170 3622 40226
rect 3678 40170 3774 40226
rect 3154 40102 3774 40170
rect 3154 40046 3250 40102
rect 3306 40046 3374 40102
rect 3430 40046 3498 40102
rect 3554 40046 3622 40102
rect 3678 40046 3774 40102
rect 3154 39978 3774 40046
rect 3154 39922 3250 39978
rect 3306 39922 3374 39978
rect 3430 39922 3498 39978
rect 3554 39922 3622 39978
rect 3678 39922 3774 39978
rect 3154 22350 3774 39922
rect 3154 22294 3250 22350
rect 3306 22294 3374 22350
rect 3430 22294 3498 22350
rect 3554 22294 3622 22350
rect 3678 22294 3774 22350
rect 3154 22226 3774 22294
rect 3154 22170 3250 22226
rect 3306 22170 3374 22226
rect 3430 22170 3498 22226
rect 3554 22170 3622 22226
rect 3678 22170 3774 22226
rect 3154 22102 3774 22170
rect 3154 22046 3250 22102
rect 3306 22046 3374 22102
rect 3430 22046 3498 22102
rect 3554 22046 3622 22102
rect 3678 22046 3774 22102
rect 3154 21978 3774 22046
rect 3154 21922 3250 21978
rect 3306 21922 3374 21978
rect 3430 21922 3498 21978
rect 3554 21922 3622 21978
rect 3678 21922 3774 21978
rect 3154 4350 3774 21922
rect 3154 4294 3250 4350
rect 3306 4294 3374 4350
rect 3430 4294 3498 4350
rect 3554 4294 3622 4350
rect 3678 4294 3774 4350
rect 3154 4226 3774 4294
rect 3154 4170 3250 4226
rect 3306 4170 3374 4226
rect 3430 4170 3498 4226
rect 3554 4170 3622 4226
rect 3678 4170 3774 4226
rect 3154 4102 3774 4170
rect 3154 4046 3250 4102
rect 3306 4046 3374 4102
rect 3430 4046 3498 4102
rect 3554 4046 3622 4102
rect 3678 4046 3774 4102
rect 3154 3978 3774 4046
rect 3154 3922 3250 3978
rect 3306 3922 3374 3978
rect 3430 3922 3498 3978
rect 3554 3922 3622 3978
rect 3678 3922 3774 3978
rect 3154 -160 3774 3922
rect 3154 -216 3250 -160
rect 3306 -216 3374 -160
rect 3430 -216 3498 -160
rect 3554 -216 3622 -160
rect 3678 -216 3774 -160
rect 3154 -284 3774 -216
rect 3154 -340 3250 -284
rect 3306 -340 3374 -284
rect 3430 -340 3498 -284
rect 3554 -340 3622 -284
rect 3678 -340 3774 -284
rect 3154 -408 3774 -340
rect 3154 -464 3250 -408
rect 3306 -464 3374 -408
rect 3430 -464 3498 -408
rect 3554 -464 3622 -408
rect 3678 -464 3774 -408
rect 3154 -532 3774 -464
rect 3154 -588 3250 -532
rect 3306 -588 3374 -532
rect 3430 -588 3498 -532
rect 3554 -588 3622 -532
rect 3678 -588 3774 -532
rect -1916 -1176 -1820 -1120
rect -1764 -1176 -1696 -1120
rect -1640 -1176 -1572 -1120
rect -1516 -1176 -1448 -1120
rect -1392 -1176 -1296 -1120
rect -1916 -1244 -1296 -1176
rect -1916 -1300 -1820 -1244
rect -1764 -1300 -1696 -1244
rect -1640 -1300 -1572 -1244
rect -1516 -1300 -1448 -1244
rect -1392 -1300 -1296 -1244
rect -1916 -1368 -1296 -1300
rect -1916 -1424 -1820 -1368
rect -1764 -1424 -1696 -1368
rect -1640 -1424 -1572 -1368
rect -1516 -1424 -1448 -1368
rect -1392 -1424 -1296 -1368
rect -1916 -1492 -1296 -1424
rect -1916 -1548 -1820 -1492
rect -1764 -1548 -1696 -1492
rect -1640 -1548 -1572 -1492
rect -1516 -1548 -1448 -1492
rect -1392 -1548 -1296 -1492
rect -1916 -1644 -1296 -1548
rect 3154 -1644 3774 -588
rect 6874 598172 7494 598268
rect 6874 598116 6970 598172
rect 7026 598116 7094 598172
rect 7150 598116 7218 598172
rect 7274 598116 7342 598172
rect 7398 598116 7494 598172
rect 6874 598048 7494 598116
rect 6874 597992 6970 598048
rect 7026 597992 7094 598048
rect 7150 597992 7218 598048
rect 7274 597992 7342 598048
rect 7398 597992 7494 598048
rect 6874 597924 7494 597992
rect 6874 597868 6970 597924
rect 7026 597868 7094 597924
rect 7150 597868 7218 597924
rect 7274 597868 7342 597924
rect 7398 597868 7494 597924
rect 6874 597800 7494 597868
rect 6874 597744 6970 597800
rect 7026 597744 7094 597800
rect 7150 597744 7218 597800
rect 7274 597744 7342 597800
rect 7398 597744 7494 597800
rect 6874 586350 7494 597744
rect 21154 597212 21774 598268
rect 21154 597156 21250 597212
rect 21306 597156 21374 597212
rect 21430 597156 21498 597212
rect 21554 597156 21622 597212
rect 21678 597156 21774 597212
rect 21154 597088 21774 597156
rect 21154 597032 21250 597088
rect 21306 597032 21374 597088
rect 21430 597032 21498 597088
rect 21554 597032 21622 597088
rect 21678 597032 21774 597088
rect 21154 596964 21774 597032
rect 21154 596908 21250 596964
rect 21306 596908 21374 596964
rect 21430 596908 21498 596964
rect 21554 596908 21622 596964
rect 21678 596908 21774 596964
rect 21154 596840 21774 596908
rect 21154 596784 21250 596840
rect 21306 596784 21374 596840
rect 21430 596784 21498 596840
rect 21554 596784 21622 596840
rect 21678 596784 21774 596840
rect 6874 586294 6970 586350
rect 7026 586294 7094 586350
rect 7150 586294 7218 586350
rect 7274 586294 7342 586350
rect 7398 586294 7494 586350
rect 6874 586226 7494 586294
rect 6874 586170 6970 586226
rect 7026 586170 7094 586226
rect 7150 586170 7218 586226
rect 7274 586170 7342 586226
rect 7398 586170 7494 586226
rect 6874 586102 7494 586170
rect 6874 586046 6970 586102
rect 7026 586046 7094 586102
rect 7150 586046 7218 586102
rect 7274 586046 7342 586102
rect 7398 586046 7494 586102
rect 6874 585978 7494 586046
rect 6874 585922 6970 585978
rect 7026 585922 7094 585978
rect 7150 585922 7218 585978
rect 7274 585922 7342 585978
rect 7398 585922 7494 585978
rect 6874 568350 7494 585922
rect 6874 568294 6970 568350
rect 7026 568294 7094 568350
rect 7150 568294 7218 568350
rect 7274 568294 7342 568350
rect 7398 568294 7494 568350
rect 6874 568226 7494 568294
rect 6874 568170 6970 568226
rect 7026 568170 7094 568226
rect 7150 568170 7218 568226
rect 7274 568170 7342 568226
rect 7398 568170 7494 568226
rect 6874 568102 7494 568170
rect 6874 568046 6970 568102
rect 7026 568046 7094 568102
rect 7150 568046 7218 568102
rect 7274 568046 7342 568102
rect 7398 568046 7494 568102
rect 6874 567978 7494 568046
rect 6874 567922 6970 567978
rect 7026 567922 7094 567978
rect 7150 567922 7218 567978
rect 7274 567922 7342 567978
rect 7398 567922 7494 567978
rect 6874 550350 7494 567922
rect 9996 587972 10052 587982
rect 6874 550294 6970 550350
rect 7026 550294 7094 550350
rect 7150 550294 7218 550350
rect 7274 550294 7342 550350
rect 7398 550294 7494 550350
rect 6874 550226 7494 550294
rect 6874 550170 6970 550226
rect 7026 550170 7094 550226
rect 7150 550170 7218 550226
rect 7274 550170 7342 550226
rect 7398 550170 7494 550226
rect 6874 550102 7494 550170
rect 6874 550046 6970 550102
rect 7026 550046 7094 550102
rect 7150 550046 7218 550102
rect 7274 550046 7342 550102
rect 7398 550046 7494 550102
rect 6874 549978 7494 550046
rect 6874 549922 6970 549978
rect 7026 549922 7094 549978
rect 7150 549922 7218 549978
rect 7274 549922 7342 549978
rect 7398 549922 7494 549978
rect 6874 532350 7494 549922
rect 6874 532294 6970 532350
rect 7026 532294 7094 532350
rect 7150 532294 7218 532350
rect 7274 532294 7342 532350
rect 7398 532294 7494 532350
rect 6874 532226 7494 532294
rect 6874 532170 6970 532226
rect 7026 532170 7094 532226
rect 7150 532170 7218 532226
rect 7274 532170 7342 532226
rect 7398 532170 7494 532226
rect 6874 532102 7494 532170
rect 6874 532046 6970 532102
rect 7026 532046 7094 532102
rect 7150 532046 7218 532102
rect 7274 532046 7342 532102
rect 7398 532046 7494 532102
rect 6874 531978 7494 532046
rect 6874 531922 6970 531978
rect 7026 531922 7094 531978
rect 7150 531922 7218 531978
rect 7274 531922 7342 531978
rect 7398 531922 7494 531978
rect 6874 514350 7494 531922
rect 6874 514294 6970 514350
rect 7026 514294 7094 514350
rect 7150 514294 7218 514350
rect 7274 514294 7342 514350
rect 7398 514294 7494 514350
rect 6874 514226 7494 514294
rect 6874 514170 6970 514226
rect 7026 514170 7094 514226
rect 7150 514170 7218 514226
rect 7274 514170 7342 514226
rect 7398 514170 7494 514226
rect 6874 514102 7494 514170
rect 6874 514046 6970 514102
rect 7026 514046 7094 514102
rect 7150 514046 7218 514102
rect 7274 514046 7342 514102
rect 7398 514046 7494 514102
rect 6874 513978 7494 514046
rect 6874 513922 6970 513978
rect 7026 513922 7094 513978
rect 7150 513922 7218 513978
rect 7274 513922 7342 513978
rect 7398 513922 7494 513978
rect 6874 496350 7494 513922
rect 6874 496294 6970 496350
rect 7026 496294 7094 496350
rect 7150 496294 7218 496350
rect 7274 496294 7342 496350
rect 7398 496294 7494 496350
rect 6874 496226 7494 496294
rect 6874 496170 6970 496226
rect 7026 496170 7094 496226
rect 7150 496170 7218 496226
rect 7274 496170 7342 496226
rect 7398 496170 7494 496226
rect 6874 496102 7494 496170
rect 6874 496046 6970 496102
rect 7026 496046 7094 496102
rect 7150 496046 7218 496102
rect 7274 496046 7342 496102
rect 7398 496046 7494 496102
rect 6874 495978 7494 496046
rect 6874 495922 6970 495978
rect 7026 495922 7094 495978
rect 7150 495922 7218 495978
rect 7274 495922 7342 495978
rect 7398 495922 7494 495978
rect 6874 478350 7494 495922
rect 6874 478294 6970 478350
rect 7026 478294 7094 478350
rect 7150 478294 7218 478350
rect 7274 478294 7342 478350
rect 7398 478294 7494 478350
rect 6874 478226 7494 478294
rect 6874 478170 6970 478226
rect 7026 478170 7094 478226
rect 7150 478170 7218 478226
rect 7274 478170 7342 478226
rect 7398 478170 7494 478226
rect 6874 478102 7494 478170
rect 6874 478046 6970 478102
rect 7026 478046 7094 478102
rect 7150 478046 7218 478102
rect 7274 478046 7342 478102
rect 7398 478046 7494 478102
rect 6874 477978 7494 478046
rect 6874 477922 6970 477978
rect 7026 477922 7094 477978
rect 7150 477922 7218 477978
rect 7274 477922 7342 477978
rect 7398 477922 7494 477978
rect 6874 460350 7494 477922
rect 6874 460294 6970 460350
rect 7026 460294 7094 460350
rect 7150 460294 7218 460350
rect 7274 460294 7342 460350
rect 7398 460294 7494 460350
rect 6874 460226 7494 460294
rect 6874 460170 6970 460226
rect 7026 460170 7094 460226
rect 7150 460170 7218 460226
rect 7274 460170 7342 460226
rect 7398 460170 7494 460226
rect 6874 460102 7494 460170
rect 6874 460046 6970 460102
rect 7026 460046 7094 460102
rect 7150 460046 7218 460102
rect 7274 460046 7342 460102
rect 7398 460046 7494 460102
rect 6874 459978 7494 460046
rect 6874 459922 6970 459978
rect 7026 459922 7094 459978
rect 7150 459922 7218 459978
rect 7274 459922 7342 459978
rect 7398 459922 7494 459978
rect 6874 442350 7494 459922
rect 6874 442294 6970 442350
rect 7026 442294 7094 442350
rect 7150 442294 7218 442350
rect 7274 442294 7342 442350
rect 7398 442294 7494 442350
rect 6874 442226 7494 442294
rect 6874 442170 6970 442226
rect 7026 442170 7094 442226
rect 7150 442170 7218 442226
rect 7274 442170 7342 442226
rect 7398 442170 7494 442226
rect 6874 442102 7494 442170
rect 6874 442046 6970 442102
rect 7026 442046 7094 442102
rect 7150 442046 7218 442102
rect 7274 442046 7342 442102
rect 7398 442046 7494 442102
rect 6874 441978 7494 442046
rect 6874 441922 6970 441978
rect 7026 441922 7094 441978
rect 7150 441922 7218 441978
rect 7274 441922 7342 441978
rect 7398 441922 7494 441978
rect 6874 424350 7494 441922
rect 6874 424294 6970 424350
rect 7026 424294 7094 424350
rect 7150 424294 7218 424350
rect 7274 424294 7342 424350
rect 7398 424294 7494 424350
rect 6874 424226 7494 424294
rect 6874 424170 6970 424226
rect 7026 424170 7094 424226
rect 7150 424170 7218 424226
rect 7274 424170 7342 424226
rect 7398 424170 7494 424226
rect 6874 424102 7494 424170
rect 6874 424046 6970 424102
rect 7026 424046 7094 424102
rect 7150 424046 7218 424102
rect 7274 424046 7342 424102
rect 7398 424046 7494 424102
rect 6874 423978 7494 424046
rect 6874 423922 6970 423978
rect 7026 423922 7094 423978
rect 7150 423922 7218 423978
rect 7274 423922 7342 423978
rect 7398 423922 7494 423978
rect 6874 406350 7494 423922
rect 6874 406294 6970 406350
rect 7026 406294 7094 406350
rect 7150 406294 7218 406350
rect 7274 406294 7342 406350
rect 7398 406294 7494 406350
rect 6874 406226 7494 406294
rect 6874 406170 6970 406226
rect 7026 406170 7094 406226
rect 7150 406170 7218 406226
rect 7274 406170 7342 406226
rect 7398 406170 7494 406226
rect 6874 406102 7494 406170
rect 6874 406046 6970 406102
rect 7026 406046 7094 406102
rect 7150 406046 7218 406102
rect 7274 406046 7342 406102
rect 7398 406046 7494 406102
rect 6874 405978 7494 406046
rect 6874 405922 6970 405978
rect 7026 405922 7094 405978
rect 7150 405922 7218 405978
rect 7274 405922 7342 405978
rect 7398 405922 7494 405978
rect 6874 388350 7494 405922
rect 6874 388294 6970 388350
rect 7026 388294 7094 388350
rect 7150 388294 7218 388350
rect 7274 388294 7342 388350
rect 7398 388294 7494 388350
rect 6874 388226 7494 388294
rect 6874 388170 6970 388226
rect 7026 388170 7094 388226
rect 7150 388170 7218 388226
rect 7274 388170 7342 388226
rect 7398 388170 7494 388226
rect 6874 388102 7494 388170
rect 6874 388046 6970 388102
rect 7026 388046 7094 388102
rect 7150 388046 7218 388102
rect 7274 388046 7342 388102
rect 7398 388046 7494 388102
rect 6874 387978 7494 388046
rect 6874 387922 6970 387978
rect 7026 387922 7094 387978
rect 7150 387922 7218 387978
rect 7274 387922 7342 387978
rect 7398 387922 7494 387978
rect 6874 370350 7494 387922
rect 6874 370294 6970 370350
rect 7026 370294 7094 370350
rect 7150 370294 7218 370350
rect 7274 370294 7342 370350
rect 7398 370294 7494 370350
rect 6874 370226 7494 370294
rect 6874 370170 6970 370226
rect 7026 370170 7094 370226
rect 7150 370170 7218 370226
rect 7274 370170 7342 370226
rect 7398 370170 7494 370226
rect 6874 370102 7494 370170
rect 6874 370046 6970 370102
rect 7026 370046 7094 370102
rect 7150 370046 7218 370102
rect 7274 370046 7342 370102
rect 7398 370046 7494 370102
rect 6874 369978 7494 370046
rect 6874 369922 6970 369978
rect 7026 369922 7094 369978
rect 7150 369922 7218 369978
rect 7274 369922 7342 369978
rect 7398 369922 7494 369978
rect 6874 352350 7494 369922
rect 6874 352294 6970 352350
rect 7026 352294 7094 352350
rect 7150 352294 7218 352350
rect 7274 352294 7342 352350
rect 7398 352294 7494 352350
rect 6874 352226 7494 352294
rect 6874 352170 6970 352226
rect 7026 352170 7094 352226
rect 7150 352170 7218 352226
rect 7274 352170 7342 352226
rect 7398 352170 7494 352226
rect 6874 352102 7494 352170
rect 6874 352046 6970 352102
rect 7026 352046 7094 352102
rect 7150 352046 7218 352102
rect 7274 352046 7342 352102
rect 7398 352046 7494 352102
rect 6874 351978 7494 352046
rect 6874 351922 6970 351978
rect 7026 351922 7094 351978
rect 7150 351922 7218 351978
rect 7274 351922 7342 351978
rect 7398 351922 7494 351978
rect 6874 334350 7494 351922
rect 6874 334294 6970 334350
rect 7026 334294 7094 334350
rect 7150 334294 7218 334350
rect 7274 334294 7342 334350
rect 7398 334294 7494 334350
rect 6874 334226 7494 334294
rect 6874 334170 6970 334226
rect 7026 334170 7094 334226
rect 7150 334170 7218 334226
rect 7274 334170 7342 334226
rect 7398 334170 7494 334226
rect 6874 334102 7494 334170
rect 6874 334046 6970 334102
rect 7026 334046 7094 334102
rect 7150 334046 7218 334102
rect 7274 334046 7342 334102
rect 7398 334046 7494 334102
rect 6874 333978 7494 334046
rect 6874 333922 6970 333978
rect 7026 333922 7094 333978
rect 7150 333922 7218 333978
rect 7274 333922 7342 333978
rect 7398 333922 7494 333978
rect 6874 316350 7494 333922
rect 6874 316294 6970 316350
rect 7026 316294 7094 316350
rect 7150 316294 7218 316350
rect 7274 316294 7342 316350
rect 7398 316294 7494 316350
rect 6874 316226 7494 316294
rect 6874 316170 6970 316226
rect 7026 316170 7094 316226
rect 7150 316170 7218 316226
rect 7274 316170 7342 316226
rect 7398 316170 7494 316226
rect 6874 316102 7494 316170
rect 6874 316046 6970 316102
rect 7026 316046 7094 316102
rect 7150 316046 7218 316102
rect 7274 316046 7342 316102
rect 7398 316046 7494 316102
rect 6874 315978 7494 316046
rect 6874 315922 6970 315978
rect 7026 315922 7094 315978
rect 7150 315922 7218 315978
rect 7274 315922 7342 315978
rect 7398 315922 7494 315978
rect 6874 298350 7494 315922
rect 6874 298294 6970 298350
rect 7026 298294 7094 298350
rect 7150 298294 7218 298350
rect 7274 298294 7342 298350
rect 7398 298294 7494 298350
rect 6874 298226 7494 298294
rect 6874 298170 6970 298226
rect 7026 298170 7094 298226
rect 7150 298170 7218 298226
rect 7274 298170 7342 298226
rect 7398 298170 7494 298226
rect 6874 298102 7494 298170
rect 6874 298046 6970 298102
rect 7026 298046 7094 298102
rect 7150 298046 7218 298102
rect 7274 298046 7342 298102
rect 7398 298046 7494 298102
rect 6874 297978 7494 298046
rect 6874 297922 6970 297978
rect 7026 297922 7094 297978
rect 7150 297922 7218 297978
rect 7274 297922 7342 297978
rect 7398 297922 7494 297978
rect 6874 280350 7494 297922
rect 6874 280294 6970 280350
rect 7026 280294 7094 280350
rect 7150 280294 7218 280350
rect 7274 280294 7342 280350
rect 7398 280294 7494 280350
rect 6874 280226 7494 280294
rect 6874 280170 6970 280226
rect 7026 280170 7094 280226
rect 7150 280170 7218 280226
rect 7274 280170 7342 280226
rect 7398 280170 7494 280226
rect 6874 280102 7494 280170
rect 6874 280046 6970 280102
rect 7026 280046 7094 280102
rect 7150 280046 7218 280102
rect 7274 280046 7342 280102
rect 7398 280046 7494 280102
rect 6874 279978 7494 280046
rect 6874 279922 6970 279978
rect 7026 279922 7094 279978
rect 7150 279922 7218 279978
rect 7274 279922 7342 279978
rect 7398 279922 7494 279978
rect 6874 262350 7494 279922
rect 6874 262294 6970 262350
rect 7026 262294 7094 262350
rect 7150 262294 7218 262350
rect 7274 262294 7342 262350
rect 7398 262294 7494 262350
rect 6874 262226 7494 262294
rect 6874 262170 6970 262226
rect 7026 262170 7094 262226
rect 7150 262170 7218 262226
rect 7274 262170 7342 262226
rect 7398 262170 7494 262226
rect 6874 262102 7494 262170
rect 6874 262046 6970 262102
rect 7026 262046 7094 262102
rect 7150 262046 7218 262102
rect 7274 262046 7342 262102
rect 7398 262046 7494 262102
rect 6874 261978 7494 262046
rect 6874 261922 6970 261978
rect 7026 261922 7094 261978
rect 7150 261922 7218 261978
rect 7274 261922 7342 261978
rect 7398 261922 7494 261978
rect 6874 244350 7494 261922
rect 6874 244294 6970 244350
rect 7026 244294 7094 244350
rect 7150 244294 7218 244350
rect 7274 244294 7342 244350
rect 7398 244294 7494 244350
rect 6874 244226 7494 244294
rect 6874 244170 6970 244226
rect 7026 244170 7094 244226
rect 7150 244170 7218 244226
rect 7274 244170 7342 244226
rect 7398 244170 7494 244226
rect 6874 244102 7494 244170
rect 6874 244046 6970 244102
rect 7026 244046 7094 244102
rect 7150 244046 7218 244102
rect 7274 244046 7342 244102
rect 7398 244046 7494 244102
rect 6874 243978 7494 244046
rect 6874 243922 6970 243978
rect 7026 243922 7094 243978
rect 7150 243922 7218 243978
rect 7274 243922 7342 243978
rect 7398 243922 7494 243978
rect 6874 226350 7494 243922
rect 6874 226294 6970 226350
rect 7026 226294 7094 226350
rect 7150 226294 7218 226350
rect 7274 226294 7342 226350
rect 7398 226294 7494 226350
rect 6874 226226 7494 226294
rect 6874 226170 6970 226226
rect 7026 226170 7094 226226
rect 7150 226170 7218 226226
rect 7274 226170 7342 226226
rect 7398 226170 7494 226226
rect 6874 226102 7494 226170
rect 6874 226046 6970 226102
rect 7026 226046 7094 226102
rect 7150 226046 7218 226102
rect 7274 226046 7342 226102
rect 7398 226046 7494 226102
rect 6874 225978 7494 226046
rect 6874 225922 6970 225978
rect 7026 225922 7094 225978
rect 7150 225922 7218 225978
rect 7274 225922 7342 225978
rect 7398 225922 7494 225978
rect 6874 208350 7494 225922
rect 6874 208294 6970 208350
rect 7026 208294 7094 208350
rect 7150 208294 7218 208350
rect 7274 208294 7342 208350
rect 7398 208294 7494 208350
rect 6874 208226 7494 208294
rect 6874 208170 6970 208226
rect 7026 208170 7094 208226
rect 7150 208170 7218 208226
rect 7274 208170 7342 208226
rect 7398 208170 7494 208226
rect 6874 208102 7494 208170
rect 6874 208046 6970 208102
rect 7026 208046 7094 208102
rect 7150 208046 7218 208102
rect 7274 208046 7342 208102
rect 7398 208046 7494 208102
rect 6874 207978 7494 208046
rect 6874 207922 6970 207978
rect 7026 207922 7094 207978
rect 7150 207922 7218 207978
rect 7274 207922 7342 207978
rect 7398 207922 7494 207978
rect 6874 190350 7494 207922
rect 6874 190294 6970 190350
rect 7026 190294 7094 190350
rect 7150 190294 7218 190350
rect 7274 190294 7342 190350
rect 7398 190294 7494 190350
rect 6874 190226 7494 190294
rect 6874 190170 6970 190226
rect 7026 190170 7094 190226
rect 7150 190170 7218 190226
rect 7274 190170 7342 190226
rect 7398 190170 7494 190226
rect 6874 190102 7494 190170
rect 6874 190046 6970 190102
rect 7026 190046 7094 190102
rect 7150 190046 7218 190102
rect 7274 190046 7342 190102
rect 7398 190046 7494 190102
rect 6874 189978 7494 190046
rect 6874 189922 6970 189978
rect 7026 189922 7094 189978
rect 7150 189922 7218 189978
rect 7274 189922 7342 189978
rect 7398 189922 7494 189978
rect 6874 172350 7494 189922
rect 6874 172294 6970 172350
rect 7026 172294 7094 172350
rect 7150 172294 7218 172350
rect 7274 172294 7342 172350
rect 7398 172294 7494 172350
rect 6874 172226 7494 172294
rect 6874 172170 6970 172226
rect 7026 172170 7094 172226
rect 7150 172170 7218 172226
rect 7274 172170 7342 172226
rect 7398 172170 7494 172226
rect 6874 172102 7494 172170
rect 6874 172046 6970 172102
rect 7026 172046 7094 172102
rect 7150 172046 7218 172102
rect 7274 172046 7342 172102
rect 7398 172046 7494 172102
rect 6874 171978 7494 172046
rect 6874 171922 6970 171978
rect 7026 171922 7094 171978
rect 7150 171922 7218 171978
rect 7274 171922 7342 171978
rect 7398 171922 7494 171978
rect 6874 154350 7494 171922
rect 6874 154294 6970 154350
rect 7026 154294 7094 154350
rect 7150 154294 7218 154350
rect 7274 154294 7342 154350
rect 7398 154294 7494 154350
rect 6874 154226 7494 154294
rect 6874 154170 6970 154226
rect 7026 154170 7094 154226
rect 7150 154170 7218 154226
rect 7274 154170 7342 154226
rect 7398 154170 7494 154226
rect 6874 154102 7494 154170
rect 6874 154046 6970 154102
rect 7026 154046 7094 154102
rect 7150 154046 7218 154102
rect 7274 154046 7342 154102
rect 7398 154046 7494 154102
rect 6874 153978 7494 154046
rect 6874 153922 6970 153978
rect 7026 153922 7094 153978
rect 7150 153922 7218 153978
rect 7274 153922 7342 153978
rect 7398 153922 7494 153978
rect 6874 136350 7494 153922
rect 6874 136294 6970 136350
rect 7026 136294 7094 136350
rect 7150 136294 7218 136350
rect 7274 136294 7342 136350
rect 7398 136294 7494 136350
rect 6874 136226 7494 136294
rect 6874 136170 6970 136226
rect 7026 136170 7094 136226
rect 7150 136170 7218 136226
rect 7274 136170 7342 136226
rect 7398 136170 7494 136226
rect 6874 136102 7494 136170
rect 6874 136046 6970 136102
rect 7026 136046 7094 136102
rect 7150 136046 7218 136102
rect 7274 136046 7342 136102
rect 7398 136046 7494 136102
rect 6874 135978 7494 136046
rect 6874 135922 6970 135978
rect 7026 135922 7094 135978
rect 7150 135922 7218 135978
rect 7274 135922 7342 135978
rect 7398 135922 7494 135978
rect 6874 118350 7494 135922
rect 6874 118294 6970 118350
rect 7026 118294 7094 118350
rect 7150 118294 7218 118350
rect 7274 118294 7342 118350
rect 7398 118294 7494 118350
rect 6874 118226 7494 118294
rect 6874 118170 6970 118226
rect 7026 118170 7094 118226
rect 7150 118170 7218 118226
rect 7274 118170 7342 118226
rect 7398 118170 7494 118226
rect 6874 118102 7494 118170
rect 6874 118046 6970 118102
rect 7026 118046 7094 118102
rect 7150 118046 7218 118102
rect 7274 118046 7342 118102
rect 7398 118046 7494 118102
rect 6874 117978 7494 118046
rect 6874 117922 6970 117978
rect 7026 117922 7094 117978
rect 7150 117922 7218 117978
rect 7274 117922 7342 117978
rect 7398 117922 7494 117978
rect 6874 100350 7494 117922
rect 6874 100294 6970 100350
rect 7026 100294 7094 100350
rect 7150 100294 7218 100350
rect 7274 100294 7342 100350
rect 7398 100294 7494 100350
rect 6874 100226 7494 100294
rect 6874 100170 6970 100226
rect 7026 100170 7094 100226
rect 7150 100170 7218 100226
rect 7274 100170 7342 100226
rect 7398 100170 7494 100226
rect 6874 100102 7494 100170
rect 6874 100046 6970 100102
rect 7026 100046 7094 100102
rect 7150 100046 7218 100102
rect 7274 100046 7342 100102
rect 7398 100046 7494 100102
rect 6874 99978 7494 100046
rect 6874 99922 6970 99978
rect 7026 99922 7094 99978
rect 7150 99922 7218 99978
rect 7274 99922 7342 99978
rect 7398 99922 7494 99978
rect 6874 82350 7494 99922
rect 6874 82294 6970 82350
rect 7026 82294 7094 82350
rect 7150 82294 7218 82350
rect 7274 82294 7342 82350
rect 7398 82294 7494 82350
rect 6874 82226 7494 82294
rect 6874 82170 6970 82226
rect 7026 82170 7094 82226
rect 7150 82170 7218 82226
rect 7274 82170 7342 82226
rect 7398 82170 7494 82226
rect 6874 82102 7494 82170
rect 6874 82046 6970 82102
rect 7026 82046 7094 82102
rect 7150 82046 7218 82102
rect 7274 82046 7342 82102
rect 7398 82046 7494 82102
rect 6874 81978 7494 82046
rect 6874 81922 6970 81978
rect 7026 81922 7094 81978
rect 7150 81922 7218 81978
rect 7274 81922 7342 81978
rect 7398 81922 7494 81978
rect 6874 64350 7494 81922
rect 6874 64294 6970 64350
rect 7026 64294 7094 64350
rect 7150 64294 7218 64350
rect 7274 64294 7342 64350
rect 7398 64294 7494 64350
rect 6874 64226 7494 64294
rect 6874 64170 6970 64226
rect 7026 64170 7094 64226
rect 7150 64170 7218 64226
rect 7274 64170 7342 64226
rect 7398 64170 7494 64226
rect 6874 64102 7494 64170
rect 6874 64046 6970 64102
rect 7026 64046 7094 64102
rect 7150 64046 7218 64102
rect 7274 64046 7342 64102
rect 7398 64046 7494 64102
rect 6874 63978 7494 64046
rect 6874 63922 6970 63978
rect 7026 63922 7094 63978
rect 7150 63922 7218 63978
rect 7274 63922 7342 63978
rect 7398 63922 7494 63978
rect 6874 46350 7494 63922
rect 6874 46294 6970 46350
rect 7026 46294 7094 46350
rect 7150 46294 7218 46350
rect 7274 46294 7342 46350
rect 7398 46294 7494 46350
rect 6874 46226 7494 46294
rect 6874 46170 6970 46226
rect 7026 46170 7094 46226
rect 7150 46170 7218 46226
rect 7274 46170 7342 46226
rect 7398 46170 7494 46226
rect 6874 46102 7494 46170
rect 6874 46046 6970 46102
rect 7026 46046 7094 46102
rect 7150 46046 7218 46102
rect 7274 46046 7342 46102
rect 7398 46046 7494 46102
rect 6874 45978 7494 46046
rect 6874 45922 6970 45978
rect 7026 45922 7094 45978
rect 7150 45922 7218 45978
rect 7274 45922 7342 45978
rect 7398 45922 7494 45978
rect 6874 28350 7494 45922
rect 6874 28294 6970 28350
rect 7026 28294 7094 28350
rect 7150 28294 7218 28350
rect 7274 28294 7342 28350
rect 7398 28294 7494 28350
rect 6874 28226 7494 28294
rect 6874 28170 6970 28226
rect 7026 28170 7094 28226
rect 7150 28170 7218 28226
rect 7274 28170 7342 28226
rect 7398 28170 7494 28226
rect 6874 28102 7494 28170
rect 6874 28046 6970 28102
rect 7026 28046 7094 28102
rect 7150 28046 7218 28102
rect 7274 28046 7342 28102
rect 7398 28046 7494 28102
rect 6874 27978 7494 28046
rect 6874 27922 6970 27978
rect 7026 27922 7094 27978
rect 7150 27922 7218 27978
rect 7274 27922 7342 27978
rect 7398 27922 7494 27978
rect 6874 10350 7494 27922
rect 7644 551236 7700 551246
rect 7644 16772 7700 551180
rect 9884 316820 9940 316830
rect 9772 313460 9828 313470
rect 9660 303380 9716 303390
rect 9660 150388 9716 303324
rect 9772 154532 9828 313404
rect 9772 154466 9828 154476
rect 9660 150322 9716 150332
rect 9884 147028 9940 316764
rect 9884 146962 9940 146972
rect 9996 18452 10052 587916
rect 21154 580350 21774 596784
rect 21154 580294 21250 580350
rect 21306 580294 21374 580350
rect 21430 580294 21498 580350
rect 21554 580294 21622 580350
rect 21678 580294 21774 580350
rect 21154 580226 21774 580294
rect 21154 580170 21250 580226
rect 21306 580170 21374 580226
rect 21430 580170 21498 580226
rect 21554 580170 21622 580226
rect 21678 580170 21774 580226
rect 21154 580102 21774 580170
rect 21154 580046 21250 580102
rect 21306 580046 21374 580102
rect 21430 580046 21498 580102
rect 21554 580046 21622 580102
rect 21678 580046 21774 580102
rect 21154 579978 21774 580046
rect 21154 579922 21250 579978
rect 21306 579922 21374 579978
rect 21430 579922 21498 579978
rect 21554 579922 21622 579978
rect 21678 579922 21774 579978
rect 21154 562350 21774 579922
rect 21154 562294 21250 562350
rect 21306 562294 21374 562350
rect 21430 562294 21498 562350
rect 21554 562294 21622 562350
rect 21678 562294 21774 562350
rect 21154 562226 21774 562294
rect 21154 562170 21250 562226
rect 21306 562170 21374 562226
rect 21430 562170 21498 562226
rect 21554 562170 21622 562226
rect 21678 562170 21774 562226
rect 21154 562102 21774 562170
rect 21154 562046 21250 562102
rect 21306 562046 21374 562102
rect 21430 562046 21498 562102
rect 21554 562046 21622 562102
rect 21678 562046 21774 562102
rect 21154 561978 21774 562046
rect 21154 561922 21250 561978
rect 21306 561922 21374 561978
rect 21430 561922 21498 561978
rect 21554 561922 21622 561978
rect 21678 561922 21774 561978
rect 21154 544350 21774 561922
rect 21154 544294 21250 544350
rect 21306 544294 21374 544350
rect 21430 544294 21498 544350
rect 21554 544294 21622 544350
rect 21678 544294 21774 544350
rect 21154 544226 21774 544294
rect 21154 544170 21250 544226
rect 21306 544170 21374 544226
rect 21430 544170 21498 544226
rect 21554 544170 21622 544226
rect 21678 544170 21774 544226
rect 21154 544102 21774 544170
rect 21154 544046 21250 544102
rect 21306 544046 21374 544102
rect 21430 544046 21498 544102
rect 21554 544046 21622 544102
rect 21678 544046 21774 544102
rect 21154 543978 21774 544046
rect 21154 543922 21250 543978
rect 21306 543922 21374 543978
rect 21430 543922 21498 543978
rect 21554 543922 21622 543978
rect 21678 543922 21774 543978
rect 21154 526350 21774 543922
rect 21154 526294 21250 526350
rect 21306 526294 21374 526350
rect 21430 526294 21498 526350
rect 21554 526294 21622 526350
rect 21678 526294 21774 526350
rect 21154 526226 21774 526294
rect 21154 526170 21250 526226
rect 21306 526170 21374 526226
rect 21430 526170 21498 526226
rect 21554 526170 21622 526226
rect 21678 526170 21774 526226
rect 21154 526102 21774 526170
rect 21154 526046 21250 526102
rect 21306 526046 21374 526102
rect 21430 526046 21498 526102
rect 21554 526046 21622 526102
rect 21678 526046 21774 526102
rect 21154 525978 21774 526046
rect 21154 525922 21250 525978
rect 21306 525922 21374 525978
rect 21430 525922 21498 525978
rect 21554 525922 21622 525978
rect 21678 525922 21774 525978
rect 21154 508350 21774 525922
rect 21154 508294 21250 508350
rect 21306 508294 21374 508350
rect 21430 508294 21498 508350
rect 21554 508294 21622 508350
rect 21678 508294 21774 508350
rect 21154 508226 21774 508294
rect 21154 508170 21250 508226
rect 21306 508170 21374 508226
rect 21430 508170 21498 508226
rect 21554 508170 21622 508226
rect 21678 508170 21774 508226
rect 21154 508102 21774 508170
rect 21154 508046 21250 508102
rect 21306 508046 21374 508102
rect 21430 508046 21498 508102
rect 21554 508046 21622 508102
rect 21678 508046 21774 508102
rect 21154 507978 21774 508046
rect 21154 507922 21250 507978
rect 21306 507922 21374 507978
rect 21430 507922 21498 507978
rect 21554 507922 21622 507978
rect 21678 507922 21774 507978
rect 21154 490350 21774 507922
rect 21154 490294 21250 490350
rect 21306 490294 21374 490350
rect 21430 490294 21498 490350
rect 21554 490294 21622 490350
rect 21678 490294 21774 490350
rect 21154 490226 21774 490294
rect 21154 490170 21250 490226
rect 21306 490170 21374 490226
rect 21430 490170 21498 490226
rect 21554 490170 21622 490226
rect 21678 490170 21774 490226
rect 21154 490102 21774 490170
rect 21154 490046 21250 490102
rect 21306 490046 21374 490102
rect 21430 490046 21498 490102
rect 21554 490046 21622 490102
rect 21678 490046 21774 490102
rect 21154 489978 21774 490046
rect 21154 489922 21250 489978
rect 21306 489922 21374 489978
rect 21430 489922 21498 489978
rect 21554 489922 21622 489978
rect 21678 489922 21774 489978
rect 21154 472350 21774 489922
rect 21154 472294 21250 472350
rect 21306 472294 21374 472350
rect 21430 472294 21498 472350
rect 21554 472294 21622 472350
rect 21678 472294 21774 472350
rect 21154 472226 21774 472294
rect 21154 472170 21250 472226
rect 21306 472170 21374 472226
rect 21430 472170 21498 472226
rect 21554 472170 21622 472226
rect 21678 472170 21774 472226
rect 21154 472102 21774 472170
rect 21154 472046 21250 472102
rect 21306 472046 21374 472102
rect 21430 472046 21498 472102
rect 21554 472046 21622 472102
rect 21678 472046 21774 472102
rect 21154 471978 21774 472046
rect 21154 471922 21250 471978
rect 21306 471922 21374 471978
rect 21430 471922 21498 471978
rect 21554 471922 21622 471978
rect 21678 471922 21774 471978
rect 21154 458342 21774 471922
rect 24874 598172 25494 598268
rect 24874 598116 24970 598172
rect 25026 598116 25094 598172
rect 25150 598116 25218 598172
rect 25274 598116 25342 598172
rect 25398 598116 25494 598172
rect 24874 598048 25494 598116
rect 24874 597992 24970 598048
rect 25026 597992 25094 598048
rect 25150 597992 25218 598048
rect 25274 597992 25342 598048
rect 25398 597992 25494 598048
rect 24874 597924 25494 597992
rect 24874 597868 24970 597924
rect 25026 597868 25094 597924
rect 25150 597868 25218 597924
rect 25274 597868 25342 597924
rect 25398 597868 25494 597924
rect 24874 597800 25494 597868
rect 24874 597744 24970 597800
rect 25026 597744 25094 597800
rect 25150 597744 25218 597800
rect 25274 597744 25342 597800
rect 25398 597744 25494 597800
rect 24874 586350 25494 597744
rect 24874 586294 24970 586350
rect 25026 586294 25094 586350
rect 25150 586294 25218 586350
rect 25274 586294 25342 586350
rect 25398 586294 25494 586350
rect 24874 586226 25494 586294
rect 24874 586170 24970 586226
rect 25026 586170 25094 586226
rect 25150 586170 25218 586226
rect 25274 586170 25342 586226
rect 25398 586170 25494 586226
rect 24874 586102 25494 586170
rect 24874 586046 24970 586102
rect 25026 586046 25094 586102
rect 25150 586046 25218 586102
rect 25274 586046 25342 586102
rect 25398 586046 25494 586102
rect 24874 585978 25494 586046
rect 24874 585922 24970 585978
rect 25026 585922 25094 585978
rect 25150 585922 25218 585978
rect 25274 585922 25342 585978
rect 25398 585922 25494 585978
rect 24874 568350 25494 585922
rect 24874 568294 24970 568350
rect 25026 568294 25094 568350
rect 25150 568294 25218 568350
rect 25274 568294 25342 568350
rect 25398 568294 25494 568350
rect 24874 568226 25494 568294
rect 24874 568170 24970 568226
rect 25026 568170 25094 568226
rect 25150 568170 25218 568226
rect 25274 568170 25342 568226
rect 25398 568170 25494 568226
rect 24874 568102 25494 568170
rect 24874 568046 24970 568102
rect 25026 568046 25094 568102
rect 25150 568046 25218 568102
rect 25274 568046 25342 568102
rect 25398 568046 25494 568102
rect 24874 567978 25494 568046
rect 24874 567922 24970 567978
rect 25026 567922 25094 567978
rect 25150 567922 25218 567978
rect 25274 567922 25342 567978
rect 25398 567922 25494 567978
rect 24874 550350 25494 567922
rect 24874 550294 24970 550350
rect 25026 550294 25094 550350
rect 25150 550294 25218 550350
rect 25274 550294 25342 550350
rect 25398 550294 25494 550350
rect 24874 550226 25494 550294
rect 24874 550170 24970 550226
rect 25026 550170 25094 550226
rect 25150 550170 25218 550226
rect 25274 550170 25342 550226
rect 25398 550170 25494 550226
rect 24874 550102 25494 550170
rect 24874 550046 24970 550102
rect 25026 550046 25094 550102
rect 25150 550046 25218 550102
rect 25274 550046 25342 550102
rect 25398 550046 25494 550102
rect 24874 549978 25494 550046
rect 24874 549922 24970 549978
rect 25026 549922 25094 549978
rect 25150 549922 25218 549978
rect 25274 549922 25342 549978
rect 25398 549922 25494 549978
rect 24874 532350 25494 549922
rect 24874 532294 24970 532350
rect 25026 532294 25094 532350
rect 25150 532294 25218 532350
rect 25274 532294 25342 532350
rect 25398 532294 25494 532350
rect 24874 532226 25494 532294
rect 24874 532170 24970 532226
rect 25026 532170 25094 532226
rect 25150 532170 25218 532226
rect 25274 532170 25342 532226
rect 25398 532170 25494 532226
rect 24874 532102 25494 532170
rect 24874 532046 24970 532102
rect 25026 532046 25094 532102
rect 25150 532046 25218 532102
rect 25274 532046 25342 532102
rect 25398 532046 25494 532102
rect 24874 531978 25494 532046
rect 24874 531922 24970 531978
rect 25026 531922 25094 531978
rect 25150 531922 25218 531978
rect 25274 531922 25342 531978
rect 25398 531922 25494 531978
rect 24874 514350 25494 531922
rect 24874 514294 24970 514350
rect 25026 514294 25094 514350
rect 25150 514294 25218 514350
rect 25274 514294 25342 514350
rect 25398 514294 25494 514350
rect 24874 514226 25494 514294
rect 24874 514170 24970 514226
rect 25026 514170 25094 514226
rect 25150 514170 25218 514226
rect 25274 514170 25342 514226
rect 25398 514170 25494 514226
rect 24874 514102 25494 514170
rect 24874 514046 24970 514102
rect 25026 514046 25094 514102
rect 25150 514046 25218 514102
rect 25274 514046 25342 514102
rect 25398 514046 25494 514102
rect 24874 513978 25494 514046
rect 24874 513922 24970 513978
rect 25026 513922 25094 513978
rect 25150 513922 25218 513978
rect 25274 513922 25342 513978
rect 25398 513922 25494 513978
rect 24874 496350 25494 513922
rect 24874 496294 24970 496350
rect 25026 496294 25094 496350
rect 25150 496294 25218 496350
rect 25274 496294 25342 496350
rect 25398 496294 25494 496350
rect 24874 496226 25494 496294
rect 24874 496170 24970 496226
rect 25026 496170 25094 496226
rect 25150 496170 25218 496226
rect 25274 496170 25342 496226
rect 25398 496170 25494 496226
rect 24874 496102 25494 496170
rect 24874 496046 24970 496102
rect 25026 496046 25094 496102
rect 25150 496046 25218 496102
rect 25274 496046 25342 496102
rect 25398 496046 25494 496102
rect 24874 495978 25494 496046
rect 24874 495922 24970 495978
rect 25026 495922 25094 495978
rect 25150 495922 25218 495978
rect 25274 495922 25342 495978
rect 25398 495922 25494 495978
rect 24874 478350 25494 495922
rect 24874 478294 24970 478350
rect 25026 478294 25094 478350
rect 25150 478294 25218 478350
rect 25274 478294 25342 478350
rect 25398 478294 25494 478350
rect 24874 478226 25494 478294
rect 24874 478170 24970 478226
rect 25026 478170 25094 478226
rect 25150 478170 25218 478226
rect 25274 478170 25342 478226
rect 25398 478170 25494 478226
rect 24874 478102 25494 478170
rect 24874 478046 24970 478102
rect 25026 478046 25094 478102
rect 25150 478046 25218 478102
rect 25274 478046 25342 478102
rect 25398 478046 25494 478102
rect 24874 477978 25494 478046
rect 24874 477922 24970 477978
rect 25026 477922 25094 477978
rect 25150 477922 25218 477978
rect 25274 477922 25342 477978
rect 25398 477922 25494 477978
rect 24874 460350 25494 477922
rect 24874 460294 24970 460350
rect 25026 460294 25094 460350
rect 25150 460294 25218 460350
rect 25274 460294 25342 460350
rect 25398 460294 25494 460350
rect 24874 460226 25494 460294
rect 24874 460170 24970 460226
rect 25026 460170 25094 460226
rect 25150 460170 25218 460226
rect 25274 460170 25342 460226
rect 25398 460170 25494 460226
rect 24874 460102 25494 460170
rect 24874 460046 24970 460102
rect 25026 460046 25094 460102
rect 25150 460046 25218 460102
rect 25274 460046 25342 460102
rect 25398 460046 25494 460102
rect 24874 459978 25494 460046
rect 24874 459922 24970 459978
rect 25026 459922 25094 459978
rect 25150 459922 25218 459978
rect 25274 459922 25342 459978
rect 25398 459922 25494 459978
rect 24874 458342 25494 459922
rect 39154 597212 39774 598268
rect 39154 597156 39250 597212
rect 39306 597156 39374 597212
rect 39430 597156 39498 597212
rect 39554 597156 39622 597212
rect 39678 597156 39774 597212
rect 39154 597088 39774 597156
rect 39154 597032 39250 597088
rect 39306 597032 39374 597088
rect 39430 597032 39498 597088
rect 39554 597032 39622 597088
rect 39678 597032 39774 597088
rect 39154 596964 39774 597032
rect 39154 596908 39250 596964
rect 39306 596908 39374 596964
rect 39430 596908 39498 596964
rect 39554 596908 39622 596964
rect 39678 596908 39774 596964
rect 39154 596840 39774 596908
rect 39154 596784 39250 596840
rect 39306 596784 39374 596840
rect 39430 596784 39498 596840
rect 39554 596784 39622 596840
rect 39678 596784 39774 596840
rect 39154 580350 39774 596784
rect 39154 580294 39250 580350
rect 39306 580294 39374 580350
rect 39430 580294 39498 580350
rect 39554 580294 39622 580350
rect 39678 580294 39774 580350
rect 39154 580226 39774 580294
rect 39154 580170 39250 580226
rect 39306 580170 39374 580226
rect 39430 580170 39498 580226
rect 39554 580170 39622 580226
rect 39678 580170 39774 580226
rect 39154 580102 39774 580170
rect 39154 580046 39250 580102
rect 39306 580046 39374 580102
rect 39430 580046 39498 580102
rect 39554 580046 39622 580102
rect 39678 580046 39774 580102
rect 39154 579978 39774 580046
rect 39154 579922 39250 579978
rect 39306 579922 39374 579978
rect 39430 579922 39498 579978
rect 39554 579922 39622 579978
rect 39678 579922 39774 579978
rect 39154 562350 39774 579922
rect 39154 562294 39250 562350
rect 39306 562294 39374 562350
rect 39430 562294 39498 562350
rect 39554 562294 39622 562350
rect 39678 562294 39774 562350
rect 39154 562226 39774 562294
rect 39154 562170 39250 562226
rect 39306 562170 39374 562226
rect 39430 562170 39498 562226
rect 39554 562170 39622 562226
rect 39678 562170 39774 562226
rect 39154 562102 39774 562170
rect 39154 562046 39250 562102
rect 39306 562046 39374 562102
rect 39430 562046 39498 562102
rect 39554 562046 39622 562102
rect 39678 562046 39774 562102
rect 39154 561978 39774 562046
rect 39154 561922 39250 561978
rect 39306 561922 39374 561978
rect 39430 561922 39498 561978
rect 39554 561922 39622 561978
rect 39678 561922 39774 561978
rect 39154 544350 39774 561922
rect 39154 544294 39250 544350
rect 39306 544294 39374 544350
rect 39430 544294 39498 544350
rect 39554 544294 39622 544350
rect 39678 544294 39774 544350
rect 39154 544226 39774 544294
rect 39154 544170 39250 544226
rect 39306 544170 39374 544226
rect 39430 544170 39498 544226
rect 39554 544170 39622 544226
rect 39678 544170 39774 544226
rect 39154 544102 39774 544170
rect 39154 544046 39250 544102
rect 39306 544046 39374 544102
rect 39430 544046 39498 544102
rect 39554 544046 39622 544102
rect 39678 544046 39774 544102
rect 39154 543978 39774 544046
rect 39154 543922 39250 543978
rect 39306 543922 39374 543978
rect 39430 543922 39498 543978
rect 39554 543922 39622 543978
rect 39678 543922 39774 543978
rect 39154 526350 39774 543922
rect 39154 526294 39250 526350
rect 39306 526294 39374 526350
rect 39430 526294 39498 526350
rect 39554 526294 39622 526350
rect 39678 526294 39774 526350
rect 39154 526226 39774 526294
rect 39154 526170 39250 526226
rect 39306 526170 39374 526226
rect 39430 526170 39498 526226
rect 39554 526170 39622 526226
rect 39678 526170 39774 526226
rect 39154 526102 39774 526170
rect 39154 526046 39250 526102
rect 39306 526046 39374 526102
rect 39430 526046 39498 526102
rect 39554 526046 39622 526102
rect 39678 526046 39774 526102
rect 39154 525978 39774 526046
rect 39154 525922 39250 525978
rect 39306 525922 39374 525978
rect 39430 525922 39498 525978
rect 39554 525922 39622 525978
rect 39678 525922 39774 525978
rect 39154 508350 39774 525922
rect 39154 508294 39250 508350
rect 39306 508294 39374 508350
rect 39430 508294 39498 508350
rect 39554 508294 39622 508350
rect 39678 508294 39774 508350
rect 39154 508226 39774 508294
rect 39154 508170 39250 508226
rect 39306 508170 39374 508226
rect 39430 508170 39498 508226
rect 39554 508170 39622 508226
rect 39678 508170 39774 508226
rect 39154 508102 39774 508170
rect 39154 508046 39250 508102
rect 39306 508046 39374 508102
rect 39430 508046 39498 508102
rect 39554 508046 39622 508102
rect 39678 508046 39774 508102
rect 39154 507978 39774 508046
rect 39154 507922 39250 507978
rect 39306 507922 39374 507978
rect 39430 507922 39498 507978
rect 39554 507922 39622 507978
rect 39678 507922 39774 507978
rect 39154 490350 39774 507922
rect 39154 490294 39250 490350
rect 39306 490294 39374 490350
rect 39430 490294 39498 490350
rect 39554 490294 39622 490350
rect 39678 490294 39774 490350
rect 39154 490226 39774 490294
rect 39154 490170 39250 490226
rect 39306 490170 39374 490226
rect 39430 490170 39498 490226
rect 39554 490170 39622 490226
rect 39678 490170 39774 490226
rect 39154 490102 39774 490170
rect 39154 490046 39250 490102
rect 39306 490046 39374 490102
rect 39430 490046 39498 490102
rect 39554 490046 39622 490102
rect 39678 490046 39774 490102
rect 39154 489978 39774 490046
rect 39154 489922 39250 489978
rect 39306 489922 39374 489978
rect 39430 489922 39498 489978
rect 39554 489922 39622 489978
rect 39678 489922 39774 489978
rect 39154 472350 39774 489922
rect 39154 472294 39250 472350
rect 39306 472294 39374 472350
rect 39430 472294 39498 472350
rect 39554 472294 39622 472350
rect 39678 472294 39774 472350
rect 39154 472226 39774 472294
rect 39154 472170 39250 472226
rect 39306 472170 39374 472226
rect 39430 472170 39498 472226
rect 39554 472170 39622 472226
rect 39678 472170 39774 472226
rect 39154 472102 39774 472170
rect 39154 472046 39250 472102
rect 39306 472046 39374 472102
rect 39430 472046 39498 472102
rect 39554 472046 39622 472102
rect 39678 472046 39774 472102
rect 39154 471978 39774 472046
rect 39154 471922 39250 471978
rect 39306 471922 39374 471978
rect 39430 471922 39498 471978
rect 39554 471922 39622 471978
rect 39678 471922 39774 471978
rect 39154 458342 39774 471922
rect 42874 598172 43494 598268
rect 42874 598116 42970 598172
rect 43026 598116 43094 598172
rect 43150 598116 43218 598172
rect 43274 598116 43342 598172
rect 43398 598116 43494 598172
rect 42874 598048 43494 598116
rect 42874 597992 42970 598048
rect 43026 597992 43094 598048
rect 43150 597992 43218 598048
rect 43274 597992 43342 598048
rect 43398 597992 43494 598048
rect 42874 597924 43494 597992
rect 42874 597868 42970 597924
rect 43026 597868 43094 597924
rect 43150 597868 43218 597924
rect 43274 597868 43342 597924
rect 43398 597868 43494 597924
rect 42874 597800 43494 597868
rect 42874 597744 42970 597800
rect 43026 597744 43094 597800
rect 43150 597744 43218 597800
rect 43274 597744 43342 597800
rect 43398 597744 43494 597800
rect 42874 586350 43494 597744
rect 42874 586294 42970 586350
rect 43026 586294 43094 586350
rect 43150 586294 43218 586350
rect 43274 586294 43342 586350
rect 43398 586294 43494 586350
rect 42874 586226 43494 586294
rect 42874 586170 42970 586226
rect 43026 586170 43094 586226
rect 43150 586170 43218 586226
rect 43274 586170 43342 586226
rect 43398 586170 43494 586226
rect 42874 586102 43494 586170
rect 42874 586046 42970 586102
rect 43026 586046 43094 586102
rect 43150 586046 43218 586102
rect 43274 586046 43342 586102
rect 43398 586046 43494 586102
rect 42874 585978 43494 586046
rect 42874 585922 42970 585978
rect 43026 585922 43094 585978
rect 43150 585922 43218 585978
rect 43274 585922 43342 585978
rect 43398 585922 43494 585978
rect 42874 568350 43494 585922
rect 42874 568294 42970 568350
rect 43026 568294 43094 568350
rect 43150 568294 43218 568350
rect 43274 568294 43342 568350
rect 43398 568294 43494 568350
rect 42874 568226 43494 568294
rect 42874 568170 42970 568226
rect 43026 568170 43094 568226
rect 43150 568170 43218 568226
rect 43274 568170 43342 568226
rect 43398 568170 43494 568226
rect 42874 568102 43494 568170
rect 42874 568046 42970 568102
rect 43026 568046 43094 568102
rect 43150 568046 43218 568102
rect 43274 568046 43342 568102
rect 43398 568046 43494 568102
rect 42874 567978 43494 568046
rect 42874 567922 42970 567978
rect 43026 567922 43094 567978
rect 43150 567922 43218 567978
rect 43274 567922 43342 567978
rect 43398 567922 43494 567978
rect 42874 550350 43494 567922
rect 42874 550294 42970 550350
rect 43026 550294 43094 550350
rect 43150 550294 43218 550350
rect 43274 550294 43342 550350
rect 43398 550294 43494 550350
rect 42874 550226 43494 550294
rect 42874 550170 42970 550226
rect 43026 550170 43094 550226
rect 43150 550170 43218 550226
rect 43274 550170 43342 550226
rect 43398 550170 43494 550226
rect 42874 550102 43494 550170
rect 42874 550046 42970 550102
rect 43026 550046 43094 550102
rect 43150 550046 43218 550102
rect 43274 550046 43342 550102
rect 43398 550046 43494 550102
rect 42874 549978 43494 550046
rect 42874 549922 42970 549978
rect 43026 549922 43094 549978
rect 43150 549922 43218 549978
rect 43274 549922 43342 549978
rect 43398 549922 43494 549978
rect 42874 532350 43494 549922
rect 42874 532294 42970 532350
rect 43026 532294 43094 532350
rect 43150 532294 43218 532350
rect 43274 532294 43342 532350
rect 43398 532294 43494 532350
rect 42874 532226 43494 532294
rect 42874 532170 42970 532226
rect 43026 532170 43094 532226
rect 43150 532170 43218 532226
rect 43274 532170 43342 532226
rect 43398 532170 43494 532226
rect 42874 532102 43494 532170
rect 42874 532046 42970 532102
rect 43026 532046 43094 532102
rect 43150 532046 43218 532102
rect 43274 532046 43342 532102
rect 43398 532046 43494 532102
rect 42874 531978 43494 532046
rect 42874 531922 42970 531978
rect 43026 531922 43094 531978
rect 43150 531922 43218 531978
rect 43274 531922 43342 531978
rect 43398 531922 43494 531978
rect 42874 514350 43494 531922
rect 42874 514294 42970 514350
rect 43026 514294 43094 514350
rect 43150 514294 43218 514350
rect 43274 514294 43342 514350
rect 43398 514294 43494 514350
rect 42874 514226 43494 514294
rect 42874 514170 42970 514226
rect 43026 514170 43094 514226
rect 43150 514170 43218 514226
rect 43274 514170 43342 514226
rect 43398 514170 43494 514226
rect 42874 514102 43494 514170
rect 42874 514046 42970 514102
rect 43026 514046 43094 514102
rect 43150 514046 43218 514102
rect 43274 514046 43342 514102
rect 43398 514046 43494 514102
rect 42874 513978 43494 514046
rect 42874 513922 42970 513978
rect 43026 513922 43094 513978
rect 43150 513922 43218 513978
rect 43274 513922 43342 513978
rect 43398 513922 43494 513978
rect 42874 496350 43494 513922
rect 42874 496294 42970 496350
rect 43026 496294 43094 496350
rect 43150 496294 43218 496350
rect 43274 496294 43342 496350
rect 43398 496294 43494 496350
rect 42874 496226 43494 496294
rect 42874 496170 42970 496226
rect 43026 496170 43094 496226
rect 43150 496170 43218 496226
rect 43274 496170 43342 496226
rect 43398 496170 43494 496226
rect 42874 496102 43494 496170
rect 42874 496046 42970 496102
rect 43026 496046 43094 496102
rect 43150 496046 43218 496102
rect 43274 496046 43342 496102
rect 43398 496046 43494 496102
rect 42874 495978 43494 496046
rect 42874 495922 42970 495978
rect 43026 495922 43094 495978
rect 43150 495922 43218 495978
rect 43274 495922 43342 495978
rect 43398 495922 43494 495978
rect 42874 478350 43494 495922
rect 42874 478294 42970 478350
rect 43026 478294 43094 478350
rect 43150 478294 43218 478350
rect 43274 478294 43342 478350
rect 43398 478294 43494 478350
rect 42874 478226 43494 478294
rect 42874 478170 42970 478226
rect 43026 478170 43094 478226
rect 43150 478170 43218 478226
rect 43274 478170 43342 478226
rect 43398 478170 43494 478226
rect 42874 478102 43494 478170
rect 42874 478046 42970 478102
rect 43026 478046 43094 478102
rect 43150 478046 43218 478102
rect 43274 478046 43342 478102
rect 43398 478046 43494 478102
rect 42874 477978 43494 478046
rect 42874 477922 42970 477978
rect 43026 477922 43094 477978
rect 43150 477922 43218 477978
rect 43274 477922 43342 477978
rect 43398 477922 43494 477978
rect 42874 460350 43494 477922
rect 42874 460294 42970 460350
rect 43026 460294 43094 460350
rect 43150 460294 43218 460350
rect 43274 460294 43342 460350
rect 43398 460294 43494 460350
rect 42874 460226 43494 460294
rect 42874 460170 42970 460226
rect 43026 460170 43094 460226
rect 43150 460170 43218 460226
rect 43274 460170 43342 460226
rect 43398 460170 43494 460226
rect 42874 460102 43494 460170
rect 42874 460046 42970 460102
rect 43026 460046 43094 460102
rect 43150 460046 43218 460102
rect 43274 460046 43342 460102
rect 43398 460046 43494 460102
rect 42874 459978 43494 460046
rect 42874 459922 42970 459978
rect 43026 459922 43094 459978
rect 43150 459922 43218 459978
rect 43274 459922 43342 459978
rect 43398 459922 43494 459978
rect 42874 458342 43494 459922
rect 57154 597212 57774 598268
rect 57154 597156 57250 597212
rect 57306 597156 57374 597212
rect 57430 597156 57498 597212
rect 57554 597156 57622 597212
rect 57678 597156 57774 597212
rect 57154 597088 57774 597156
rect 57154 597032 57250 597088
rect 57306 597032 57374 597088
rect 57430 597032 57498 597088
rect 57554 597032 57622 597088
rect 57678 597032 57774 597088
rect 57154 596964 57774 597032
rect 57154 596908 57250 596964
rect 57306 596908 57374 596964
rect 57430 596908 57498 596964
rect 57554 596908 57622 596964
rect 57678 596908 57774 596964
rect 57154 596840 57774 596908
rect 57154 596784 57250 596840
rect 57306 596784 57374 596840
rect 57430 596784 57498 596840
rect 57554 596784 57622 596840
rect 57678 596784 57774 596840
rect 57154 580350 57774 596784
rect 57154 580294 57250 580350
rect 57306 580294 57374 580350
rect 57430 580294 57498 580350
rect 57554 580294 57622 580350
rect 57678 580294 57774 580350
rect 57154 580226 57774 580294
rect 57154 580170 57250 580226
rect 57306 580170 57374 580226
rect 57430 580170 57498 580226
rect 57554 580170 57622 580226
rect 57678 580170 57774 580226
rect 57154 580102 57774 580170
rect 57154 580046 57250 580102
rect 57306 580046 57374 580102
rect 57430 580046 57498 580102
rect 57554 580046 57622 580102
rect 57678 580046 57774 580102
rect 57154 579978 57774 580046
rect 57154 579922 57250 579978
rect 57306 579922 57374 579978
rect 57430 579922 57498 579978
rect 57554 579922 57622 579978
rect 57678 579922 57774 579978
rect 57154 562350 57774 579922
rect 57154 562294 57250 562350
rect 57306 562294 57374 562350
rect 57430 562294 57498 562350
rect 57554 562294 57622 562350
rect 57678 562294 57774 562350
rect 57154 562226 57774 562294
rect 57154 562170 57250 562226
rect 57306 562170 57374 562226
rect 57430 562170 57498 562226
rect 57554 562170 57622 562226
rect 57678 562170 57774 562226
rect 57154 562102 57774 562170
rect 57154 562046 57250 562102
rect 57306 562046 57374 562102
rect 57430 562046 57498 562102
rect 57554 562046 57622 562102
rect 57678 562046 57774 562102
rect 57154 561978 57774 562046
rect 57154 561922 57250 561978
rect 57306 561922 57374 561978
rect 57430 561922 57498 561978
rect 57554 561922 57622 561978
rect 57678 561922 57774 561978
rect 57154 544350 57774 561922
rect 57154 544294 57250 544350
rect 57306 544294 57374 544350
rect 57430 544294 57498 544350
rect 57554 544294 57622 544350
rect 57678 544294 57774 544350
rect 57154 544226 57774 544294
rect 57154 544170 57250 544226
rect 57306 544170 57374 544226
rect 57430 544170 57498 544226
rect 57554 544170 57622 544226
rect 57678 544170 57774 544226
rect 57154 544102 57774 544170
rect 57154 544046 57250 544102
rect 57306 544046 57374 544102
rect 57430 544046 57498 544102
rect 57554 544046 57622 544102
rect 57678 544046 57774 544102
rect 57154 543978 57774 544046
rect 57154 543922 57250 543978
rect 57306 543922 57374 543978
rect 57430 543922 57498 543978
rect 57554 543922 57622 543978
rect 57678 543922 57774 543978
rect 57154 526350 57774 543922
rect 57154 526294 57250 526350
rect 57306 526294 57374 526350
rect 57430 526294 57498 526350
rect 57554 526294 57622 526350
rect 57678 526294 57774 526350
rect 57154 526226 57774 526294
rect 57154 526170 57250 526226
rect 57306 526170 57374 526226
rect 57430 526170 57498 526226
rect 57554 526170 57622 526226
rect 57678 526170 57774 526226
rect 57154 526102 57774 526170
rect 57154 526046 57250 526102
rect 57306 526046 57374 526102
rect 57430 526046 57498 526102
rect 57554 526046 57622 526102
rect 57678 526046 57774 526102
rect 57154 525978 57774 526046
rect 57154 525922 57250 525978
rect 57306 525922 57374 525978
rect 57430 525922 57498 525978
rect 57554 525922 57622 525978
rect 57678 525922 57774 525978
rect 57154 508350 57774 525922
rect 57154 508294 57250 508350
rect 57306 508294 57374 508350
rect 57430 508294 57498 508350
rect 57554 508294 57622 508350
rect 57678 508294 57774 508350
rect 57154 508226 57774 508294
rect 57154 508170 57250 508226
rect 57306 508170 57374 508226
rect 57430 508170 57498 508226
rect 57554 508170 57622 508226
rect 57678 508170 57774 508226
rect 57154 508102 57774 508170
rect 57154 508046 57250 508102
rect 57306 508046 57374 508102
rect 57430 508046 57498 508102
rect 57554 508046 57622 508102
rect 57678 508046 57774 508102
rect 57154 507978 57774 508046
rect 57154 507922 57250 507978
rect 57306 507922 57374 507978
rect 57430 507922 57498 507978
rect 57554 507922 57622 507978
rect 57678 507922 57774 507978
rect 57154 490350 57774 507922
rect 57154 490294 57250 490350
rect 57306 490294 57374 490350
rect 57430 490294 57498 490350
rect 57554 490294 57622 490350
rect 57678 490294 57774 490350
rect 57154 490226 57774 490294
rect 57154 490170 57250 490226
rect 57306 490170 57374 490226
rect 57430 490170 57498 490226
rect 57554 490170 57622 490226
rect 57678 490170 57774 490226
rect 57154 490102 57774 490170
rect 57154 490046 57250 490102
rect 57306 490046 57374 490102
rect 57430 490046 57498 490102
rect 57554 490046 57622 490102
rect 57678 490046 57774 490102
rect 57154 489978 57774 490046
rect 57154 489922 57250 489978
rect 57306 489922 57374 489978
rect 57430 489922 57498 489978
rect 57554 489922 57622 489978
rect 57678 489922 57774 489978
rect 57154 472350 57774 489922
rect 57154 472294 57250 472350
rect 57306 472294 57374 472350
rect 57430 472294 57498 472350
rect 57554 472294 57622 472350
rect 57678 472294 57774 472350
rect 57154 472226 57774 472294
rect 57154 472170 57250 472226
rect 57306 472170 57374 472226
rect 57430 472170 57498 472226
rect 57554 472170 57622 472226
rect 57678 472170 57774 472226
rect 57154 472102 57774 472170
rect 57154 472046 57250 472102
rect 57306 472046 57374 472102
rect 57430 472046 57498 472102
rect 57554 472046 57622 472102
rect 57678 472046 57774 472102
rect 57154 471978 57774 472046
rect 57154 471922 57250 471978
rect 57306 471922 57374 471978
rect 57430 471922 57498 471978
rect 57554 471922 57622 471978
rect 57678 471922 57774 471978
rect 57154 458342 57774 471922
rect 60874 598172 61494 598268
rect 60874 598116 60970 598172
rect 61026 598116 61094 598172
rect 61150 598116 61218 598172
rect 61274 598116 61342 598172
rect 61398 598116 61494 598172
rect 60874 598048 61494 598116
rect 60874 597992 60970 598048
rect 61026 597992 61094 598048
rect 61150 597992 61218 598048
rect 61274 597992 61342 598048
rect 61398 597992 61494 598048
rect 60874 597924 61494 597992
rect 60874 597868 60970 597924
rect 61026 597868 61094 597924
rect 61150 597868 61218 597924
rect 61274 597868 61342 597924
rect 61398 597868 61494 597924
rect 60874 597800 61494 597868
rect 60874 597744 60970 597800
rect 61026 597744 61094 597800
rect 61150 597744 61218 597800
rect 61274 597744 61342 597800
rect 61398 597744 61494 597800
rect 60874 586350 61494 597744
rect 60874 586294 60970 586350
rect 61026 586294 61094 586350
rect 61150 586294 61218 586350
rect 61274 586294 61342 586350
rect 61398 586294 61494 586350
rect 60874 586226 61494 586294
rect 60874 586170 60970 586226
rect 61026 586170 61094 586226
rect 61150 586170 61218 586226
rect 61274 586170 61342 586226
rect 61398 586170 61494 586226
rect 60874 586102 61494 586170
rect 60874 586046 60970 586102
rect 61026 586046 61094 586102
rect 61150 586046 61218 586102
rect 61274 586046 61342 586102
rect 61398 586046 61494 586102
rect 60874 585978 61494 586046
rect 60874 585922 60970 585978
rect 61026 585922 61094 585978
rect 61150 585922 61218 585978
rect 61274 585922 61342 585978
rect 61398 585922 61494 585978
rect 60874 568350 61494 585922
rect 60874 568294 60970 568350
rect 61026 568294 61094 568350
rect 61150 568294 61218 568350
rect 61274 568294 61342 568350
rect 61398 568294 61494 568350
rect 60874 568226 61494 568294
rect 60874 568170 60970 568226
rect 61026 568170 61094 568226
rect 61150 568170 61218 568226
rect 61274 568170 61342 568226
rect 61398 568170 61494 568226
rect 60874 568102 61494 568170
rect 60874 568046 60970 568102
rect 61026 568046 61094 568102
rect 61150 568046 61218 568102
rect 61274 568046 61342 568102
rect 61398 568046 61494 568102
rect 60874 567978 61494 568046
rect 60874 567922 60970 567978
rect 61026 567922 61094 567978
rect 61150 567922 61218 567978
rect 61274 567922 61342 567978
rect 61398 567922 61494 567978
rect 60874 550350 61494 567922
rect 60874 550294 60970 550350
rect 61026 550294 61094 550350
rect 61150 550294 61218 550350
rect 61274 550294 61342 550350
rect 61398 550294 61494 550350
rect 60874 550226 61494 550294
rect 60874 550170 60970 550226
rect 61026 550170 61094 550226
rect 61150 550170 61218 550226
rect 61274 550170 61342 550226
rect 61398 550170 61494 550226
rect 60874 550102 61494 550170
rect 60874 550046 60970 550102
rect 61026 550046 61094 550102
rect 61150 550046 61218 550102
rect 61274 550046 61342 550102
rect 61398 550046 61494 550102
rect 60874 549978 61494 550046
rect 60874 549922 60970 549978
rect 61026 549922 61094 549978
rect 61150 549922 61218 549978
rect 61274 549922 61342 549978
rect 61398 549922 61494 549978
rect 60874 532350 61494 549922
rect 60874 532294 60970 532350
rect 61026 532294 61094 532350
rect 61150 532294 61218 532350
rect 61274 532294 61342 532350
rect 61398 532294 61494 532350
rect 60874 532226 61494 532294
rect 60874 532170 60970 532226
rect 61026 532170 61094 532226
rect 61150 532170 61218 532226
rect 61274 532170 61342 532226
rect 61398 532170 61494 532226
rect 60874 532102 61494 532170
rect 60874 532046 60970 532102
rect 61026 532046 61094 532102
rect 61150 532046 61218 532102
rect 61274 532046 61342 532102
rect 61398 532046 61494 532102
rect 60874 531978 61494 532046
rect 60874 531922 60970 531978
rect 61026 531922 61094 531978
rect 61150 531922 61218 531978
rect 61274 531922 61342 531978
rect 61398 531922 61494 531978
rect 60874 514350 61494 531922
rect 60874 514294 60970 514350
rect 61026 514294 61094 514350
rect 61150 514294 61218 514350
rect 61274 514294 61342 514350
rect 61398 514294 61494 514350
rect 60874 514226 61494 514294
rect 60874 514170 60970 514226
rect 61026 514170 61094 514226
rect 61150 514170 61218 514226
rect 61274 514170 61342 514226
rect 61398 514170 61494 514226
rect 60874 514102 61494 514170
rect 60874 514046 60970 514102
rect 61026 514046 61094 514102
rect 61150 514046 61218 514102
rect 61274 514046 61342 514102
rect 61398 514046 61494 514102
rect 60874 513978 61494 514046
rect 60874 513922 60970 513978
rect 61026 513922 61094 513978
rect 61150 513922 61218 513978
rect 61274 513922 61342 513978
rect 61398 513922 61494 513978
rect 60874 496350 61494 513922
rect 60874 496294 60970 496350
rect 61026 496294 61094 496350
rect 61150 496294 61218 496350
rect 61274 496294 61342 496350
rect 61398 496294 61494 496350
rect 60874 496226 61494 496294
rect 60874 496170 60970 496226
rect 61026 496170 61094 496226
rect 61150 496170 61218 496226
rect 61274 496170 61342 496226
rect 61398 496170 61494 496226
rect 60874 496102 61494 496170
rect 60874 496046 60970 496102
rect 61026 496046 61094 496102
rect 61150 496046 61218 496102
rect 61274 496046 61342 496102
rect 61398 496046 61494 496102
rect 60874 495978 61494 496046
rect 60874 495922 60970 495978
rect 61026 495922 61094 495978
rect 61150 495922 61218 495978
rect 61274 495922 61342 495978
rect 61398 495922 61494 495978
rect 60874 478350 61494 495922
rect 60874 478294 60970 478350
rect 61026 478294 61094 478350
rect 61150 478294 61218 478350
rect 61274 478294 61342 478350
rect 61398 478294 61494 478350
rect 60874 478226 61494 478294
rect 60874 478170 60970 478226
rect 61026 478170 61094 478226
rect 61150 478170 61218 478226
rect 61274 478170 61342 478226
rect 61398 478170 61494 478226
rect 60874 478102 61494 478170
rect 60874 478046 60970 478102
rect 61026 478046 61094 478102
rect 61150 478046 61218 478102
rect 61274 478046 61342 478102
rect 61398 478046 61494 478102
rect 60874 477978 61494 478046
rect 60874 477922 60970 477978
rect 61026 477922 61094 477978
rect 61150 477922 61218 477978
rect 61274 477922 61342 477978
rect 61398 477922 61494 477978
rect 60874 460350 61494 477922
rect 60874 460294 60970 460350
rect 61026 460294 61094 460350
rect 61150 460294 61218 460350
rect 61274 460294 61342 460350
rect 61398 460294 61494 460350
rect 60874 460226 61494 460294
rect 60874 460170 60970 460226
rect 61026 460170 61094 460226
rect 61150 460170 61218 460226
rect 61274 460170 61342 460226
rect 61398 460170 61494 460226
rect 60874 460102 61494 460170
rect 60874 460046 60970 460102
rect 61026 460046 61094 460102
rect 61150 460046 61218 460102
rect 61274 460046 61342 460102
rect 61398 460046 61494 460102
rect 60874 459978 61494 460046
rect 60874 459922 60970 459978
rect 61026 459922 61094 459978
rect 61150 459922 61218 459978
rect 61274 459922 61342 459978
rect 61398 459922 61494 459978
rect 60874 458342 61494 459922
rect 75154 597212 75774 598268
rect 75154 597156 75250 597212
rect 75306 597156 75374 597212
rect 75430 597156 75498 597212
rect 75554 597156 75622 597212
rect 75678 597156 75774 597212
rect 75154 597088 75774 597156
rect 75154 597032 75250 597088
rect 75306 597032 75374 597088
rect 75430 597032 75498 597088
rect 75554 597032 75622 597088
rect 75678 597032 75774 597088
rect 75154 596964 75774 597032
rect 75154 596908 75250 596964
rect 75306 596908 75374 596964
rect 75430 596908 75498 596964
rect 75554 596908 75622 596964
rect 75678 596908 75774 596964
rect 75154 596840 75774 596908
rect 75154 596784 75250 596840
rect 75306 596784 75374 596840
rect 75430 596784 75498 596840
rect 75554 596784 75622 596840
rect 75678 596784 75774 596840
rect 75154 580350 75774 596784
rect 75154 580294 75250 580350
rect 75306 580294 75374 580350
rect 75430 580294 75498 580350
rect 75554 580294 75622 580350
rect 75678 580294 75774 580350
rect 75154 580226 75774 580294
rect 75154 580170 75250 580226
rect 75306 580170 75374 580226
rect 75430 580170 75498 580226
rect 75554 580170 75622 580226
rect 75678 580170 75774 580226
rect 75154 580102 75774 580170
rect 75154 580046 75250 580102
rect 75306 580046 75374 580102
rect 75430 580046 75498 580102
rect 75554 580046 75622 580102
rect 75678 580046 75774 580102
rect 75154 579978 75774 580046
rect 75154 579922 75250 579978
rect 75306 579922 75374 579978
rect 75430 579922 75498 579978
rect 75554 579922 75622 579978
rect 75678 579922 75774 579978
rect 75154 562350 75774 579922
rect 75154 562294 75250 562350
rect 75306 562294 75374 562350
rect 75430 562294 75498 562350
rect 75554 562294 75622 562350
rect 75678 562294 75774 562350
rect 75154 562226 75774 562294
rect 75154 562170 75250 562226
rect 75306 562170 75374 562226
rect 75430 562170 75498 562226
rect 75554 562170 75622 562226
rect 75678 562170 75774 562226
rect 75154 562102 75774 562170
rect 75154 562046 75250 562102
rect 75306 562046 75374 562102
rect 75430 562046 75498 562102
rect 75554 562046 75622 562102
rect 75678 562046 75774 562102
rect 75154 561978 75774 562046
rect 75154 561922 75250 561978
rect 75306 561922 75374 561978
rect 75430 561922 75498 561978
rect 75554 561922 75622 561978
rect 75678 561922 75774 561978
rect 75154 544350 75774 561922
rect 75154 544294 75250 544350
rect 75306 544294 75374 544350
rect 75430 544294 75498 544350
rect 75554 544294 75622 544350
rect 75678 544294 75774 544350
rect 75154 544226 75774 544294
rect 75154 544170 75250 544226
rect 75306 544170 75374 544226
rect 75430 544170 75498 544226
rect 75554 544170 75622 544226
rect 75678 544170 75774 544226
rect 75154 544102 75774 544170
rect 75154 544046 75250 544102
rect 75306 544046 75374 544102
rect 75430 544046 75498 544102
rect 75554 544046 75622 544102
rect 75678 544046 75774 544102
rect 75154 543978 75774 544046
rect 75154 543922 75250 543978
rect 75306 543922 75374 543978
rect 75430 543922 75498 543978
rect 75554 543922 75622 543978
rect 75678 543922 75774 543978
rect 75154 526350 75774 543922
rect 75154 526294 75250 526350
rect 75306 526294 75374 526350
rect 75430 526294 75498 526350
rect 75554 526294 75622 526350
rect 75678 526294 75774 526350
rect 75154 526226 75774 526294
rect 75154 526170 75250 526226
rect 75306 526170 75374 526226
rect 75430 526170 75498 526226
rect 75554 526170 75622 526226
rect 75678 526170 75774 526226
rect 75154 526102 75774 526170
rect 75154 526046 75250 526102
rect 75306 526046 75374 526102
rect 75430 526046 75498 526102
rect 75554 526046 75622 526102
rect 75678 526046 75774 526102
rect 75154 525978 75774 526046
rect 75154 525922 75250 525978
rect 75306 525922 75374 525978
rect 75430 525922 75498 525978
rect 75554 525922 75622 525978
rect 75678 525922 75774 525978
rect 75154 508350 75774 525922
rect 75154 508294 75250 508350
rect 75306 508294 75374 508350
rect 75430 508294 75498 508350
rect 75554 508294 75622 508350
rect 75678 508294 75774 508350
rect 75154 508226 75774 508294
rect 75154 508170 75250 508226
rect 75306 508170 75374 508226
rect 75430 508170 75498 508226
rect 75554 508170 75622 508226
rect 75678 508170 75774 508226
rect 75154 508102 75774 508170
rect 75154 508046 75250 508102
rect 75306 508046 75374 508102
rect 75430 508046 75498 508102
rect 75554 508046 75622 508102
rect 75678 508046 75774 508102
rect 75154 507978 75774 508046
rect 75154 507922 75250 507978
rect 75306 507922 75374 507978
rect 75430 507922 75498 507978
rect 75554 507922 75622 507978
rect 75678 507922 75774 507978
rect 75154 490350 75774 507922
rect 75154 490294 75250 490350
rect 75306 490294 75374 490350
rect 75430 490294 75498 490350
rect 75554 490294 75622 490350
rect 75678 490294 75774 490350
rect 75154 490226 75774 490294
rect 75154 490170 75250 490226
rect 75306 490170 75374 490226
rect 75430 490170 75498 490226
rect 75554 490170 75622 490226
rect 75678 490170 75774 490226
rect 75154 490102 75774 490170
rect 75154 490046 75250 490102
rect 75306 490046 75374 490102
rect 75430 490046 75498 490102
rect 75554 490046 75622 490102
rect 75678 490046 75774 490102
rect 75154 489978 75774 490046
rect 75154 489922 75250 489978
rect 75306 489922 75374 489978
rect 75430 489922 75498 489978
rect 75554 489922 75622 489978
rect 75678 489922 75774 489978
rect 75154 472350 75774 489922
rect 75154 472294 75250 472350
rect 75306 472294 75374 472350
rect 75430 472294 75498 472350
rect 75554 472294 75622 472350
rect 75678 472294 75774 472350
rect 75154 472226 75774 472294
rect 75154 472170 75250 472226
rect 75306 472170 75374 472226
rect 75430 472170 75498 472226
rect 75554 472170 75622 472226
rect 75678 472170 75774 472226
rect 75154 472102 75774 472170
rect 75154 472046 75250 472102
rect 75306 472046 75374 472102
rect 75430 472046 75498 472102
rect 75554 472046 75622 472102
rect 75678 472046 75774 472102
rect 75154 471978 75774 472046
rect 75154 471922 75250 471978
rect 75306 471922 75374 471978
rect 75430 471922 75498 471978
rect 75554 471922 75622 471978
rect 75678 471922 75774 471978
rect 75154 458342 75774 471922
rect 78874 598172 79494 598268
rect 78874 598116 78970 598172
rect 79026 598116 79094 598172
rect 79150 598116 79218 598172
rect 79274 598116 79342 598172
rect 79398 598116 79494 598172
rect 78874 598048 79494 598116
rect 78874 597992 78970 598048
rect 79026 597992 79094 598048
rect 79150 597992 79218 598048
rect 79274 597992 79342 598048
rect 79398 597992 79494 598048
rect 78874 597924 79494 597992
rect 78874 597868 78970 597924
rect 79026 597868 79094 597924
rect 79150 597868 79218 597924
rect 79274 597868 79342 597924
rect 79398 597868 79494 597924
rect 78874 597800 79494 597868
rect 78874 597744 78970 597800
rect 79026 597744 79094 597800
rect 79150 597744 79218 597800
rect 79274 597744 79342 597800
rect 79398 597744 79494 597800
rect 78874 586350 79494 597744
rect 78874 586294 78970 586350
rect 79026 586294 79094 586350
rect 79150 586294 79218 586350
rect 79274 586294 79342 586350
rect 79398 586294 79494 586350
rect 78874 586226 79494 586294
rect 78874 586170 78970 586226
rect 79026 586170 79094 586226
rect 79150 586170 79218 586226
rect 79274 586170 79342 586226
rect 79398 586170 79494 586226
rect 78874 586102 79494 586170
rect 78874 586046 78970 586102
rect 79026 586046 79094 586102
rect 79150 586046 79218 586102
rect 79274 586046 79342 586102
rect 79398 586046 79494 586102
rect 78874 585978 79494 586046
rect 78874 585922 78970 585978
rect 79026 585922 79094 585978
rect 79150 585922 79218 585978
rect 79274 585922 79342 585978
rect 79398 585922 79494 585978
rect 78874 568350 79494 585922
rect 78874 568294 78970 568350
rect 79026 568294 79094 568350
rect 79150 568294 79218 568350
rect 79274 568294 79342 568350
rect 79398 568294 79494 568350
rect 78874 568226 79494 568294
rect 78874 568170 78970 568226
rect 79026 568170 79094 568226
rect 79150 568170 79218 568226
rect 79274 568170 79342 568226
rect 79398 568170 79494 568226
rect 78874 568102 79494 568170
rect 78874 568046 78970 568102
rect 79026 568046 79094 568102
rect 79150 568046 79218 568102
rect 79274 568046 79342 568102
rect 79398 568046 79494 568102
rect 78874 567978 79494 568046
rect 78874 567922 78970 567978
rect 79026 567922 79094 567978
rect 79150 567922 79218 567978
rect 79274 567922 79342 567978
rect 79398 567922 79494 567978
rect 78874 550350 79494 567922
rect 78874 550294 78970 550350
rect 79026 550294 79094 550350
rect 79150 550294 79218 550350
rect 79274 550294 79342 550350
rect 79398 550294 79494 550350
rect 78874 550226 79494 550294
rect 78874 550170 78970 550226
rect 79026 550170 79094 550226
rect 79150 550170 79218 550226
rect 79274 550170 79342 550226
rect 79398 550170 79494 550226
rect 78874 550102 79494 550170
rect 78874 550046 78970 550102
rect 79026 550046 79094 550102
rect 79150 550046 79218 550102
rect 79274 550046 79342 550102
rect 79398 550046 79494 550102
rect 78874 549978 79494 550046
rect 78874 549922 78970 549978
rect 79026 549922 79094 549978
rect 79150 549922 79218 549978
rect 79274 549922 79342 549978
rect 79398 549922 79494 549978
rect 78874 532350 79494 549922
rect 78874 532294 78970 532350
rect 79026 532294 79094 532350
rect 79150 532294 79218 532350
rect 79274 532294 79342 532350
rect 79398 532294 79494 532350
rect 78874 532226 79494 532294
rect 78874 532170 78970 532226
rect 79026 532170 79094 532226
rect 79150 532170 79218 532226
rect 79274 532170 79342 532226
rect 79398 532170 79494 532226
rect 78874 532102 79494 532170
rect 78874 532046 78970 532102
rect 79026 532046 79094 532102
rect 79150 532046 79218 532102
rect 79274 532046 79342 532102
rect 79398 532046 79494 532102
rect 78874 531978 79494 532046
rect 78874 531922 78970 531978
rect 79026 531922 79094 531978
rect 79150 531922 79218 531978
rect 79274 531922 79342 531978
rect 79398 531922 79494 531978
rect 78874 514350 79494 531922
rect 78874 514294 78970 514350
rect 79026 514294 79094 514350
rect 79150 514294 79218 514350
rect 79274 514294 79342 514350
rect 79398 514294 79494 514350
rect 78874 514226 79494 514294
rect 78874 514170 78970 514226
rect 79026 514170 79094 514226
rect 79150 514170 79218 514226
rect 79274 514170 79342 514226
rect 79398 514170 79494 514226
rect 78874 514102 79494 514170
rect 78874 514046 78970 514102
rect 79026 514046 79094 514102
rect 79150 514046 79218 514102
rect 79274 514046 79342 514102
rect 79398 514046 79494 514102
rect 78874 513978 79494 514046
rect 78874 513922 78970 513978
rect 79026 513922 79094 513978
rect 79150 513922 79218 513978
rect 79274 513922 79342 513978
rect 79398 513922 79494 513978
rect 78874 496350 79494 513922
rect 78874 496294 78970 496350
rect 79026 496294 79094 496350
rect 79150 496294 79218 496350
rect 79274 496294 79342 496350
rect 79398 496294 79494 496350
rect 78874 496226 79494 496294
rect 78874 496170 78970 496226
rect 79026 496170 79094 496226
rect 79150 496170 79218 496226
rect 79274 496170 79342 496226
rect 79398 496170 79494 496226
rect 78874 496102 79494 496170
rect 78874 496046 78970 496102
rect 79026 496046 79094 496102
rect 79150 496046 79218 496102
rect 79274 496046 79342 496102
rect 79398 496046 79494 496102
rect 78874 495978 79494 496046
rect 78874 495922 78970 495978
rect 79026 495922 79094 495978
rect 79150 495922 79218 495978
rect 79274 495922 79342 495978
rect 79398 495922 79494 495978
rect 78874 478350 79494 495922
rect 78874 478294 78970 478350
rect 79026 478294 79094 478350
rect 79150 478294 79218 478350
rect 79274 478294 79342 478350
rect 79398 478294 79494 478350
rect 78874 478226 79494 478294
rect 78874 478170 78970 478226
rect 79026 478170 79094 478226
rect 79150 478170 79218 478226
rect 79274 478170 79342 478226
rect 79398 478170 79494 478226
rect 78874 478102 79494 478170
rect 78874 478046 78970 478102
rect 79026 478046 79094 478102
rect 79150 478046 79218 478102
rect 79274 478046 79342 478102
rect 79398 478046 79494 478102
rect 78874 477978 79494 478046
rect 78874 477922 78970 477978
rect 79026 477922 79094 477978
rect 79150 477922 79218 477978
rect 79274 477922 79342 477978
rect 79398 477922 79494 477978
rect 78874 460350 79494 477922
rect 78874 460294 78970 460350
rect 79026 460294 79094 460350
rect 79150 460294 79218 460350
rect 79274 460294 79342 460350
rect 79398 460294 79494 460350
rect 78874 460226 79494 460294
rect 78874 460170 78970 460226
rect 79026 460170 79094 460226
rect 79150 460170 79218 460226
rect 79274 460170 79342 460226
rect 79398 460170 79494 460226
rect 78874 460102 79494 460170
rect 78874 460046 78970 460102
rect 79026 460046 79094 460102
rect 79150 460046 79218 460102
rect 79274 460046 79342 460102
rect 79398 460046 79494 460102
rect 78874 459978 79494 460046
rect 78874 459922 78970 459978
rect 79026 459922 79094 459978
rect 79150 459922 79218 459978
rect 79274 459922 79342 459978
rect 79398 459922 79494 459978
rect 78874 458342 79494 459922
rect 93154 597212 93774 598268
rect 93154 597156 93250 597212
rect 93306 597156 93374 597212
rect 93430 597156 93498 597212
rect 93554 597156 93622 597212
rect 93678 597156 93774 597212
rect 93154 597088 93774 597156
rect 93154 597032 93250 597088
rect 93306 597032 93374 597088
rect 93430 597032 93498 597088
rect 93554 597032 93622 597088
rect 93678 597032 93774 597088
rect 93154 596964 93774 597032
rect 93154 596908 93250 596964
rect 93306 596908 93374 596964
rect 93430 596908 93498 596964
rect 93554 596908 93622 596964
rect 93678 596908 93774 596964
rect 93154 596840 93774 596908
rect 93154 596784 93250 596840
rect 93306 596784 93374 596840
rect 93430 596784 93498 596840
rect 93554 596784 93622 596840
rect 93678 596784 93774 596840
rect 93154 580350 93774 596784
rect 93154 580294 93250 580350
rect 93306 580294 93374 580350
rect 93430 580294 93498 580350
rect 93554 580294 93622 580350
rect 93678 580294 93774 580350
rect 93154 580226 93774 580294
rect 93154 580170 93250 580226
rect 93306 580170 93374 580226
rect 93430 580170 93498 580226
rect 93554 580170 93622 580226
rect 93678 580170 93774 580226
rect 93154 580102 93774 580170
rect 93154 580046 93250 580102
rect 93306 580046 93374 580102
rect 93430 580046 93498 580102
rect 93554 580046 93622 580102
rect 93678 580046 93774 580102
rect 93154 579978 93774 580046
rect 93154 579922 93250 579978
rect 93306 579922 93374 579978
rect 93430 579922 93498 579978
rect 93554 579922 93622 579978
rect 93678 579922 93774 579978
rect 93154 562350 93774 579922
rect 93154 562294 93250 562350
rect 93306 562294 93374 562350
rect 93430 562294 93498 562350
rect 93554 562294 93622 562350
rect 93678 562294 93774 562350
rect 93154 562226 93774 562294
rect 93154 562170 93250 562226
rect 93306 562170 93374 562226
rect 93430 562170 93498 562226
rect 93554 562170 93622 562226
rect 93678 562170 93774 562226
rect 93154 562102 93774 562170
rect 93154 562046 93250 562102
rect 93306 562046 93374 562102
rect 93430 562046 93498 562102
rect 93554 562046 93622 562102
rect 93678 562046 93774 562102
rect 93154 561978 93774 562046
rect 93154 561922 93250 561978
rect 93306 561922 93374 561978
rect 93430 561922 93498 561978
rect 93554 561922 93622 561978
rect 93678 561922 93774 561978
rect 93154 544350 93774 561922
rect 93154 544294 93250 544350
rect 93306 544294 93374 544350
rect 93430 544294 93498 544350
rect 93554 544294 93622 544350
rect 93678 544294 93774 544350
rect 93154 544226 93774 544294
rect 93154 544170 93250 544226
rect 93306 544170 93374 544226
rect 93430 544170 93498 544226
rect 93554 544170 93622 544226
rect 93678 544170 93774 544226
rect 93154 544102 93774 544170
rect 93154 544046 93250 544102
rect 93306 544046 93374 544102
rect 93430 544046 93498 544102
rect 93554 544046 93622 544102
rect 93678 544046 93774 544102
rect 93154 543978 93774 544046
rect 93154 543922 93250 543978
rect 93306 543922 93374 543978
rect 93430 543922 93498 543978
rect 93554 543922 93622 543978
rect 93678 543922 93774 543978
rect 93154 526350 93774 543922
rect 93154 526294 93250 526350
rect 93306 526294 93374 526350
rect 93430 526294 93498 526350
rect 93554 526294 93622 526350
rect 93678 526294 93774 526350
rect 93154 526226 93774 526294
rect 93154 526170 93250 526226
rect 93306 526170 93374 526226
rect 93430 526170 93498 526226
rect 93554 526170 93622 526226
rect 93678 526170 93774 526226
rect 93154 526102 93774 526170
rect 93154 526046 93250 526102
rect 93306 526046 93374 526102
rect 93430 526046 93498 526102
rect 93554 526046 93622 526102
rect 93678 526046 93774 526102
rect 93154 525978 93774 526046
rect 93154 525922 93250 525978
rect 93306 525922 93374 525978
rect 93430 525922 93498 525978
rect 93554 525922 93622 525978
rect 93678 525922 93774 525978
rect 93154 508350 93774 525922
rect 93154 508294 93250 508350
rect 93306 508294 93374 508350
rect 93430 508294 93498 508350
rect 93554 508294 93622 508350
rect 93678 508294 93774 508350
rect 93154 508226 93774 508294
rect 93154 508170 93250 508226
rect 93306 508170 93374 508226
rect 93430 508170 93498 508226
rect 93554 508170 93622 508226
rect 93678 508170 93774 508226
rect 93154 508102 93774 508170
rect 93154 508046 93250 508102
rect 93306 508046 93374 508102
rect 93430 508046 93498 508102
rect 93554 508046 93622 508102
rect 93678 508046 93774 508102
rect 93154 507978 93774 508046
rect 93154 507922 93250 507978
rect 93306 507922 93374 507978
rect 93430 507922 93498 507978
rect 93554 507922 93622 507978
rect 93678 507922 93774 507978
rect 93154 490350 93774 507922
rect 93154 490294 93250 490350
rect 93306 490294 93374 490350
rect 93430 490294 93498 490350
rect 93554 490294 93622 490350
rect 93678 490294 93774 490350
rect 93154 490226 93774 490294
rect 93154 490170 93250 490226
rect 93306 490170 93374 490226
rect 93430 490170 93498 490226
rect 93554 490170 93622 490226
rect 93678 490170 93774 490226
rect 93154 490102 93774 490170
rect 93154 490046 93250 490102
rect 93306 490046 93374 490102
rect 93430 490046 93498 490102
rect 93554 490046 93622 490102
rect 93678 490046 93774 490102
rect 93154 489978 93774 490046
rect 93154 489922 93250 489978
rect 93306 489922 93374 489978
rect 93430 489922 93498 489978
rect 93554 489922 93622 489978
rect 93678 489922 93774 489978
rect 93154 472350 93774 489922
rect 93154 472294 93250 472350
rect 93306 472294 93374 472350
rect 93430 472294 93498 472350
rect 93554 472294 93622 472350
rect 93678 472294 93774 472350
rect 93154 472226 93774 472294
rect 93154 472170 93250 472226
rect 93306 472170 93374 472226
rect 93430 472170 93498 472226
rect 93554 472170 93622 472226
rect 93678 472170 93774 472226
rect 93154 472102 93774 472170
rect 93154 472046 93250 472102
rect 93306 472046 93374 472102
rect 93430 472046 93498 472102
rect 93554 472046 93622 472102
rect 93678 472046 93774 472102
rect 93154 471978 93774 472046
rect 93154 471922 93250 471978
rect 93306 471922 93374 471978
rect 93430 471922 93498 471978
rect 93554 471922 93622 471978
rect 93678 471922 93774 471978
rect 93154 458342 93774 471922
rect 96874 598172 97494 598268
rect 96874 598116 96970 598172
rect 97026 598116 97094 598172
rect 97150 598116 97218 598172
rect 97274 598116 97342 598172
rect 97398 598116 97494 598172
rect 96874 598048 97494 598116
rect 96874 597992 96970 598048
rect 97026 597992 97094 598048
rect 97150 597992 97218 598048
rect 97274 597992 97342 598048
rect 97398 597992 97494 598048
rect 96874 597924 97494 597992
rect 96874 597868 96970 597924
rect 97026 597868 97094 597924
rect 97150 597868 97218 597924
rect 97274 597868 97342 597924
rect 97398 597868 97494 597924
rect 96874 597800 97494 597868
rect 96874 597744 96970 597800
rect 97026 597744 97094 597800
rect 97150 597744 97218 597800
rect 97274 597744 97342 597800
rect 97398 597744 97494 597800
rect 96874 586350 97494 597744
rect 96874 586294 96970 586350
rect 97026 586294 97094 586350
rect 97150 586294 97218 586350
rect 97274 586294 97342 586350
rect 97398 586294 97494 586350
rect 96874 586226 97494 586294
rect 96874 586170 96970 586226
rect 97026 586170 97094 586226
rect 97150 586170 97218 586226
rect 97274 586170 97342 586226
rect 97398 586170 97494 586226
rect 96874 586102 97494 586170
rect 96874 586046 96970 586102
rect 97026 586046 97094 586102
rect 97150 586046 97218 586102
rect 97274 586046 97342 586102
rect 97398 586046 97494 586102
rect 96874 585978 97494 586046
rect 96874 585922 96970 585978
rect 97026 585922 97094 585978
rect 97150 585922 97218 585978
rect 97274 585922 97342 585978
rect 97398 585922 97494 585978
rect 96874 568350 97494 585922
rect 96874 568294 96970 568350
rect 97026 568294 97094 568350
rect 97150 568294 97218 568350
rect 97274 568294 97342 568350
rect 97398 568294 97494 568350
rect 96874 568226 97494 568294
rect 96874 568170 96970 568226
rect 97026 568170 97094 568226
rect 97150 568170 97218 568226
rect 97274 568170 97342 568226
rect 97398 568170 97494 568226
rect 96874 568102 97494 568170
rect 96874 568046 96970 568102
rect 97026 568046 97094 568102
rect 97150 568046 97218 568102
rect 97274 568046 97342 568102
rect 97398 568046 97494 568102
rect 96874 567978 97494 568046
rect 96874 567922 96970 567978
rect 97026 567922 97094 567978
rect 97150 567922 97218 567978
rect 97274 567922 97342 567978
rect 97398 567922 97494 567978
rect 96874 550350 97494 567922
rect 96874 550294 96970 550350
rect 97026 550294 97094 550350
rect 97150 550294 97218 550350
rect 97274 550294 97342 550350
rect 97398 550294 97494 550350
rect 96874 550226 97494 550294
rect 96874 550170 96970 550226
rect 97026 550170 97094 550226
rect 97150 550170 97218 550226
rect 97274 550170 97342 550226
rect 97398 550170 97494 550226
rect 96874 550102 97494 550170
rect 96874 550046 96970 550102
rect 97026 550046 97094 550102
rect 97150 550046 97218 550102
rect 97274 550046 97342 550102
rect 97398 550046 97494 550102
rect 96874 549978 97494 550046
rect 96874 549922 96970 549978
rect 97026 549922 97094 549978
rect 97150 549922 97218 549978
rect 97274 549922 97342 549978
rect 97398 549922 97494 549978
rect 96874 532350 97494 549922
rect 96874 532294 96970 532350
rect 97026 532294 97094 532350
rect 97150 532294 97218 532350
rect 97274 532294 97342 532350
rect 97398 532294 97494 532350
rect 96874 532226 97494 532294
rect 96874 532170 96970 532226
rect 97026 532170 97094 532226
rect 97150 532170 97218 532226
rect 97274 532170 97342 532226
rect 97398 532170 97494 532226
rect 96874 532102 97494 532170
rect 96874 532046 96970 532102
rect 97026 532046 97094 532102
rect 97150 532046 97218 532102
rect 97274 532046 97342 532102
rect 97398 532046 97494 532102
rect 96874 531978 97494 532046
rect 96874 531922 96970 531978
rect 97026 531922 97094 531978
rect 97150 531922 97218 531978
rect 97274 531922 97342 531978
rect 97398 531922 97494 531978
rect 96874 514350 97494 531922
rect 96874 514294 96970 514350
rect 97026 514294 97094 514350
rect 97150 514294 97218 514350
rect 97274 514294 97342 514350
rect 97398 514294 97494 514350
rect 96874 514226 97494 514294
rect 96874 514170 96970 514226
rect 97026 514170 97094 514226
rect 97150 514170 97218 514226
rect 97274 514170 97342 514226
rect 97398 514170 97494 514226
rect 96874 514102 97494 514170
rect 96874 514046 96970 514102
rect 97026 514046 97094 514102
rect 97150 514046 97218 514102
rect 97274 514046 97342 514102
rect 97398 514046 97494 514102
rect 96874 513978 97494 514046
rect 96874 513922 96970 513978
rect 97026 513922 97094 513978
rect 97150 513922 97218 513978
rect 97274 513922 97342 513978
rect 97398 513922 97494 513978
rect 96874 496350 97494 513922
rect 96874 496294 96970 496350
rect 97026 496294 97094 496350
rect 97150 496294 97218 496350
rect 97274 496294 97342 496350
rect 97398 496294 97494 496350
rect 96874 496226 97494 496294
rect 96874 496170 96970 496226
rect 97026 496170 97094 496226
rect 97150 496170 97218 496226
rect 97274 496170 97342 496226
rect 97398 496170 97494 496226
rect 96874 496102 97494 496170
rect 96874 496046 96970 496102
rect 97026 496046 97094 496102
rect 97150 496046 97218 496102
rect 97274 496046 97342 496102
rect 97398 496046 97494 496102
rect 96874 495978 97494 496046
rect 96874 495922 96970 495978
rect 97026 495922 97094 495978
rect 97150 495922 97218 495978
rect 97274 495922 97342 495978
rect 97398 495922 97494 495978
rect 96874 478350 97494 495922
rect 96874 478294 96970 478350
rect 97026 478294 97094 478350
rect 97150 478294 97218 478350
rect 97274 478294 97342 478350
rect 97398 478294 97494 478350
rect 96874 478226 97494 478294
rect 96874 478170 96970 478226
rect 97026 478170 97094 478226
rect 97150 478170 97218 478226
rect 97274 478170 97342 478226
rect 97398 478170 97494 478226
rect 96874 478102 97494 478170
rect 96874 478046 96970 478102
rect 97026 478046 97094 478102
rect 97150 478046 97218 478102
rect 97274 478046 97342 478102
rect 97398 478046 97494 478102
rect 96874 477978 97494 478046
rect 96874 477922 96970 477978
rect 97026 477922 97094 477978
rect 97150 477922 97218 477978
rect 97274 477922 97342 477978
rect 97398 477922 97494 477978
rect 96874 460350 97494 477922
rect 96874 460294 96970 460350
rect 97026 460294 97094 460350
rect 97150 460294 97218 460350
rect 97274 460294 97342 460350
rect 97398 460294 97494 460350
rect 96874 460226 97494 460294
rect 96874 460170 96970 460226
rect 97026 460170 97094 460226
rect 97150 460170 97218 460226
rect 97274 460170 97342 460226
rect 97398 460170 97494 460226
rect 96874 460102 97494 460170
rect 96874 460046 96970 460102
rect 97026 460046 97094 460102
rect 97150 460046 97218 460102
rect 97274 460046 97342 460102
rect 97398 460046 97494 460102
rect 96874 459978 97494 460046
rect 96874 459922 96970 459978
rect 97026 459922 97094 459978
rect 97150 459922 97218 459978
rect 97274 459922 97342 459978
rect 97398 459922 97494 459978
rect 96874 458342 97494 459922
rect 111154 597212 111774 598268
rect 111154 597156 111250 597212
rect 111306 597156 111374 597212
rect 111430 597156 111498 597212
rect 111554 597156 111622 597212
rect 111678 597156 111774 597212
rect 111154 597088 111774 597156
rect 111154 597032 111250 597088
rect 111306 597032 111374 597088
rect 111430 597032 111498 597088
rect 111554 597032 111622 597088
rect 111678 597032 111774 597088
rect 111154 596964 111774 597032
rect 111154 596908 111250 596964
rect 111306 596908 111374 596964
rect 111430 596908 111498 596964
rect 111554 596908 111622 596964
rect 111678 596908 111774 596964
rect 111154 596840 111774 596908
rect 111154 596784 111250 596840
rect 111306 596784 111374 596840
rect 111430 596784 111498 596840
rect 111554 596784 111622 596840
rect 111678 596784 111774 596840
rect 111154 580350 111774 596784
rect 111154 580294 111250 580350
rect 111306 580294 111374 580350
rect 111430 580294 111498 580350
rect 111554 580294 111622 580350
rect 111678 580294 111774 580350
rect 111154 580226 111774 580294
rect 111154 580170 111250 580226
rect 111306 580170 111374 580226
rect 111430 580170 111498 580226
rect 111554 580170 111622 580226
rect 111678 580170 111774 580226
rect 111154 580102 111774 580170
rect 111154 580046 111250 580102
rect 111306 580046 111374 580102
rect 111430 580046 111498 580102
rect 111554 580046 111622 580102
rect 111678 580046 111774 580102
rect 111154 579978 111774 580046
rect 111154 579922 111250 579978
rect 111306 579922 111374 579978
rect 111430 579922 111498 579978
rect 111554 579922 111622 579978
rect 111678 579922 111774 579978
rect 111154 562350 111774 579922
rect 111154 562294 111250 562350
rect 111306 562294 111374 562350
rect 111430 562294 111498 562350
rect 111554 562294 111622 562350
rect 111678 562294 111774 562350
rect 111154 562226 111774 562294
rect 111154 562170 111250 562226
rect 111306 562170 111374 562226
rect 111430 562170 111498 562226
rect 111554 562170 111622 562226
rect 111678 562170 111774 562226
rect 111154 562102 111774 562170
rect 111154 562046 111250 562102
rect 111306 562046 111374 562102
rect 111430 562046 111498 562102
rect 111554 562046 111622 562102
rect 111678 562046 111774 562102
rect 111154 561978 111774 562046
rect 111154 561922 111250 561978
rect 111306 561922 111374 561978
rect 111430 561922 111498 561978
rect 111554 561922 111622 561978
rect 111678 561922 111774 561978
rect 111154 544350 111774 561922
rect 111154 544294 111250 544350
rect 111306 544294 111374 544350
rect 111430 544294 111498 544350
rect 111554 544294 111622 544350
rect 111678 544294 111774 544350
rect 111154 544226 111774 544294
rect 111154 544170 111250 544226
rect 111306 544170 111374 544226
rect 111430 544170 111498 544226
rect 111554 544170 111622 544226
rect 111678 544170 111774 544226
rect 111154 544102 111774 544170
rect 111154 544046 111250 544102
rect 111306 544046 111374 544102
rect 111430 544046 111498 544102
rect 111554 544046 111622 544102
rect 111678 544046 111774 544102
rect 111154 543978 111774 544046
rect 111154 543922 111250 543978
rect 111306 543922 111374 543978
rect 111430 543922 111498 543978
rect 111554 543922 111622 543978
rect 111678 543922 111774 543978
rect 111154 526350 111774 543922
rect 111154 526294 111250 526350
rect 111306 526294 111374 526350
rect 111430 526294 111498 526350
rect 111554 526294 111622 526350
rect 111678 526294 111774 526350
rect 111154 526226 111774 526294
rect 111154 526170 111250 526226
rect 111306 526170 111374 526226
rect 111430 526170 111498 526226
rect 111554 526170 111622 526226
rect 111678 526170 111774 526226
rect 111154 526102 111774 526170
rect 111154 526046 111250 526102
rect 111306 526046 111374 526102
rect 111430 526046 111498 526102
rect 111554 526046 111622 526102
rect 111678 526046 111774 526102
rect 111154 525978 111774 526046
rect 111154 525922 111250 525978
rect 111306 525922 111374 525978
rect 111430 525922 111498 525978
rect 111554 525922 111622 525978
rect 111678 525922 111774 525978
rect 111154 508350 111774 525922
rect 111154 508294 111250 508350
rect 111306 508294 111374 508350
rect 111430 508294 111498 508350
rect 111554 508294 111622 508350
rect 111678 508294 111774 508350
rect 111154 508226 111774 508294
rect 111154 508170 111250 508226
rect 111306 508170 111374 508226
rect 111430 508170 111498 508226
rect 111554 508170 111622 508226
rect 111678 508170 111774 508226
rect 111154 508102 111774 508170
rect 111154 508046 111250 508102
rect 111306 508046 111374 508102
rect 111430 508046 111498 508102
rect 111554 508046 111622 508102
rect 111678 508046 111774 508102
rect 111154 507978 111774 508046
rect 111154 507922 111250 507978
rect 111306 507922 111374 507978
rect 111430 507922 111498 507978
rect 111554 507922 111622 507978
rect 111678 507922 111774 507978
rect 111154 490350 111774 507922
rect 111154 490294 111250 490350
rect 111306 490294 111374 490350
rect 111430 490294 111498 490350
rect 111554 490294 111622 490350
rect 111678 490294 111774 490350
rect 111154 490226 111774 490294
rect 111154 490170 111250 490226
rect 111306 490170 111374 490226
rect 111430 490170 111498 490226
rect 111554 490170 111622 490226
rect 111678 490170 111774 490226
rect 111154 490102 111774 490170
rect 111154 490046 111250 490102
rect 111306 490046 111374 490102
rect 111430 490046 111498 490102
rect 111554 490046 111622 490102
rect 111678 490046 111774 490102
rect 111154 489978 111774 490046
rect 111154 489922 111250 489978
rect 111306 489922 111374 489978
rect 111430 489922 111498 489978
rect 111554 489922 111622 489978
rect 111678 489922 111774 489978
rect 111154 472350 111774 489922
rect 111154 472294 111250 472350
rect 111306 472294 111374 472350
rect 111430 472294 111498 472350
rect 111554 472294 111622 472350
rect 111678 472294 111774 472350
rect 111154 472226 111774 472294
rect 111154 472170 111250 472226
rect 111306 472170 111374 472226
rect 111430 472170 111498 472226
rect 111554 472170 111622 472226
rect 111678 472170 111774 472226
rect 111154 472102 111774 472170
rect 111154 472046 111250 472102
rect 111306 472046 111374 472102
rect 111430 472046 111498 472102
rect 111554 472046 111622 472102
rect 111678 472046 111774 472102
rect 111154 471978 111774 472046
rect 111154 471922 111250 471978
rect 111306 471922 111374 471978
rect 111430 471922 111498 471978
rect 111554 471922 111622 471978
rect 111678 471922 111774 471978
rect 111154 458342 111774 471922
rect 114874 598172 115494 598268
rect 114874 598116 114970 598172
rect 115026 598116 115094 598172
rect 115150 598116 115218 598172
rect 115274 598116 115342 598172
rect 115398 598116 115494 598172
rect 114874 598048 115494 598116
rect 114874 597992 114970 598048
rect 115026 597992 115094 598048
rect 115150 597992 115218 598048
rect 115274 597992 115342 598048
rect 115398 597992 115494 598048
rect 114874 597924 115494 597992
rect 114874 597868 114970 597924
rect 115026 597868 115094 597924
rect 115150 597868 115218 597924
rect 115274 597868 115342 597924
rect 115398 597868 115494 597924
rect 114874 597800 115494 597868
rect 114874 597744 114970 597800
rect 115026 597744 115094 597800
rect 115150 597744 115218 597800
rect 115274 597744 115342 597800
rect 115398 597744 115494 597800
rect 114874 586350 115494 597744
rect 114874 586294 114970 586350
rect 115026 586294 115094 586350
rect 115150 586294 115218 586350
rect 115274 586294 115342 586350
rect 115398 586294 115494 586350
rect 114874 586226 115494 586294
rect 114874 586170 114970 586226
rect 115026 586170 115094 586226
rect 115150 586170 115218 586226
rect 115274 586170 115342 586226
rect 115398 586170 115494 586226
rect 114874 586102 115494 586170
rect 114874 586046 114970 586102
rect 115026 586046 115094 586102
rect 115150 586046 115218 586102
rect 115274 586046 115342 586102
rect 115398 586046 115494 586102
rect 114874 585978 115494 586046
rect 114874 585922 114970 585978
rect 115026 585922 115094 585978
rect 115150 585922 115218 585978
rect 115274 585922 115342 585978
rect 115398 585922 115494 585978
rect 114874 568350 115494 585922
rect 114874 568294 114970 568350
rect 115026 568294 115094 568350
rect 115150 568294 115218 568350
rect 115274 568294 115342 568350
rect 115398 568294 115494 568350
rect 114874 568226 115494 568294
rect 114874 568170 114970 568226
rect 115026 568170 115094 568226
rect 115150 568170 115218 568226
rect 115274 568170 115342 568226
rect 115398 568170 115494 568226
rect 114874 568102 115494 568170
rect 114874 568046 114970 568102
rect 115026 568046 115094 568102
rect 115150 568046 115218 568102
rect 115274 568046 115342 568102
rect 115398 568046 115494 568102
rect 114874 567978 115494 568046
rect 114874 567922 114970 567978
rect 115026 567922 115094 567978
rect 115150 567922 115218 567978
rect 115274 567922 115342 567978
rect 115398 567922 115494 567978
rect 114874 550350 115494 567922
rect 114874 550294 114970 550350
rect 115026 550294 115094 550350
rect 115150 550294 115218 550350
rect 115274 550294 115342 550350
rect 115398 550294 115494 550350
rect 114874 550226 115494 550294
rect 114874 550170 114970 550226
rect 115026 550170 115094 550226
rect 115150 550170 115218 550226
rect 115274 550170 115342 550226
rect 115398 550170 115494 550226
rect 114874 550102 115494 550170
rect 114874 550046 114970 550102
rect 115026 550046 115094 550102
rect 115150 550046 115218 550102
rect 115274 550046 115342 550102
rect 115398 550046 115494 550102
rect 114874 549978 115494 550046
rect 114874 549922 114970 549978
rect 115026 549922 115094 549978
rect 115150 549922 115218 549978
rect 115274 549922 115342 549978
rect 115398 549922 115494 549978
rect 114874 532350 115494 549922
rect 114874 532294 114970 532350
rect 115026 532294 115094 532350
rect 115150 532294 115218 532350
rect 115274 532294 115342 532350
rect 115398 532294 115494 532350
rect 114874 532226 115494 532294
rect 114874 532170 114970 532226
rect 115026 532170 115094 532226
rect 115150 532170 115218 532226
rect 115274 532170 115342 532226
rect 115398 532170 115494 532226
rect 114874 532102 115494 532170
rect 114874 532046 114970 532102
rect 115026 532046 115094 532102
rect 115150 532046 115218 532102
rect 115274 532046 115342 532102
rect 115398 532046 115494 532102
rect 114874 531978 115494 532046
rect 114874 531922 114970 531978
rect 115026 531922 115094 531978
rect 115150 531922 115218 531978
rect 115274 531922 115342 531978
rect 115398 531922 115494 531978
rect 114874 514350 115494 531922
rect 114874 514294 114970 514350
rect 115026 514294 115094 514350
rect 115150 514294 115218 514350
rect 115274 514294 115342 514350
rect 115398 514294 115494 514350
rect 114874 514226 115494 514294
rect 114874 514170 114970 514226
rect 115026 514170 115094 514226
rect 115150 514170 115218 514226
rect 115274 514170 115342 514226
rect 115398 514170 115494 514226
rect 114874 514102 115494 514170
rect 114874 514046 114970 514102
rect 115026 514046 115094 514102
rect 115150 514046 115218 514102
rect 115274 514046 115342 514102
rect 115398 514046 115494 514102
rect 114874 513978 115494 514046
rect 114874 513922 114970 513978
rect 115026 513922 115094 513978
rect 115150 513922 115218 513978
rect 115274 513922 115342 513978
rect 115398 513922 115494 513978
rect 114874 496350 115494 513922
rect 114874 496294 114970 496350
rect 115026 496294 115094 496350
rect 115150 496294 115218 496350
rect 115274 496294 115342 496350
rect 115398 496294 115494 496350
rect 114874 496226 115494 496294
rect 114874 496170 114970 496226
rect 115026 496170 115094 496226
rect 115150 496170 115218 496226
rect 115274 496170 115342 496226
rect 115398 496170 115494 496226
rect 114874 496102 115494 496170
rect 114874 496046 114970 496102
rect 115026 496046 115094 496102
rect 115150 496046 115218 496102
rect 115274 496046 115342 496102
rect 115398 496046 115494 496102
rect 114874 495978 115494 496046
rect 114874 495922 114970 495978
rect 115026 495922 115094 495978
rect 115150 495922 115218 495978
rect 115274 495922 115342 495978
rect 115398 495922 115494 495978
rect 114874 478350 115494 495922
rect 114874 478294 114970 478350
rect 115026 478294 115094 478350
rect 115150 478294 115218 478350
rect 115274 478294 115342 478350
rect 115398 478294 115494 478350
rect 114874 478226 115494 478294
rect 114874 478170 114970 478226
rect 115026 478170 115094 478226
rect 115150 478170 115218 478226
rect 115274 478170 115342 478226
rect 115398 478170 115494 478226
rect 114874 478102 115494 478170
rect 114874 478046 114970 478102
rect 115026 478046 115094 478102
rect 115150 478046 115218 478102
rect 115274 478046 115342 478102
rect 115398 478046 115494 478102
rect 114874 477978 115494 478046
rect 114874 477922 114970 477978
rect 115026 477922 115094 477978
rect 115150 477922 115218 477978
rect 115274 477922 115342 477978
rect 115398 477922 115494 477978
rect 114874 460350 115494 477922
rect 114874 460294 114970 460350
rect 115026 460294 115094 460350
rect 115150 460294 115218 460350
rect 115274 460294 115342 460350
rect 115398 460294 115494 460350
rect 114874 460226 115494 460294
rect 114874 460170 114970 460226
rect 115026 460170 115094 460226
rect 115150 460170 115218 460226
rect 115274 460170 115342 460226
rect 115398 460170 115494 460226
rect 114874 460102 115494 460170
rect 114874 460046 114970 460102
rect 115026 460046 115094 460102
rect 115150 460046 115218 460102
rect 115274 460046 115342 460102
rect 115398 460046 115494 460102
rect 114874 459978 115494 460046
rect 114874 459922 114970 459978
rect 115026 459922 115094 459978
rect 115150 459922 115218 459978
rect 115274 459922 115342 459978
rect 115398 459922 115494 459978
rect 114874 458342 115494 459922
rect 129154 597212 129774 598268
rect 129154 597156 129250 597212
rect 129306 597156 129374 597212
rect 129430 597156 129498 597212
rect 129554 597156 129622 597212
rect 129678 597156 129774 597212
rect 129154 597088 129774 597156
rect 129154 597032 129250 597088
rect 129306 597032 129374 597088
rect 129430 597032 129498 597088
rect 129554 597032 129622 597088
rect 129678 597032 129774 597088
rect 129154 596964 129774 597032
rect 129154 596908 129250 596964
rect 129306 596908 129374 596964
rect 129430 596908 129498 596964
rect 129554 596908 129622 596964
rect 129678 596908 129774 596964
rect 129154 596840 129774 596908
rect 129154 596784 129250 596840
rect 129306 596784 129374 596840
rect 129430 596784 129498 596840
rect 129554 596784 129622 596840
rect 129678 596784 129774 596840
rect 129154 580350 129774 596784
rect 129154 580294 129250 580350
rect 129306 580294 129374 580350
rect 129430 580294 129498 580350
rect 129554 580294 129622 580350
rect 129678 580294 129774 580350
rect 129154 580226 129774 580294
rect 129154 580170 129250 580226
rect 129306 580170 129374 580226
rect 129430 580170 129498 580226
rect 129554 580170 129622 580226
rect 129678 580170 129774 580226
rect 129154 580102 129774 580170
rect 129154 580046 129250 580102
rect 129306 580046 129374 580102
rect 129430 580046 129498 580102
rect 129554 580046 129622 580102
rect 129678 580046 129774 580102
rect 129154 579978 129774 580046
rect 129154 579922 129250 579978
rect 129306 579922 129374 579978
rect 129430 579922 129498 579978
rect 129554 579922 129622 579978
rect 129678 579922 129774 579978
rect 129154 562350 129774 579922
rect 129154 562294 129250 562350
rect 129306 562294 129374 562350
rect 129430 562294 129498 562350
rect 129554 562294 129622 562350
rect 129678 562294 129774 562350
rect 129154 562226 129774 562294
rect 129154 562170 129250 562226
rect 129306 562170 129374 562226
rect 129430 562170 129498 562226
rect 129554 562170 129622 562226
rect 129678 562170 129774 562226
rect 129154 562102 129774 562170
rect 129154 562046 129250 562102
rect 129306 562046 129374 562102
rect 129430 562046 129498 562102
rect 129554 562046 129622 562102
rect 129678 562046 129774 562102
rect 129154 561978 129774 562046
rect 129154 561922 129250 561978
rect 129306 561922 129374 561978
rect 129430 561922 129498 561978
rect 129554 561922 129622 561978
rect 129678 561922 129774 561978
rect 129154 544350 129774 561922
rect 129154 544294 129250 544350
rect 129306 544294 129374 544350
rect 129430 544294 129498 544350
rect 129554 544294 129622 544350
rect 129678 544294 129774 544350
rect 129154 544226 129774 544294
rect 129154 544170 129250 544226
rect 129306 544170 129374 544226
rect 129430 544170 129498 544226
rect 129554 544170 129622 544226
rect 129678 544170 129774 544226
rect 129154 544102 129774 544170
rect 129154 544046 129250 544102
rect 129306 544046 129374 544102
rect 129430 544046 129498 544102
rect 129554 544046 129622 544102
rect 129678 544046 129774 544102
rect 129154 543978 129774 544046
rect 129154 543922 129250 543978
rect 129306 543922 129374 543978
rect 129430 543922 129498 543978
rect 129554 543922 129622 543978
rect 129678 543922 129774 543978
rect 129154 526350 129774 543922
rect 129154 526294 129250 526350
rect 129306 526294 129374 526350
rect 129430 526294 129498 526350
rect 129554 526294 129622 526350
rect 129678 526294 129774 526350
rect 129154 526226 129774 526294
rect 129154 526170 129250 526226
rect 129306 526170 129374 526226
rect 129430 526170 129498 526226
rect 129554 526170 129622 526226
rect 129678 526170 129774 526226
rect 129154 526102 129774 526170
rect 129154 526046 129250 526102
rect 129306 526046 129374 526102
rect 129430 526046 129498 526102
rect 129554 526046 129622 526102
rect 129678 526046 129774 526102
rect 129154 525978 129774 526046
rect 129154 525922 129250 525978
rect 129306 525922 129374 525978
rect 129430 525922 129498 525978
rect 129554 525922 129622 525978
rect 129678 525922 129774 525978
rect 129154 508350 129774 525922
rect 129154 508294 129250 508350
rect 129306 508294 129374 508350
rect 129430 508294 129498 508350
rect 129554 508294 129622 508350
rect 129678 508294 129774 508350
rect 129154 508226 129774 508294
rect 129154 508170 129250 508226
rect 129306 508170 129374 508226
rect 129430 508170 129498 508226
rect 129554 508170 129622 508226
rect 129678 508170 129774 508226
rect 129154 508102 129774 508170
rect 129154 508046 129250 508102
rect 129306 508046 129374 508102
rect 129430 508046 129498 508102
rect 129554 508046 129622 508102
rect 129678 508046 129774 508102
rect 129154 507978 129774 508046
rect 129154 507922 129250 507978
rect 129306 507922 129374 507978
rect 129430 507922 129498 507978
rect 129554 507922 129622 507978
rect 129678 507922 129774 507978
rect 129154 490350 129774 507922
rect 129154 490294 129250 490350
rect 129306 490294 129374 490350
rect 129430 490294 129498 490350
rect 129554 490294 129622 490350
rect 129678 490294 129774 490350
rect 129154 490226 129774 490294
rect 129154 490170 129250 490226
rect 129306 490170 129374 490226
rect 129430 490170 129498 490226
rect 129554 490170 129622 490226
rect 129678 490170 129774 490226
rect 129154 490102 129774 490170
rect 129154 490046 129250 490102
rect 129306 490046 129374 490102
rect 129430 490046 129498 490102
rect 129554 490046 129622 490102
rect 129678 490046 129774 490102
rect 129154 489978 129774 490046
rect 129154 489922 129250 489978
rect 129306 489922 129374 489978
rect 129430 489922 129498 489978
rect 129554 489922 129622 489978
rect 129678 489922 129774 489978
rect 129154 472350 129774 489922
rect 129154 472294 129250 472350
rect 129306 472294 129374 472350
rect 129430 472294 129498 472350
rect 129554 472294 129622 472350
rect 129678 472294 129774 472350
rect 129154 472226 129774 472294
rect 129154 472170 129250 472226
rect 129306 472170 129374 472226
rect 129430 472170 129498 472226
rect 129554 472170 129622 472226
rect 129678 472170 129774 472226
rect 129154 472102 129774 472170
rect 129154 472046 129250 472102
rect 129306 472046 129374 472102
rect 129430 472046 129498 472102
rect 129554 472046 129622 472102
rect 129678 472046 129774 472102
rect 129154 471978 129774 472046
rect 129154 471922 129250 471978
rect 129306 471922 129374 471978
rect 129430 471922 129498 471978
rect 129554 471922 129622 471978
rect 129678 471922 129774 471978
rect 129154 458342 129774 471922
rect 132874 598172 133494 598268
rect 132874 598116 132970 598172
rect 133026 598116 133094 598172
rect 133150 598116 133218 598172
rect 133274 598116 133342 598172
rect 133398 598116 133494 598172
rect 132874 598048 133494 598116
rect 132874 597992 132970 598048
rect 133026 597992 133094 598048
rect 133150 597992 133218 598048
rect 133274 597992 133342 598048
rect 133398 597992 133494 598048
rect 132874 597924 133494 597992
rect 132874 597868 132970 597924
rect 133026 597868 133094 597924
rect 133150 597868 133218 597924
rect 133274 597868 133342 597924
rect 133398 597868 133494 597924
rect 132874 597800 133494 597868
rect 132874 597744 132970 597800
rect 133026 597744 133094 597800
rect 133150 597744 133218 597800
rect 133274 597744 133342 597800
rect 133398 597744 133494 597800
rect 132874 586350 133494 597744
rect 132874 586294 132970 586350
rect 133026 586294 133094 586350
rect 133150 586294 133218 586350
rect 133274 586294 133342 586350
rect 133398 586294 133494 586350
rect 132874 586226 133494 586294
rect 132874 586170 132970 586226
rect 133026 586170 133094 586226
rect 133150 586170 133218 586226
rect 133274 586170 133342 586226
rect 133398 586170 133494 586226
rect 132874 586102 133494 586170
rect 132874 586046 132970 586102
rect 133026 586046 133094 586102
rect 133150 586046 133218 586102
rect 133274 586046 133342 586102
rect 133398 586046 133494 586102
rect 132874 585978 133494 586046
rect 132874 585922 132970 585978
rect 133026 585922 133094 585978
rect 133150 585922 133218 585978
rect 133274 585922 133342 585978
rect 133398 585922 133494 585978
rect 132874 568350 133494 585922
rect 132874 568294 132970 568350
rect 133026 568294 133094 568350
rect 133150 568294 133218 568350
rect 133274 568294 133342 568350
rect 133398 568294 133494 568350
rect 132874 568226 133494 568294
rect 132874 568170 132970 568226
rect 133026 568170 133094 568226
rect 133150 568170 133218 568226
rect 133274 568170 133342 568226
rect 133398 568170 133494 568226
rect 132874 568102 133494 568170
rect 132874 568046 132970 568102
rect 133026 568046 133094 568102
rect 133150 568046 133218 568102
rect 133274 568046 133342 568102
rect 133398 568046 133494 568102
rect 132874 567978 133494 568046
rect 132874 567922 132970 567978
rect 133026 567922 133094 567978
rect 133150 567922 133218 567978
rect 133274 567922 133342 567978
rect 133398 567922 133494 567978
rect 132874 550350 133494 567922
rect 132874 550294 132970 550350
rect 133026 550294 133094 550350
rect 133150 550294 133218 550350
rect 133274 550294 133342 550350
rect 133398 550294 133494 550350
rect 132874 550226 133494 550294
rect 132874 550170 132970 550226
rect 133026 550170 133094 550226
rect 133150 550170 133218 550226
rect 133274 550170 133342 550226
rect 133398 550170 133494 550226
rect 132874 550102 133494 550170
rect 132874 550046 132970 550102
rect 133026 550046 133094 550102
rect 133150 550046 133218 550102
rect 133274 550046 133342 550102
rect 133398 550046 133494 550102
rect 132874 549978 133494 550046
rect 132874 549922 132970 549978
rect 133026 549922 133094 549978
rect 133150 549922 133218 549978
rect 133274 549922 133342 549978
rect 133398 549922 133494 549978
rect 132874 532350 133494 549922
rect 132874 532294 132970 532350
rect 133026 532294 133094 532350
rect 133150 532294 133218 532350
rect 133274 532294 133342 532350
rect 133398 532294 133494 532350
rect 132874 532226 133494 532294
rect 132874 532170 132970 532226
rect 133026 532170 133094 532226
rect 133150 532170 133218 532226
rect 133274 532170 133342 532226
rect 133398 532170 133494 532226
rect 132874 532102 133494 532170
rect 132874 532046 132970 532102
rect 133026 532046 133094 532102
rect 133150 532046 133218 532102
rect 133274 532046 133342 532102
rect 133398 532046 133494 532102
rect 132874 531978 133494 532046
rect 132874 531922 132970 531978
rect 133026 531922 133094 531978
rect 133150 531922 133218 531978
rect 133274 531922 133342 531978
rect 133398 531922 133494 531978
rect 132874 514350 133494 531922
rect 132874 514294 132970 514350
rect 133026 514294 133094 514350
rect 133150 514294 133218 514350
rect 133274 514294 133342 514350
rect 133398 514294 133494 514350
rect 132874 514226 133494 514294
rect 132874 514170 132970 514226
rect 133026 514170 133094 514226
rect 133150 514170 133218 514226
rect 133274 514170 133342 514226
rect 133398 514170 133494 514226
rect 132874 514102 133494 514170
rect 132874 514046 132970 514102
rect 133026 514046 133094 514102
rect 133150 514046 133218 514102
rect 133274 514046 133342 514102
rect 133398 514046 133494 514102
rect 132874 513978 133494 514046
rect 132874 513922 132970 513978
rect 133026 513922 133094 513978
rect 133150 513922 133218 513978
rect 133274 513922 133342 513978
rect 133398 513922 133494 513978
rect 132874 496350 133494 513922
rect 132874 496294 132970 496350
rect 133026 496294 133094 496350
rect 133150 496294 133218 496350
rect 133274 496294 133342 496350
rect 133398 496294 133494 496350
rect 132874 496226 133494 496294
rect 132874 496170 132970 496226
rect 133026 496170 133094 496226
rect 133150 496170 133218 496226
rect 133274 496170 133342 496226
rect 133398 496170 133494 496226
rect 132874 496102 133494 496170
rect 132874 496046 132970 496102
rect 133026 496046 133094 496102
rect 133150 496046 133218 496102
rect 133274 496046 133342 496102
rect 133398 496046 133494 496102
rect 132874 495978 133494 496046
rect 132874 495922 132970 495978
rect 133026 495922 133094 495978
rect 133150 495922 133218 495978
rect 133274 495922 133342 495978
rect 133398 495922 133494 495978
rect 132874 478350 133494 495922
rect 132874 478294 132970 478350
rect 133026 478294 133094 478350
rect 133150 478294 133218 478350
rect 133274 478294 133342 478350
rect 133398 478294 133494 478350
rect 132874 478226 133494 478294
rect 132874 478170 132970 478226
rect 133026 478170 133094 478226
rect 133150 478170 133218 478226
rect 133274 478170 133342 478226
rect 133398 478170 133494 478226
rect 132874 478102 133494 478170
rect 132874 478046 132970 478102
rect 133026 478046 133094 478102
rect 133150 478046 133218 478102
rect 133274 478046 133342 478102
rect 133398 478046 133494 478102
rect 132874 477978 133494 478046
rect 132874 477922 132970 477978
rect 133026 477922 133094 477978
rect 133150 477922 133218 477978
rect 133274 477922 133342 477978
rect 133398 477922 133494 477978
rect 132874 460350 133494 477922
rect 132874 460294 132970 460350
rect 133026 460294 133094 460350
rect 133150 460294 133218 460350
rect 133274 460294 133342 460350
rect 133398 460294 133494 460350
rect 132874 460226 133494 460294
rect 132874 460170 132970 460226
rect 133026 460170 133094 460226
rect 133150 460170 133218 460226
rect 133274 460170 133342 460226
rect 133398 460170 133494 460226
rect 132874 460102 133494 460170
rect 132874 460046 132970 460102
rect 133026 460046 133094 460102
rect 133150 460046 133218 460102
rect 133274 460046 133342 460102
rect 133398 460046 133494 460102
rect 132874 459978 133494 460046
rect 132874 459922 132970 459978
rect 133026 459922 133094 459978
rect 133150 459922 133218 459978
rect 133274 459922 133342 459978
rect 133398 459922 133494 459978
rect 132874 458342 133494 459922
rect 147154 597212 147774 598268
rect 147154 597156 147250 597212
rect 147306 597156 147374 597212
rect 147430 597156 147498 597212
rect 147554 597156 147622 597212
rect 147678 597156 147774 597212
rect 147154 597088 147774 597156
rect 147154 597032 147250 597088
rect 147306 597032 147374 597088
rect 147430 597032 147498 597088
rect 147554 597032 147622 597088
rect 147678 597032 147774 597088
rect 147154 596964 147774 597032
rect 147154 596908 147250 596964
rect 147306 596908 147374 596964
rect 147430 596908 147498 596964
rect 147554 596908 147622 596964
rect 147678 596908 147774 596964
rect 147154 596840 147774 596908
rect 147154 596784 147250 596840
rect 147306 596784 147374 596840
rect 147430 596784 147498 596840
rect 147554 596784 147622 596840
rect 147678 596784 147774 596840
rect 147154 580350 147774 596784
rect 147154 580294 147250 580350
rect 147306 580294 147374 580350
rect 147430 580294 147498 580350
rect 147554 580294 147622 580350
rect 147678 580294 147774 580350
rect 147154 580226 147774 580294
rect 147154 580170 147250 580226
rect 147306 580170 147374 580226
rect 147430 580170 147498 580226
rect 147554 580170 147622 580226
rect 147678 580170 147774 580226
rect 147154 580102 147774 580170
rect 147154 580046 147250 580102
rect 147306 580046 147374 580102
rect 147430 580046 147498 580102
rect 147554 580046 147622 580102
rect 147678 580046 147774 580102
rect 147154 579978 147774 580046
rect 147154 579922 147250 579978
rect 147306 579922 147374 579978
rect 147430 579922 147498 579978
rect 147554 579922 147622 579978
rect 147678 579922 147774 579978
rect 147154 562350 147774 579922
rect 147154 562294 147250 562350
rect 147306 562294 147374 562350
rect 147430 562294 147498 562350
rect 147554 562294 147622 562350
rect 147678 562294 147774 562350
rect 147154 562226 147774 562294
rect 147154 562170 147250 562226
rect 147306 562170 147374 562226
rect 147430 562170 147498 562226
rect 147554 562170 147622 562226
rect 147678 562170 147774 562226
rect 147154 562102 147774 562170
rect 147154 562046 147250 562102
rect 147306 562046 147374 562102
rect 147430 562046 147498 562102
rect 147554 562046 147622 562102
rect 147678 562046 147774 562102
rect 147154 561978 147774 562046
rect 147154 561922 147250 561978
rect 147306 561922 147374 561978
rect 147430 561922 147498 561978
rect 147554 561922 147622 561978
rect 147678 561922 147774 561978
rect 147154 544350 147774 561922
rect 147154 544294 147250 544350
rect 147306 544294 147374 544350
rect 147430 544294 147498 544350
rect 147554 544294 147622 544350
rect 147678 544294 147774 544350
rect 147154 544226 147774 544294
rect 147154 544170 147250 544226
rect 147306 544170 147374 544226
rect 147430 544170 147498 544226
rect 147554 544170 147622 544226
rect 147678 544170 147774 544226
rect 147154 544102 147774 544170
rect 147154 544046 147250 544102
rect 147306 544046 147374 544102
rect 147430 544046 147498 544102
rect 147554 544046 147622 544102
rect 147678 544046 147774 544102
rect 147154 543978 147774 544046
rect 147154 543922 147250 543978
rect 147306 543922 147374 543978
rect 147430 543922 147498 543978
rect 147554 543922 147622 543978
rect 147678 543922 147774 543978
rect 147154 526350 147774 543922
rect 147154 526294 147250 526350
rect 147306 526294 147374 526350
rect 147430 526294 147498 526350
rect 147554 526294 147622 526350
rect 147678 526294 147774 526350
rect 147154 526226 147774 526294
rect 147154 526170 147250 526226
rect 147306 526170 147374 526226
rect 147430 526170 147498 526226
rect 147554 526170 147622 526226
rect 147678 526170 147774 526226
rect 147154 526102 147774 526170
rect 147154 526046 147250 526102
rect 147306 526046 147374 526102
rect 147430 526046 147498 526102
rect 147554 526046 147622 526102
rect 147678 526046 147774 526102
rect 147154 525978 147774 526046
rect 147154 525922 147250 525978
rect 147306 525922 147374 525978
rect 147430 525922 147498 525978
rect 147554 525922 147622 525978
rect 147678 525922 147774 525978
rect 147154 508350 147774 525922
rect 147154 508294 147250 508350
rect 147306 508294 147374 508350
rect 147430 508294 147498 508350
rect 147554 508294 147622 508350
rect 147678 508294 147774 508350
rect 147154 508226 147774 508294
rect 147154 508170 147250 508226
rect 147306 508170 147374 508226
rect 147430 508170 147498 508226
rect 147554 508170 147622 508226
rect 147678 508170 147774 508226
rect 147154 508102 147774 508170
rect 147154 508046 147250 508102
rect 147306 508046 147374 508102
rect 147430 508046 147498 508102
rect 147554 508046 147622 508102
rect 147678 508046 147774 508102
rect 147154 507978 147774 508046
rect 147154 507922 147250 507978
rect 147306 507922 147374 507978
rect 147430 507922 147498 507978
rect 147554 507922 147622 507978
rect 147678 507922 147774 507978
rect 147154 490350 147774 507922
rect 147154 490294 147250 490350
rect 147306 490294 147374 490350
rect 147430 490294 147498 490350
rect 147554 490294 147622 490350
rect 147678 490294 147774 490350
rect 147154 490226 147774 490294
rect 147154 490170 147250 490226
rect 147306 490170 147374 490226
rect 147430 490170 147498 490226
rect 147554 490170 147622 490226
rect 147678 490170 147774 490226
rect 147154 490102 147774 490170
rect 147154 490046 147250 490102
rect 147306 490046 147374 490102
rect 147430 490046 147498 490102
rect 147554 490046 147622 490102
rect 147678 490046 147774 490102
rect 147154 489978 147774 490046
rect 147154 489922 147250 489978
rect 147306 489922 147374 489978
rect 147430 489922 147498 489978
rect 147554 489922 147622 489978
rect 147678 489922 147774 489978
rect 147154 472350 147774 489922
rect 147154 472294 147250 472350
rect 147306 472294 147374 472350
rect 147430 472294 147498 472350
rect 147554 472294 147622 472350
rect 147678 472294 147774 472350
rect 147154 472226 147774 472294
rect 147154 472170 147250 472226
rect 147306 472170 147374 472226
rect 147430 472170 147498 472226
rect 147554 472170 147622 472226
rect 147678 472170 147774 472226
rect 147154 472102 147774 472170
rect 147154 472046 147250 472102
rect 147306 472046 147374 472102
rect 147430 472046 147498 472102
rect 147554 472046 147622 472102
rect 147678 472046 147774 472102
rect 147154 471978 147774 472046
rect 147154 471922 147250 471978
rect 147306 471922 147374 471978
rect 147430 471922 147498 471978
rect 147554 471922 147622 471978
rect 147678 471922 147774 471978
rect 147154 458342 147774 471922
rect 150874 598172 151494 598268
rect 150874 598116 150970 598172
rect 151026 598116 151094 598172
rect 151150 598116 151218 598172
rect 151274 598116 151342 598172
rect 151398 598116 151494 598172
rect 150874 598048 151494 598116
rect 150874 597992 150970 598048
rect 151026 597992 151094 598048
rect 151150 597992 151218 598048
rect 151274 597992 151342 598048
rect 151398 597992 151494 598048
rect 150874 597924 151494 597992
rect 150874 597868 150970 597924
rect 151026 597868 151094 597924
rect 151150 597868 151218 597924
rect 151274 597868 151342 597924
rect 151398 597868 151494 597924
rect 150874 597800 151494 597868
rect 150874 597744 150970 597800
rect 151026 597744 151094 597800
rect 151150 597744 151218 597800
rect 151274 597744 151342 597800
rect 151398 597744 151494 597800
rect 150874 586350 151494 597744
rect 150874 586294 150970 586350
rect 151026 586294 151094 586350
rect 151150 586294 151218 586350
rect 151274 586294 151342 586350
rect 151398 586294 151494 586350
rect 150874 586226 151494 586294
rect 150874 586170 150970 586226
rect 151026 586170 151094 586226
rect 151150 586170 151218 586226
rect 151274 586170 151342 586226
rect 151398 586170 151494 586226
rect 150874 586102 151494 586170
rect 150874 586046 150970 586102
rect 151026 586046 151094 586102
rect 151150 586046 151218 586102
rect 151274 586046 151342 586102
rect 151398 586046 151494 586102
rect 150874 585978 151494 586046
rect 150874 585922 150970 585978
rect 151026 585922 151094 585978
rect 151150 585922 151218 585978
rect 151274 585922 151342 585978
rect 151398 585922 151494 585978
rect 150874 568350 151494 585922
rect 150874 568294 150970 568350
rect 151026 568294 151094 568350
rect 151150 568294 151218 568350
rect 151274 568294 151342 568350
rect 151398 568294 151494 568350
rect 150874 568226 151494 568294
rect 150874 568170 150970 568226
rect 151026 568170 151094 568226
rect 151150 568170 151218 568226
rect 151274 568170 151342 568226
rect 151398 568170 151494 568226
rect 150874 568102 151494 568170
rect 150874 568046 150970 568102
rect 151026 568046 151094 568102
rect 151150 568046 151218 568102
rect 151274 568046 151342 568102
rect 151398 568046 151494 568102
rect 150874 567978 151494 568046
rect 150874 567922 150970 567978
rect 151026 567922 151094 567978
rect 151150 567922 151218 567978
rect 151274 567922 151342 567978
rect 151398 567922 151494 567978
rect 150874 550350 151494 567922
rect 150874 550294 150970 550350
rect 151026 550294 151094 550350
rect 151150 550294 151218 550350
rect 151274 550294 151342 550350
rect 151398 550294 151494 550350
rect 150874 550226 151494 550294
rect 150874 550170 150970 550226
rect 151026 550170 151094 550226
rect 151150 550170 151218 550226
rect 151274 550170 151342 550226
rect 151398 550170 151494 550226
rect 150874 550102 151494 550170
rect 150874 550046 150970 550102
rect 151026 550046 151094 550102
rect 151150 550046 151218 550102
rect 151274 550046 151342 550102
rect 151398 550046 151494 550102
rect 150874 549978 151494 550046
rect 150874 549922 150970 549978
rect 151026 549922 151094 549978
rect 151150 549922 151218 549978
rect 151274 549922 151342 549978
rect 151398 549922 151494 549978
rect 150874 532350 151494 549922
rect 150874 532294 150970 532350
rect 151026 532294 151094 532350
rect 151150 532294 151218 532350
rect 151274 532294 151342 532350
rect 151398 532294 151494 532350
rect 150874 532226 151494 532294
rect 150874 532170 150970 532226
rect 151026 532170 151094 532226
rect 151150 532170 151218 532226
rect 151274 532170 151342 532226
rect 151398 532170 151494 532226
rect 150874 532102 151494 532170
rect 150874 532046 150970 532102
rect 151026 532046 151094 532102
rect 151150 532046 151218 532102
rect 151274 532046 151342 532102
rect 151398 532046 151494 532102
rect 150874 531978 151494 532046
rect 150874 531922 150970 531978
rect 151026 531922 151094 531978
rect 151150 531922 151218 531978
rect 151274 531922 151342 531978
rect 151398 531922 151494 531978
rect 150874 514350 151494 531922
rect 150874 514294 150970 514350
rect 151026 514294 151094 514350
rect 151150 514294 151218 514350
rect 151274 514294 151342 514350
rect 151398 514294 151494 514350
rect 150874 514226 151494 514294
rect 150874 514170 150970 514226
rect 151026 514170 151094 514226
rect 151150 514170 151218 514226
rect 151274 514170 151342 514226
rect 151398 514170 151494 514226
rect 150874 514102 151494 514170
rect 150874 514046 150970 514102
rect 151026 514046 151094 514102
rect 151150 514046 151218 514102
rect 151274 514046 151342 514102
rect 151398 514046 151494 514102
rect 150874 513978 151494 514046
rect 150874 513922 150970 513978
rect 151026 513922 151094 513978
rect 151150 513922 151218 513978
rect 151274 513922 151342 513978
rect 151398 513922 151494 513978
rect 150874 496350 151494 513922
rect 150874 496294 150970 496350
rect 151026 496294 151094 496350
rect 151150 496294 151218 496350
rect 151274 496294 151342 496350
rect 151398 496294 151494 496350
rect 150874 496226 151494 496294
rect 150874 496170 150970 496226
rect 151026 496170 151094 496226
rect 151150 496170 151218 496226
rect 151274 496170 151342 496226
rect 151398 496170 151494 496226
rect 150874 496102 151494 496170
rect 150874 496046 150970 496102
rect 151026 496046 151094 496102
rect 151150 496046 151218 496102
rect 151274 496046 151342 496102
rect 151398 496046 151494 496102
rect 150874 495978 151494 496046
rect 150874 495922 150970 495978
rect 151026 495922 151094 495978
rect 151150 495922 151218 495978
rect 151274 495922 151342 495978
rect 151398 495922 151494 495978
rect 150874 478350 151494 495922
rect 150874 478294 150970 478350
rect 151026 478294 151094 478350
rect 151150 478294 151218 478350
rect 151274 478294 151342 478350
rect 151398 478294 151494 478350
rect 150874 478226 151494 478294
rect 150874 478170 150970 478226
rect 151026 478170 151094 478226
rect 151150 478170 151218 478226
rect 151274 478170 151342 478226
rect 151398 478170 151494 478226
rect 150874 478102 151494 478170
rect 150874 478046 150970 478102
rect 151026 478046 151094 478102
rect 151150 478046 151218 478102
rect 151274 478046 151342 478102
rect 151398 478046 151494 478102
rect 150874 477978 151494 478046
rect 150874 477922 150970 477978
rect 151026 477922 151094 477978
rect 151150 477922 151218 477978
rect 151274 477922 151342 477978
rect 151398 477922 151494 477978
rect 150874 460350 151494 477922
rect 150874 460294 150970 460350
rect 151026 460294 151094 460350
rect 151150 460294 151218 460350
rect 151274 460294 151342 460350
rect 151398 460294 151494 460350
rect 150874 460226 151494 460294
rect 150874 460170 150970 460226
rect 151026 460170 151094 460226
rect 151150 460170 151218 460226
rect 151274 460170 151342 460226
rect 151398 460170 151494 460226
rect 150874 460102 151494 460170
rect 150874 460046 150970 460102
rect 151026 460046 151094 460102
rect 151150 460046 151218 460102
rect 151274 460046 151342 460102
rect 151398 460046 151494 460102
rect 150874 459978 151494 460046
rect 150874 459922 150970 459978
rect 151026 459922 151094 459978
rect 151150 459922 151218 459978
rect 151274 459922 151342 459978
rect 151398 459922 151494 459978
rect 150874 458342 151494 459922
rect 165154 597212 165774 598268
rect 165154 597156 165250 597212
rect 165306 597156 165374 597212
rect 165430 597156 165498 597212
rect 165554 597156 165622 597212
rect 165678 597156 165774 597212
rect 165154 597088 165774 597156
rect 165154 597032 165250 597088
rect 165306 597032 165374 597088
rect 165430 597032 165498 597088
rect 165554 597032 165622 597088
rect 165678 597032 165774 597088
rect 165154 596964 165774 597032
rect 165154 596908 165250 596964
rect 165306 596908 165374 596964
rect 165430 596908 165498 596964
rect 165554 596908 165622 596964
rect 165678 596908 165774 596964
rect 165154 596840 165774 596908
rect 165154 596784 165250 596840
rect 165306 596784 165374 596840
rect 165430 596784 165498 596840
rect 165554 596784 165622 596840
rect 165678 596784 165774 596840
rect 165154 580350 165774 596784
rect 165154 580294 165250 580350
rect 165306 580294 165374 580350
rect 165430 580294 165498 580350
rect 165554 580294 165622 580350
rect 165678 580294 165774 580350
rect 165154 580226 165774 580294
rect 165154 580170 165250 580226
rect 165306 580170 165374 580226
rect 165430 580170 165498 580226
rect 165554 580170 165622 580226
rect 165678 580170 165774 580226
rect 165154 580102 165774 580170
rect 165154 580046 165250 580102
rect 165306 580046 165374 580102
rect 165430 580046 165498 580102
rect 165554 580046 165622 580102
rect 165678 580046 165774 580102
rect 165154 579978 165774 580046
rect 165154 579922 165250 579978
rect 165306 579922 165374 579978
rect 165430 579922 165498 579978
rect 165554 579922 165622 579978
rect 165678 579922 165774 579978
rect 165154 562350 165774 579922
rect 165154 562294 165250 562350
rect 165306 562294 165374 562350
rect 165430 562294 165498 562350
rect 165554 562294 165622 562350
rect 165678 562294 165774 562350
rect 165154 562226 165774 562294
rect 165154 562170 165250 562226
rect 165306 562170 165374 562226
rect 165430 562170 165498 562226
rect 165554 562170 165622 562226
rect 165678 562170 165774 562226
rect 165154 562102 165774 562170
rect 165154 562046 165250 562102
rect 165306 562046 165374 562102
rect 165430 562046 165498 562102
rect 165554 562046 165622 562102
rect 165678 562046 165774 562102
rect 165154 561978 165774 562046
rect 165154 561922 165250 561978
rect 165306 561922 165374 561978
rect 165430 561922 165498 561978
rect 165554 561922 165622 561978
rect 165678 561922 165774 561978
rect 165154 544350 165774 561922
rect 165154 544294 165250 544350
rect 165306 544294 165374 544350
rect 165430 544294 165498 544350
rect 165554 544294 165622 544350
rect 165678 544294 165774 544350
rect 165154 544226 165774 544294
rect 165154 544170 165250 544226
rect 165306 544170 165374 544226
rect 165430 544170 165498 544226
rect 165554 544170 165622 544226
rect 165678 544170 165774 544226
rect 165154 544102 165774 544170
rect 165154 544046 165250 544102
rect 165306 544046 165374 544102
rect 165430 544046 165498 544102
rect 165554 544046 165622 544102
rect 165678 544046 165774 544102
rect 165154 543978 165774 544046
rect 165154 543922 165250 543978
rect 165306 543922 165374 543978
rect 165430 543922 165498 543978
rect 165554 543922 165622 543978
rect 165678 543922 165774 543978
rect 165154 526350 165774 543922
rect 165154 526294 165250 526350
rect 165306 526294 165374 526350
rect 165430 526294 165498 526350
rect 165554 526294 165622 526350
rect 165678 526294 165774 526350
rect 165154 526226 165774 526294
rect 165154 526170 165250 526226
rect 165306 526170 165374 526226
rect 165430 526170 165498 526226
rect 165554 526170 165622 526226
rect 165678 526170 165774 526226
rect 165154 526102 165774 526170
rect 165154 526046 165250 526102
rect 165306 526046 165374 526102
rect 165430 526046 165498 526102
rect 165554 526046 165622 526102
rect 165678 526046 165774 526102
rect 165154 525978 165774 526046
rect 165154 525922 165250 525978
rect 165306 525922 165374 525978
rect 165430 525922 165498 525978
rect 165554 525922 165622 525978
rect 165678 525922 165774 525978
rect 165154 508350 165774 525922
rect 165154 508294 165250 508350
rect 165306 508294 165374 508350
rect 165430 508294 165498 508350
rect 165554 508294 165622 508350
rect 165678 508294 165774 508350
rect 165154 508226 165774 508294
rect 165154 508170 165250 508226
rect 165306 508170 165374 508226
rect 165430 508170 165498 508226
rect 165554 508170 165622 508226
rect 165678 508170 165774 508226
rect 165154 508102 165774 508170
rect 165154 508046 165250 508102
rect 165306 508046 165374 508102
rect 165430 508046 165498 508102
rect 165554 508046 165622 508102
rect 165678 508046 165774 508102
rect 165154 507978 165774 508046
rect 165154 507922 165250 507978
rect 165306 507922 165374 507978
rect 165430 507922 165498 507978
rect 165554 507922 165622 507978
rect 165678 507922 165774 507978
rect 165154 490350 165774 507922
rect 165154 490294 165250 490350
rect 165306 490294 165374 490350
rect 165430 490294 165498 490350
rect 165554 490294 165622 490350
rect 165678 490294 165774 490350
rect 165154 490226 165774 490294
rect 165154 490170 165250 490226
rect 165306 490170 165374 490226
rect 165430 490170 165498 490226
rect 165554 490170 165622 490226
rect 165678 490170 165774 490226
rect 165154 490102 165774 490170
rect 165154 490046 165250 490102
rect 165306 490046 165374 490102
rect 165430 490046 165498 490102
rect 165554 490046 165622 490102
rect 165678 490046 165774 490102
rect 165154 489978 165774 490046
rect 165154 489922 165250 489978
rect 165306 489922 165374 489978
rect 165430 489922 165498 489978
rect 165554 489922 165622 489978
rect 165678 489922 165774 489978
rect 165154 472350 165774 489922
rect 165154 472294 165250 472350
rect 165306 472294 165374 472350
rect 165430 472294 165498 472350
rect 165554 472294 165622 472350
rect 165678 472294 165774 472350
rect 165154 472226 165774 472294
rect 165154 472170 165250 472226
rect 165306 472170 165374 472226
rect 165430 472170 165498 472226
rect 165554 472170 165622 472226
rect 165678 472170 165774 472226
rect 165154 472102 165774 472170
rect 165154 472046 165250 472102
rect 165306 472046 165374 472102
rect 165430 472046 165498 472102
rect 165554 472046 165622 472102
rect 165678 472046 165774 472102
rect 165154 471978 165774 472046
rect 165154 471922 165250 471978
rect 165306 471922 165374 471978
rect 165430 471922 165498 471978
rect 165554 471922 165622 471978
rect 165678 471922 165774 471978
rect 165154 458342 165774 471922
rect 168874 598172 169494 598268
rect 168874 598116 168970 598172
rect 169026 598116 169094 598172
rect 169150 598116 169218 598172
rect 169274 598116 169342 598172
rect 169398 598116 169494 598172
rect 168874 598048 169494 598116
rect 168874 597992 168970 598048
rect 169026 597992 169094 598048
rect 169150 597992 169218 598048
rect 169274 597992 169342 598048
rect 169398 597992 169494 598048
rect 168874 597924 169494 597992
rect 168874 597868 168970 597924
rect 169026 597868 169094 597924
rect 169150 597868 169218 597924
rect 169274 597868 169342 597924
rect 169398 597868 169494 597924
rect 168874 597800 169494 597868
rect 168874 597744 168970 597800
rect 169026 597744 169094 597800
rect 169150 597744 169218 597800
rect 169274 597744 169342 597800
rect 169398 597744 169494 597800
rect 168874 586350 169494 597744
rect 168874 586294 168970 586350
rect 169026 586294 169094 586350
rect 169150 586294 169218 586350
rect 169274 586294 169342 586350
rect 169398 586294 169494 586350
rect 168874 586226 169494 586294
rect 168874 586170 168970 586226
rect 169026 586170 169094 586226
rect 169150 586170 169218 586226
rect 169274 586170 169342 586226
rect 169398 586170 169494 586226
rect 168874 586102 169494 586170
rect 168874 586046 168970 586102
rect 169026 586046 169094 586102
rect 169150 586046 169218 586102
rect 169274 586046 169342 586102
rect 169398 586046 169494 586102
rect 168874 585978 169494 586046
rect 168874 585922 168970 585978
rect 169026 585922 169094 585978
rect 169150 585922 169218 585978
rect 169274 585922 169342 585978
rect 169398 585922 169494 585978
rect 168874 568350 169494 585922
rect 168874 568294 168970 568350
rect 169026 568294 169094 568350
rect 169150 568294 169218 568350
rect 169274 568294 169342 568350
rect 169398 568294 169494 568350
rect 168874 568226 169494 568294
rect 168874 568170 168970 568226
rect 169026 568170 169094 568226
rect 169150 568170 169218 568226
rect 169274 568170 169342 568226
rect 169398 568170 169494 568226
rect 168874 568102 169494 568170
rect 168874 568046 168970 568102
rect 169026 568046 169094 568102
rect 169150 568046 169218 568102
rect 169274 568046 169342 568102
rect 169398 568046 169494 568102
rect 168874 567978 169494 568046
rect 168874 567922 168970 567978
rect 169026 567922 169094 567978
rect 169150 567922 169218 567978
rect 169274 567922 169342 567978
rect 169398 567922 169494 567978
rect 168874 550350 169494 567922
rect 168874 550294 168970 550350
rect 169026 550294 169094 550350
rect 169150 550294 169218 550350
rect 169274 550294 169342 550350
rect 169398 550294 169494 550350
rect 168874 550226 169494 550294
rect 168874 550170 168970 550226
rect 169026 550170 169094 550226
rect 169150 550170 169218 550226
rect 169274 550170 169342 550226
rect 169398 550170 169494 550226
rect 168874 550102 169494 550170
rect 168874 550046 168970 550102
rect 169026 550046 169094 550102
rect 169150 550046 169218 550102
rect 169274 550046 169342 550102
rect 169398 550046 169494 550102
rect 168874 549978 169494 550046
rect 168874 549922 168970 549978
rect 169026 549922 169094 549978
rect 169150 549922 169218 549978
rect 169274 549922 169342 549978
rect 169398 549922 169494 549978
rect 168874 532350 169494 549922
rect 168874 532294 168970 532350
rect 169026 532294 169094 532350
rect 169150 532294 169218 532350
rect 169274 532294 169342 532350
rect 169398 532294 169494 532350
rect 168874 532226 169494 532294
rect 168874 532170 168970 532226
rect 169026 532170 169094 532226
rect 169150 532170 169218 532226
rect 169274 532170 169342 532226
rect 169398 532170 169494 532226
rect 168874 532102 169494 532170
rect 168874 532046 168970 532102
rect 169026 532046 169094 532102
rect 169150 532046 169218 532102
rect 169274 532046 169342 532102
rect 169398 532046 169494 532102
rect 168874 531978 169494 532046
rect 168874 531922 168970 531978
rect 169026 531922 169094 531978
rect 169150 531922 169218 531978
rect 169274 531922 169342 531978
rect 169398 531922 169494 531978
rect 168874 514350 169494 531922
rect 168874 514294 168970 514350
rect 169026 514294 169094 514350
rect 169150 514294 169218 514350
rect 169274 514294 169342 514350
rect 169398 514294 169494 514350
rect 168874 514226 169494 514294
rect 168874 514170 168970 514226
rect 169026 514170 169094 514226
rect 169150 514170 169218 514226
rect 169274 514170 169342 514226
rect 169398 514170 169494 514226
rect 168874 514102 169494 514170
rect 168874 514046 168970 514102
rect 169026 514046 169094 514102
rect 169150 514046 169218 514102
rect 169274 514046 169342 514102
rect 169398 514046 169494 514102
rect 168874 513978 169494 514046
rect 168874 513922 168970 513978
rect 169026 513922 169094 513978
rect 169150 513922 169218 513978
rect 169274 513922 169342 513978
rect 169398 513922 169494 513978
rect 168874 496350 169494 513922
rect 168874 496294 168970 496350
rect 169026 496294 169094 496350
rect 169150 496294 169218 496350
rect 169274 496294 169342 496350
rect 169398 496294 169494 496350
rect 168874 496226 169494 496294
rect 168874 496170 168970 496226
rect 169026 496170 169094 496226
rect 169150 496170 169218 496226
rect 169274 496170 169342 496226
rect 169398 496170 169494 496226
rect 168874 496102 169494 496170
rect 168874 496046 168970 496102
rect 169026 496046 169094 496102
rect 169150 496046 169218 496102
rect 169274 496046 169342 496102
rect 169398 496046 169494 496102
rect 168874 495978 169494 496046
rect 168874 495922 168970 495978
rect 169026 495922 169094 495978
rect 169150 495922 169218 495978
rect 169274 495922 169342 495978
rect 169398 495922 169494 495978
rect 168874 478350 169494 495922
rect 168874 478294 168970 478350
rect 169026 478294 169094 478350
rect 169150 478294 169218 478350
rect 169274 478294 169342 478350
rect 169398 478294 169494 478350
rect 168874 478226 169494 478294
rect 168874 478170 168970 478226
rect 169026 478170 169094 478226
rect 169150 478170 169218 478226
rect 169274 478170 169342 478226
rect 169398 478170 169494 478226
rect 168874 478102 169494 478170
rect 168874 478046 168970 478102
rect 169026 478046 169094 478102
rect 169150 478046 169218 478102
rect 169274 478046 169342 478102
rect 169398 478046 169494 478102
rect 168874 477978 169494 478046
rect 168874 477922 168970 477978
rect 169026 477922 169094 477978
rect 169150 477922 169218 477978
rect 169274 477922 169342 477978
rect 169398 477922 169494 477978
rect 168874 460350 169494 477922
rect 168874 460294 168970 460350
rect 169026 460294 169094 460350
rect 169150 460294 169218 460350
rect 169274 460294 169342 460350
rect 169398 460294 169494 460350
rect 168874 460226 169494 460294
rect 168874 460170 168970 460226
rect 169026 460170 169094 460226
rect 169150 460170 169218 460226
rect 169274 460170 169342 460226
rect 169398 460170 169494 460226
rect 168874 460102 169494 460170
rect 168874 460046 168970 460102
rect 169026 460046 169094 460102
rect 169150 460046 169218 460102
rect 169274 460046 169342 460102
rect 169398 460046 169494 460102
rect 168874 459978 169494 460046
rect 168874 459922 168970 459978
rect 169026 459922 169094 459978
rect 169150 459922 169218 459978
rect 169274 459922 169342 459978
rect 169398 459922 169494 459978
rect 168874 458342 169494 459922
rect 183154 597212 183774 598268
rect 183154 597156 183250 597212
rect 183306 597156 183374 597212
rect 183430 597156 183498 597212
rect 183554 597156 183622 597212
rect 183678 597156 183774 597212
rect 183154 597088 183774 597156
rect 183154 597032 183250 597088
rect 183306 597032 183374 597088
rect 183430 597032 183498 597088
rect 183554 597032 183622 597088
rect 183678 597032 183774 597088
rect 183154 596964 183774 597032
rect 183154 596908 183250 596964
rect 183306 596908 183374 596964
rect 183430 596908 183498 596964
rect 183554 596908 183622 596964
rect 183678 596908 183774 596964
rect 183154 596840 183774 596908
rect 183154 596784 183250 596840
rect 183306 596784 183374 596840
rect 183430 596784 183498 596840
rect 183554 596784 183622 596840
rect 183678 596784 183774 596840
rect 183154 580350 183774 596784
rect 183154 580294 183250 580350
rect 183306 580294 183374 580350
rect 183430 580294 183498 580350
rect 183554 580294 183622 580350
rect 183678 580294 183774 580350
rect 183154 580226 183774 580294
rect 183154 580170 183250 580226
rect 183306 580170 183374 580226
rect 183430 580170 183498 580226
rect 183554 580170 183622 580226
rect 183678 580170 183774 580226
rect 183154 580102 183774 580170
rect 183154 580046 183250 580102
rect 183306 580046 183374 580102
rect 183430 580046 183498 580102
rect 183554 580046 183622 580102
rect 183678 580046 183774 580102
rect 183154 579978 183774 580046
rect 183154 579922 183250 579978
rect 183306 579922 183374 579978
rect 183430 579922 183498 579978
rect 183554 579922 183622 579978
rect 183678 579922 183774 579978
rect 183154 562350 183774 579922
rect 183154 562294 183250 562350
rect 183306 562294 183374 562350
rect 183430 562294 183498 562350
rect 183554 562294 183622 562350
rect 183678 562294 183774 562350
rect 183154 562226 183774 562294
rect 183154 562170 183250 562226
rect 183306 562170 183374 562226
rect 183430 562170 183498 562226
rect 183554 562170 183622 562226
rect 183678 562170 183774 562226
rect 183154 562102 183774 562170
rect 183154 562046 183250 562102
rect 183306 562046 183374 562102
rect 183430 562046 183498 562102
rect 183554 562046 183622 562102
rect 183678 562046 183774 562102
rect 183154 561978 183774 562046
rect 183154 561922 183250 561978
rect 183306 561922 183374 561978
rect 183430 561922 183498 561978
rect 183554 561922 183622 561978
rect 183678 561922 183774 561978
rect 183154 544350 183774 561922
rect 183154 544294 183250 544350
rect 183306 544294 183374 544350
rect 183430 544294 183498 544350
rect 183554 544294 183622 544350
rect 183678 544294 183774 544350
rect 183154 544226 183774 544294
rect 183154 544170 183250 544226
rect 183306 544170 183374 544226
rect 183430 544170 183498 544226
rect 183554 544170 183622 544226
rect 183678 544170 183774 544226
rect 183154 544102 183774 544170
rect 183154 544046 183250 544102
rect 183306 544046 183374 544102
rect 183430 544046 183498 544102
rect 183554 544046 183622 544102
rect 183678 544046 183774 544102
rect 183154 543978 183774 544046
rect 183154 543922 183250 543978
rect 183306 543922 183374 543978
rect 183430 543922 183498 543978
rect 183554 543922 183622 543978
rect 183678 543922 183774 543978
rect 183154 526350 183774 543922
rect 183154 526294 183250 526350
rect 183306 526294 183374 526350
rect 183430 526294 183498 526350
rect 183554 526294 183622 526350
rect 183678 526294 183774 526350
rect 183154 526226 183774 526294
rect 183154 526170 183250 526226
rect 183306 526170 183374 526226
rect 183430 526170 183498 526226
rect 183554 526170 183622 526226
rect 183678 526170 183774 526226
rect 183154 526102 183774 526170
rect 183154 526046 183250 526102
rect 183306 526046 183374 526102
rect 183430 526046 183498 526102
rect 183554 526046 183622 526102
rect 183678 526046 183774 526102
rect 183154 525978 183774 526046
rect 183154 525922 183250 525978
rect 183306 525922 183374 525978
rect 183430 525922 183498 525978
rect 183554 525922 183622 525978
rect 183678 525922 183774 525978
rect 183154 508350 183774 525922
rect 183154 508294 183250 508350
rect 183306 508294 183374 508350
rect 183430 508294 183498 508350
rect 183554 508294 183622 508350
rect 183678 508294 183774 508350
rect 183154 508226 183774 508294
rect 183154 508170 183250 508226
rect 183306 508170 183374 508226
rect 183430 508170 183498 508226
rect 183554 508170 183622 508226
rect 183678 508170 183774 508226
rect 183154 508102 183774 508170
rect 183154 508046 183250 508102
rect 183306 508046 183374 508102
rect 183430 508046 183498 508102
rect 183554 508046 183622 508102
rect 183678 508046 183774 508102
rect 183154 507978 183774 508046
rect 183154 507922 183250 507978
rect 183306 507922 183374 507978
rect 183430 507922 183498 507978
rect 183554 507922 183622 507978
rect 183678 507922 183774 507978
rect 183154 490350 183774 507922
rect 183154 490294 183250 490350
rect 183306 490294 183374 490350
rect 183430 490294 183498 490350
rect 183554 490294 183622 490350
rect 183678 490294 183774 490350
rect 183154 490226 183774 490294
rect 183154 490170 183250 490226
rect 183306 490170 183374 490226
rect 183430 490170 183498 490226
rect 183554 490170 183622 490226
rect 183678 490170 183774 490226
rect 183154 490102 183774 490170
rect 183154 490046 183250 490102
rect 183306 490046 183374 490102
rect 183430 490046 183498 490102
rect 183554 490046 183622 490102
rect 183678 490046 183774 490102
rect 183154 489978 183774 490046
rect 183154 489922 183250 489978
rect 183306 489922 183374 489978
rect 183430 489922 183498 489978
rect 183554 489922 183622 489978
rect 183678 489922 183774 489978
rect 183154 472350 183774 489922
rect 183154 472294 183250 472350
rect 183306 472294 183374 472350
rect 183430 472294 183498 472350
rect 183554 472294 183622 472350
rect 183678 472294 183774 472350
rect 183154 472226 183774 472294
rect 183154 472170 183250 472226
rect 183306 472170 183374 472226
rect 183430 472170 183498 472226
rect 183554 472170 183622 472226
rect 183678 472170 183774 472226
rect 183154 472102 183774 472170
rect 183154 472046 183250 472102
rect 183306 472046 183374 472102
rect 183430 472046 183498 472102
rect 183554 472046 183622 472102
rect 183678 472046 183774 472102
rect 183154 471978 183774 472046
rect 183154 471922 183250 471978
rect 183306 471922 183374 471978
rect 183430 471922 183498 471978
rect 183554 471922 183622 471978
rect 183678 471922 183774 471978
rect 183154 458342 183774 471922
rect 186874 598172 187494 598268
rect 186874 598116 186970 598172
rect 187026 598116 187094 598172
rect 187150 598116 187218 598172
rect 187274 598116 187342 598172
rect 187398 598116 187494 598172
rect 186874 598048 187494 598116
rect 186874 597992 186970 598048
rect 187026 597992 187094 598048
rect 187150 597992 187218 598048
rect 187274 597992 187342 598048
rect 187398 597992 187494 598048
rect 186874 597924 187494 597992
rect 186874 597868 186970 597924
rect 187026 597868 187094 597924
rect 187150 597868 187218 597924
rect 187274 597868 187342 597924
rect 187398 597868 187494 597924
rect 186874 597800 187494 597868
rect 186874 597744 186970 597800
rect 187026 597744 187094 597800
rect 187150 597744 187218 597800
rect 187274 597744 187342 597800
rect 187398 597744 187494 597800
rect 186874 586350 187494 597744
rect 201154 597212 201774 598268
rect 201154 597156 201250 597212
rect 201306 597156 201374 597212
rect 201430 597156 201498 597212
rect 201554 597156 201622 597212
rect 201678 597156 201774 597212
rect 201154 597088 201774 597156
rect 201154 597032 201250 597088
rect 201306 597032 201374 597088
rect 201430 597032 201498 597088
rect 201554 597032 201622 597088
rect 201678 597032 201774 597088
rect 201154 596964 201774 597032
rect 201154 596908 201250 596964
rect 201306 596908 201374 596964
rect 201430 596908 201498 596964
rect 201554 596908 201622 596964
rect 201678 596908 201774 596964
rect 201154 596840 201774 596908
rect 201154 596784 201250 596840
rect 201306 596784 201374 596840
rect 201430 596784 201498 596840
rect 201554 596784 201622 596840
rect 201678 596784 201774 596840
rect 186874 586294 186970 586350
rect 187026 586294 187094 586350
rect 187150 586294 187218 586350
rect 187274 586294 187342 586350
rect 187398 586294 187494 586350
rect 186874 586226 187494 586294
rect 186874 586170 186970 586226
rect 187026 586170 187094 586226
rect 187150 586170 187218 586226
rect 187274 586170 187342 586226
rect 187398 586170 187494 586226
rect 186874 586102 187494 586170
rect 186874 586046 186970 586102
rect 187026 586046 187094 586102
rect 187150 586046 187218 586102
rect 187274 586046 187342 586102
rect 187398 586046 187494 586102
rect 186874 585978 187494 586046
rect 186874 585922 186970 585978
rect 187026 585922 187094 585978
rect 187150 585922 187218 585978
rect 187274 585922 187342 585978
rect 187398 585922 187494 585978
rect 186874 568350 187494 585922
rect 186874 568294 186970 568350
rect 187026 568294 187094 568350
rect 187150 568294 187218 568350
rect 187274 568294 187342 568350
rect 187398 568294 187494 568350
rect 186874 568226 187494 568294
rect 186874 568170 186970 568226
rect 187026 568170 187094 568226
rect 187150 568170 187218 568226
rect 187274 568170 187342 568226
rect 187398 568170 187494 568226
rect 186874 568102 187494 568170
rect 186874 568046 186970 568102
rect 187026 568046 187094 568102
rect 187150 568046 187218 568102
rect 187274 568046 187342 568102
rect 187398 568046 187494 568102
rect 186874 567978 187494 568046
rect 186874 567922 186970 567978
rect 187026 567922 187094 567978
rect 187150 567922 187218 567978
rect 187274 567922 187342 567978
rect 187398 567922 187494 567978
rect 186874 550350 187494 567922
rect 186874 550294 186970 550350
rect 187026 550294 187094 550350
rect 187150 550294 187218 550350
rect 187274 550294 187342 550350
rect 187398 550294 187494 550350
rect 186874 550226 187494 550294
rect 186874 550170 186970 550226
rect 187026 550170 187094 550226
rect 187150 550170 187218 550226
rect 187274 550170 187342 550226
rect 187398 550170 187494 550226
rect 186874 550102 187494 550170
rect 186874 550046 186970 550102
rect 187026 550046 187094 550102
rect 187150 550046 187218 550102
rect 187274 550046 187342 550102
rect 187398 550046 187494 550102
rect 186874 549978 187494 550046
rect 186874 549922 186970 549978
rect 187026 549922 187094 549978
rect 187150 549922 187218 549978
rect 187274 549922 187342 549978
rect 187398 549922 187494 549978
rect 186874 532350 187494 549922
rect 186874 532294 186970 532350
rect 187026 532294 187094 532350
rect 187150 532294 187218 532350
rect 187274 532294 187342 532350
rect 187398 532294 187494 532350
rect 186874 532226 187494 532294
rect 186874 532170 186970 532226
rect 187026 532170 187094 532226
rect 187150 532170 187218 532226
rect 187274 532170 187342 532226
rect 187398 532170 187494 532226
rect 186874 532102 187494 532170
rect 186874 532046 186970 532102
rect 187026 532046 187094 532102
rect 187150 532046 187218 532102
rect 187274 532046 187342 532102
rect 187398 532046 187494 532102
rect 186874 531978 187494 532046
rect 186874 531922 186970 531978
rect 187026 531922 187094 531978
rect 187150 531922 187218 531978
rect 187274 531922 187342 531978
rect 187398 531922 187494 531978
rect 186874 514350 187494 531922
rect 186874 514294 186970 514350
rect 187026 514294 187094 514350
rect 187150 514294 187218 514350
rect 187274 514294 187342 514350
rect 187398 514294 187494 514350
rect 186874 514226 187494 514294
rect 186874 514170 186970 514226
rect 187026 514170 187094 514226
rect 187150 514170 187218 514226
rect 187274 514170 187342 514226
rect 187398 514170 187494 514226
rect 186874 514102 187494 514170
rect 186874 514046 186970 514102
rect 187026 514046 187094 514102
rect 187150 514046 187218 514102
rect 187274 514046 187342 514102
rect 187398 514046 187494 514102
rect 186874 513978 187494 514046
rect 186874 513922 186970 513978
rect 187026 513922 187094 513978
rect 187150 513922 187218 513978
rect 187274 513922 187342 513978
rect 187398 513922 187494 513978
rect 186874 496350 187494 513922
rect 186874 496294 186970 496350
rect 187026 496294 187094 496350
rect 187150 496294 187218 496350
rect 187274 496294 187342 496350
rect 187398 496294 187494 496350
rect 186874 496226 187494 496294
rect 186874 496170 186970 496226
rect 187026 496170 187094 496226
rect 187150 496170 187218 496226
rect 187274 496170 187342 496226
rect 187398 496170 187494 496226
rect 186874 496102 187494 496170
rect 186874 496046 186970 496102
rect 187026 496046 187094 496102
rect 187150 496046 187218 496102
rect 187274 496046 187342 496102
rect 187398 496046 187494 496102
rect 186874 495978 187494 496046
rect 186874 495922 186970 495978
rect 187026 495922 187094 495978
rect 187150 495922 187218 495978
rect 187274 495922 187342 495978
rect 187398 495922 187494 495978
rect 186874 478350 187494 495922
rect 186874 478294 186970 478350
rect 187026 478294 187094 478350
rect 187150 478294 187218 478350
rect 187274 478294 187342 478350
rect 187398 478294 187494 478350
rect 186874 478226 187494 478294
rect 186874 478170 186970 478226
rect 187026 478170 187094 478226
rect 187150 478170 187218 478226
rect 187274 478170 187342 478226
rect 187398 478170 187494 478226
rect 186874 478102 187494 478170
rect 186874 478046 186970 478102
rect 187026 478046 187094 478102
rect 187150 478046 187218 478102
rect 187274 478046 187342 478102
rect 187398 478046 187494 478102
rect 186874 477978 187494 478046
rect 186874 477922 186970 477978
rect 187026 477922 187094 477978
rect 187150 477922 187218 477978
rect 187274 477922 187342 477978
rect 187398 477922 187494 477978
rect 186874 460350 187494 477922
rect 186874 460294 186970 460350
rect 187026 460294 187094 460350
rect 187150 460294 187218 460350
rect 187274 460294 187342 460350
rect 187398 460294 187494 460350
rect 186874 460226 187494 460294
rect 186874 460170 186970 460226
rect 187026 460170 187094 460226
rect 187150 460170 187218 460226
rect 187274 460170 187342 460226
rect 187398 460170 187494 460226
rect 186874 460102 187494 460170
rect 186874 460046 186970 460102
rect 187026 460046 187094 460102
rect 187150 460046 187218 460102
rect 187274 460046 187342 460102
rect 187398 460046 187494 460102
rect 186874 459978 187494 460046
rect 186874 459922 186970 459978
rect 187026 459922 187094 459978
rect 187150 459922 187218 459978
rect 187274 459922 187342 459978
rect 187398 459922 187494 459978
rect 186874 458342 187494 459922
rect 190652 587524 190708 587534
rect 24874 316350 25494 318858
rect 24874 316294 24970 316350
rect 25026 316294 25094 316350
rect 25150 316294 25218 316350
rect 25274 316294 25342 316350
rect 25398 316294 25494 316350
rect 24874 316226 25494 316294
rect 24874 316170 24970 316226
rect 25026 316170 25094 316226
rect 25150 316170 25218 316226
rect 25274 316170 25342 316226
rect 25398 316170 25494 316226
rect 24874 316102 25494 316170
rect 24874 316046 24970 316102
rect 25026 316046 25094 316102
rect 25150 316046 25218 316102
rect 25274 316046 25342 316102
rect 25398 316046 25494 316102
rect 24874 315978 25494 316046
rect 24874 315922 24970 315978
rect 25026 315922 25094 315978
rect 25150 315922 25218 315978
rect 25274 315922 25342 315978
rect 25398 315922 25494 315978
rect 24874 298422 25494 315922
rect 24874 298366 24970 298422
rect 25026 298366 25094 298422
rect 25150 298366 25218 298422
rect 25274 298366 25342 298422
rect 25398 298366 25494 298422
rect 24874 298342 25494 298366
rect 42874 316350 43494 318858
rect 42874 316294 42970 316350
rect 43026 316294 43094 316350
rect 43150 316294 43218 316350
rect 43274 316294 43342 316350
rect 43398 316294 43494 316350
rect 42874 316226 43494 316294
rect 42874 316170 42970 316226
rect 43026 316170 43094 316226
rect 43150 316170 43218 316226
rect 43274 316170 43342 316226
rect 43398 316170 43494 316226
rect 42874 316102 43494 316170
rect 42874 316046 42970 316102
rect 43026 316046 43094 316102
rect 43150 316046 43218 316102
rect 43274 316046 43342 316102
rect 43398 316046 43494 316102
rect 42874 315978 43494 316046
rect 42874 315922 42970 315978
rect 43026 315922 43094 315978
rect 43150 315922 43218 315978
rect 43274 315922 43342 315978
rect 43398 315922 43494 315978
rect 42874 298422 43494 315922
rect 42874 298366 42970 298422
rect 43026 298366 43094 298422
rect 43150 298366 43218 298422
rect 43274 298366 43342 298422
rect 43398 298366 43494 298422
rect 42874 298342 43494 298366
rect 60874 316350 61494 318858
rect 60874 316294 60970 316350
rect 61026 316294 61094 316350
rect 61150 316294 61218 316350
rect 61274 316294 61342 316350
rect 61398 316294 61494 316350
rect 60874 316226 61494 316294
rect 60874 316170 60970 316226
rect 61026 316170 61094 316226
rect 61150 316170 61218 316226
rect 61274 316170 61342 316226
rect 61398 316170 61494 316226
rect 60874 316102 61494 316170
rect 60874 316046 60970 316102
rect 61026 316046 61094 316102
rect 61150 316046 61218 316102
rect 61274 316046 61342 316102
rect 61398 316046 61494 316102
rect 60874 315978 61494 316046
rect 60874 315922 60970 315978
rect 61026 315922 61094 315978
rect 61150 315922 61218 315978
rect 61274 315922 61342 315978
rect 61398 315922 61494 315978
rect 60874 298422 61494 315922
rect 60874 298366 60970 298422
rect 61026 298366 61094 298422
rect 61150 298366 61218 298422
rect 61274 298366 61342 298422
rect 61398 298366 61494 298422
rect 60874 298342 61494 298366
rect 78874 316350 79494 318858
rect 78874 316294 78970 316350
rect 79026 316294 79094 316350
rect 79150 316294 79218 316350
rect 79274 316294 79342 316350
rect 79398 316294 79494 316350
rect 78874 316226 79494 316294
rect 78874 316170 78970 316226
rect 79026 316170 79094 316226
rect 79150 316170 79218 316226
rect 79274 316170 79342 316226
rect 79398 316170 79494 316226
rect 78874 316102 79494 316170
rect 78874 316046 78970 316102
rect 79026 316046 79094 316102
rect 79150 316046 79218 316102
rect 79274 316046 79342 316102
rect 79398 316046 79494 316102
rect 78874 315978 79494 316046
rect 78874 315922 78970 315978
rect 79026 315922 79094 315978
rect 79150 315922 79218 315978
rect 79274 315922 79342 315978
rect 79398 315922 79494 315978
rect 78874 298422 79494 315922
rect 78874 298366 78970 298422
rect 79026 298366 79094 298422
rect 79150 298366 79218 298422
rect 79274 298366 79342 298422
rect 79398 298366 79494 298422
rect 78874 298342 79494 298366
rect 96874 316350 97494 318858
rect 96874 316294 96970 316350
rect 97026 316294 97094 316350
rect 97150 316294 97218 316350
rect 97274 316294 97342 316350
rect 97398 316294 97494 316350
rect 96874 316226 97494 316294
rect 96874 316170 96970 316226
rect 97026 316170 97094 316226
rect 97150 316170 97218 316226
rect 97274 316170 97342 316226
rect 97398 316170 97494 316226
rect 96874 316102 97494 316170
rect 96874 316046 96970 316102
rect 97026 316046 97094 316102
rect 97150 316046 97218 316102
rect 97274 316046 97342 316102
rect 97398 316046 97494 316102
rect 96874 315978 97494 316046
rect 96874 315922 96970 315978
rect 97026 315922 97094 315978
rect 97150 315922 97218 315978
rect 97274 315922 97342 315978
rect 97398 315922 97494 315978
rect 96874 298422 97494 315922
rect 96874 298366 96970 298422
rect 97026 298366 97094 298422
rect 97150 298366 97218 298422
rect 97274 298366 97342 298422
rect 97398 298366 97494 298422
rect 96874 298342 97494 298366
rect 114874 316350 115494 318858
rect 114874 316294 114970 316350
rect 115026 316294 115094 316350
rect 115150 316294 115218 316350
rect 115274 316294 115342 316350
rect 115398 316294 115494 316350
rect 114874 316226 115494 316294
rect 114874 316170 114970 316226
rect 115026 316170 115094 316226
rect 115150 316170 115218 316226
rect 115274 316170 115342 316226
rect 115398 316170 115494 316226
rect 114874 316102 115494 316170
rect 114874 316046 114970 316102
rect 115026 316046 115094 316102
rect 115150 316046 115218 316102
rect 115274 316046 115342 316102
rect 115398 316046 115494 316102
rect 114874 315978 115494 316046
rect 114874 315922 114970 315978
rect 115026 315922 115094 315978
rect 115150 315922 115218 315978
rect 115274 315922 115342 315978
rect 115398 315922 115494 315978
rect 114874 298422 115494 315922
rect 114874 298366 114970 298422
rect 115026 298366 115094 298422
rect 115150 298366 115218 298422
rect 115274 298366 115342 298422
rect 115398 298366 115494 298422
rect 114874 298342 115494 298366
rect 132874 316350 133494 318858
rect 132874 316294 132970 316350
rect 133026 316294 133094 316350
rect 133150 316294 133218 316350
rect 133274 316294 133342 316350
rect 133398 316294 133494 316350
rect 132874 316226 133494 316294
rect 132874 316170 132970 316226
rect 133026 316170 133094 316226
rect 133150 316170 133218 316226
rect 133274 316170 133342 316226
rect 133398 316170 133494 316226
rect 132874 316102 133494 316170
rect 132874 316046 132970 316102
rect 133026 316046 133094 316102
rect 133150 316046 133218 316102
rect 133274 316046 133342 316102
rect 133398 316046 133494 316102
rect 132874 315978 133494 316046
rect 132874 315922 132970 315978
rect 133026 315922 133094 315978
rect 133150 315922 133218 315978
rect 133274 315922 133342 315978
rect 133398 315922 133494 315978
rect 132874 298422 133494 315922
rect 132874 298366 132970 298422
rect 133026 298366 133094 298422
rect 133150 298366 133218 298422
rect 133274 298366 133342 298422
rect 133398 298366 133494 298422
rect 132874 298342 133494 298366
rect 150874 316350 151494 318858
rect 150874 316294 150970 316350
rect 151026 316294 151094 316350
rect 151150 316294 151218 316350
rect 151274 316294 151342 316350
rect 151398 316294 151494 316350
rect 150874 316226 151494 316294
rect 150874 316170 150970 316226
rect 151026 316170 151094 316226
rect 151150 316170 151218 316226
rect 151274 316170 151342 316226
rect 151398 316170 151494 316226
rect 150874 316102 151494 316170
rect 150874 316046 150970 316102
rect 151026 316046 151094 316102
rect 151150 316046 151218 316102
rect 151274 316046 151342 316102
rect 151398 316046 151494 316102
rect 150874 315978 151494 316046
rect 150874 315922 150970 315978
rect 151026 315922 151094 315978
rect 151150 315922 151218 315978
rect 151274 315922 151342 315978
rect 151398 315922 151494 315978
rect 150874 298422 151494 315922
rect 150874 298366 150970 298422
rect 151026 298366 151094 298422
rect 151150 298366 151218 298422
rect 151274 298366 151342 298422
rect 151398 298366 151494 298422
rect 150874 298342 151494 298366
rect 168874 316350 169494 318858
rect 168874 316294 168970 316350
rect 169026 316294 169094 316350
rect 169150 316294 169218 316350
rect 169274 316294 169342 316350
rect 169398 316294 169494 316350
rect 168874 316226 169494 316294
rect 168874 316170 168970 316226
rect 169026 316170 169094 316226
rect 169150 316170 169218 316226
rect 169274 316170 169342 316226
rect 169398 316170 169494 316226
rect 168874 316102 169494 316170
rect 168874 316046 168970 316102
rect 169026 316046 169094 316102
rect 169150 316046 169218 316102
rect 169274 316046 169342 316102
rect 169398 316046 169494 316102
rect 168874 315978 169494 316046
rect 168874 315922 168970 315978
rect 169026 315922 169094 315978
rect 169150 315922 169218 315978
rect 169274 315922 169342 315978
rect 169398 315922 169494 315978
rect 168874 298422 169494 315922
rect 168874 298366 168970 298422
rect 169026 298366 169094 298422
rect 169150 298366 169218 298422
rect 169274 298366 169342 298422
rect 169398 298366 169494 298422
rect 168874 298342 169494 298366
rect 186874 316350 187494 318858
rect 186874 316294 186970 316350
rect 187026 316294 187094 316350
rect 187150 316294 187218 316350
rect 187274 316294 187342 316350
rect 187398 316294 187494 316350
rect 186874 316226 187494 316294
rect 186874 316170 186970 316226
rect 187026 316170 187094 316226
rect 187150 316170 187218 316226
rect 187274 316170 187342 316226
rect 187398 316170 187494 316226
rect 186874 316102 187494 316170
rect 186874 316046 186970 316102
rect 187026 316046 187094 316102
rect 187150 316046 187218 316102
rect 187274 316046 187342 316102
rect 187398 316046 187494 316102
rect 186874 315978 187494 316046
rect 186874 315922 186970 315978
rect 187026 315922 187094 315978
rect 187150 315922 187218 315978
rect 187274 315922 187342 315978
rect 187398 315922 187494 315978
rect 186874 298422 187494 315922
rect 189196 316820 189252 316830
rect 189084 308308 189140 308318
rect 186874 298366 186970 298422
rect 187026 298366 187094 298422
rect 187150 298366 187218 298422
rect 187274 298366 187342 298422
rect 187398 298366 187494 298422
rect 186874 298342 187494 298366
rect 188972 306628 189028 306638
rect 21154 148350 21774 158858
rect 21154 148294 21250 148350
rect 21306 148294 21374 148350
rect 21430 148294 21498 148350
rect 21554 148294 21622 148350
rect 21678 148294 21774 148350
rect 21154 148226 21774 148294
rect 21154 148170 21250 148226
rect 21306 148170 21374 148226
rect 21430 148170 21498 148226
rect 21554 148170 21622 148226
rect 21678 148170 21774 148226
rect 21154 148102 21774 148170
rect 21154 148046 21250 148102
rect 21306 148046 21374 148102
rect 21430 148046 21498 148102
rect 21554 148046 21622 148102
rect 21678 148046 21774 148102
rect 21154 147978 21774 148046
rect 21154 147922 21250 147978
rect 21306 147922 21374 147978
rect 21430 147922 21498 147978
rect 21554 147922 21622 147978
rect 21678 147922 21774 147978
rect 21154 130350 21774 147922
rect 21154 130294 21250 130350
rect 21306 130294 21374 130350
rect 21430 130294 21498 130350
rect 21554 130294 21622 130350
rect 21678 130294 21774 130350
rect 21154 130226 21774 130294
rect 21154 130170 21250 130226
rect 21306 130170 21374 130226
rect 21430 130170 21498 130226
rect 21554 130170 21622 130226
rect 21678 130170 21774 130226
rect 21154 130102 21774 130170
rect 21154 130046 21250 130102
rect 21306 130046 21374 130102
rect 21430 130046 21498 130102
rect 21554 130046 21622 130102
rect 21678 130046 21774 130102
rect 21154 129978 21774 130046
rect 21154 129922 21250 129978
rect 21306 129922 21374 129978
rect 21430 129922 21498 129978
rect 21554 129922 21622 129978
rect 21678 129922 21774 129978
rect 19516 114436 19572 114446
rect 19404 107716 19460 107726
rect 16268 102340 16324 102350
rect 16156 92932 16212 92942
rect 9996 18386 10052 18396
rect 16044 87556 16100 87566
rect 7644 16706 7700 16716
rect 6874 10294 6970 10350
rect 7026 10294 7094 10350
rect 7150 10294 7218 10350
rect 7274 10294 7342 10350
rect 7398 10294 7494 10350
rect 6874 10226 7494 10294
rect 6874 10170 6970 10226
rect 7026 10170 7094 10226
rect 7150 10170 7218 10226
rect 7274 10170 7342 10226
rect 7398 10170 7494 10226
rect 6874 10102 7494 10170
rect 6874 10046 6970 10102
rect 7026 10046 7094 10102
rect 7150 10046 7218 10102
rect 7274 10046 7342 10102
rect 7398 10046 7494 10102
rect 6874 9978 7494 10046
rect 16044 10052 16100 87500
rect 16156 14868 16212 92876
rect 16268 14980 16324 102284
rect 19180 95620 19236 95630
rect 18396 84868 18452 84878
rect 18284 70980 18340 70990
rect 16268 14914 16324 14924
rect 18172 70756 18228 70766
rect 16156 14802 16212 14812
rect 18172 12964 18228 70700
rect 18284 13300 18340 70924
rect 18396 14644 18452 84812
rect 19180 16660 19236 95564
rect 19180 16594 19236 16604
rect 18396 14578 18452 14588
rect 18284 13234 18340 13244
rect 19404 13188 19460 107660
rect 19516 68516 19572 114380
rect 21154 112350 21774 129922
rect 21154 112294 21250 112350
rect 21306 112294 21374 112350
rect 21430 112294 21498 112350
rect 21554 112294 21622 112350
rect 21678 112294 21774 112350
rect 21154 112226 21774 112294
rect 21154 112170 21250 112226
rect 21306 112170 21374 112226
rect 21430 112170 21498 112226
rect 21554 112170 21622 112226
rect 21678 112170 21774 112226
rect 21154 112102 21774 112170
rect 21154 112046 21250 112102
rect 21306 112046 21374 112102
rect 21430 112046 21498 112102
rect 21554 112046 21622 112102
rect 21678 112046 21774 112102
rect 21154 111978 21774 112046
rect 21154 111922 21250 111978
rect 21306 111922 21374 111978
rect 21430 111922 21498 111978
rect 21554 111922 21622 111978
rect 21678 111922 21774 111978
rect 19964 100996 20020 101006
rect 19740 94276 19796 94286
rect 19516 68450 19572 68460
rect 19628 90244 19684 90254
rect 19628 16436 19684 90188
rect 19740 18340 19796 94220
rect 19740 18274 19796 18284
rect 19628 16370 19684 16380
rect 19964 14756 20020 100940
rect 21154 94350 21774 111922
rect 21154 94294 21250 94350
rect 21306 94294 21374 94350
rect 21430 94294 21498 94350
rect 21554 94294 21622 94350
rect 21678 94294 21774 94350
rect 21154 94226 21774 94294
rect 21154 94170 21250 94226
rect 21306 94170 21374 94226
rect 21430 94170 21498 94226
rect 21554 94170 21622 94226
rect 21678 94170 21774 94226
rect 21154 94102 21774 94170
rect 21154 94046 21250 94102
rect 21306 94046 21374 94102
rect 21430 94046 21498 94102
rect 21554 94046 21622 94102
rect 21678 94046 21774 94102
rect 21154 93978 21774 94046
rect 21154 93922 21250 93978
rect 21306 93922 21374 93978
rect 21430 93922 21498 93978
rect 21554 93922 21622 93978
rect 21678 93922 21774 93978
rect 20076 91588 20132 91598
rect 20076 69860 20132 91532
rect 20300 83524 20356 83534
rect 20076 69794 20132 69804
rect 20188 80836 20244 80846
rect 20188 16324 20244 80780
rect 20300 19684 20356 83468
rect 21154 76350 21774 93922
rect 24874 154350 25494 158858
rect 24874 154294 24970 154350
rect 25026 154294 25094 154350
rect 25150 154294 25218 154350
rect 25274 154294 25342 154350
rect 25398 154294 25494 154350
rect 24874 154226 25494 154294
rect 24874 154170 24970 154226
rect 25026 154170 25094 154226
rect 25150 154170 25218 154226
rect 25274 154170 25342 154226
rect 25398 154170 25494 154226
rect 24874 154102 25494 154170
rect 24874 154046 24970 154102
rect 25026 154046 25094 154102
rect 25150 154046 25218 154102
rect 25274 154046 25342 154102
rect 25398 154046 25494 154102
rect 24874 153978 25494 154046
rect 24874 153922 24970 153978
rect 25026 153922 25094 153978
rect 25150 153922 25218 153978
rect 25274 153922 25342 153978
rect 25398 153922 25494 153978
rect 24874 136350 25494 153922
rect 24874 136294 24970 136350
rect 25026 136294 25094 136350
rect 25150 136294 25218 136350
rect 25274 136294 25342 136350
rect 25398 136294 25494 136350
rect 24874 136226 25494 136294
rect 24874 136170 24970 136226
rect 25026 136170 25094 136226
rect 25150 136170 25218 136226
rect 25274 136170 25342 136226
rect 25398 136170 25494 136226
rect 24874 136102 25494 136170
rect 24874 136046 24970 136102
rect 25026 136046 25094 136102
rect 25150 136046 25218 136102
rect 25274 136046 25342 136102
rect 25398 136046 25494 136102
rect 24874 135978 25494 136046
rect 24874 135922 24970 135978
rect 25026 135922 25094 135978
rect 25150 135922 25218 135978
rect 25274 135922 25342 135978
rect 25398 135922 25494 135978
rect 24874 118350 25494 135922
rect 24874 118294 24970 118350
rect 25026 118294 25094 118350
rect 25150 118294 25218 118350
rect 25274 118294 25342 118350
rect 25398 118294 25494 118350
rect 24874 118226 25494 118294
rect 24874 118170 24970 118226
rect 25026 118170 25094 118226
rect 25150 118170 25218 118226
rect 25274 118170 25342 118226
rect 25398 118170 25494 118226
rect 24874 118102 25494 118170
rect 24874 118046 24970 118102
rect 25026 118046 25094 118102
rect 25150 118046 25218 118102
rect 25274 118046 25342 118102
rect 25398 118046 25494 118102
rect 24874 117978 25494 118046
rect 24874 117922 24970 117978
rect 25026 117922 25094 117978
rect 25150 117922 25218 117978
rect 25274 117922 25342 117978
rect 25398 117922 25494 117978
rect 24874 100350 25494 117922
rect 24874 100294 24970 100350
rect 25026 100294 25094 100350
rect 25150 100294 25218 100350
rect 25274 100294 25342 100350
rect 25398 100294 25494 100350
rect 24874 100226 25494 100294
rect 24874 100170 24970 100226
rect 25026 100170 25094 100226
rect 25150 100170 25218 100226
rect 25274 100170 25342 100226
rect 25398 100170 25494 100226
rect 24874 100102 25494 100170
rect 24874 100046 24970 100102
rect 25026 100046 25094 100102
rect 25150 100046 25218 100102
rect 25274 100046 25342 100102
rect 25398 100046 25494 100102
rect 24874 99978 25494 100046
rect 24874 99922 24970 99978
rect 25026 99922 25094 99978
rect 25150 99922 25218 99978
rect 25274 99922 25342 99978
rect 25398 99922 25494 99978
rect 22204 86212 22260 86222
rect 22204 78988 22260 86156
rect 24874 82350 25494 99922
rect 24874 82294 24970 82350
rect 25026 82294 25094 82350
rect 25150 82294 25218 82350
rect 25274 82294 25342 82350
rect 25398 82294 25494 82350
rect 24874 82226 25494 82294
rect 22316 82180 22372 82190
rect 22372 82124 22820 82180
rect 22316 82114 22372 82124
rect 22204 78932 22708 78988
rect 21154 76294 21250 76350
rect 21306 76294 21374 76350
rect 21430 76294 21498 76350
rect 21554 76294 21622 76350
rect 21678 76294 21774 76350
rect 21154 76226 21774 76294
rect 21154 76170 21250 76226
rect 21306 76170 21374 76226
rect 21430 76170 21498 76226
rect 21554 76170 21622 76226
rect 21678 76170 21774 76226
rect 21154 76102 21774 76170
rect 21154 76046 21250 76102
rect 21306 76046 21374 76102
rect 21430 76046 21498 76102
rect 21554 76046 21622 76102
rect 21678 76046 21774 76102
rect 21154 75978 21774 76046
rect 21154 75922 21250 75978
rect 21306 75922 21374 75978
rect 21430 75922 21498 75978
rect 21554 75922 21622 75978
rect 21678 75922 21774 75978
rect 20300 19618 20356 19628
rect 20972 72548 21028 72558
rect 20188 16258 20244 16268
rect 19964 14690 20020 14700
rect 19404 13122 19460 13132
rect 20972 13076 21028 72492
rect 20972 13010 21028 13020
rect 21154 58350 21774 75922
rect 22092 73668 22148 73678
rect 22148 73612 22260 73668
rect 22092 73602 22148 73612
rect 21980 73556 22036 73566
rect 21980 70644 22036 73500
rect 22092 73444 22148 73454
rect 22092 70756 22148 73388
rect 22092 70690 22148 70700
rect 21980 70578 22036 70588
rect 22204 70532 22260 73612
rect 22204 70466 22260 70476
rect 21154 58294 21250 58350
rect 21306 58294 21374 58350
rect 21430 58294 21498 58350
rect 21554 58294 21622 58350
rect 21678 58294 21774 58350
rect 21154 58226 21774 58294
rect 21154 58170 21250 58226
rect 21306 58170 21374 58226
rect 21430 58170 21498 58226
rect 21554 58170 21622 58226
rect 21678 58170 21774 58226
rect 21154 58102 21774 58170
rect 21154 58046 21250 58102
rect 21306 58046 21374 58102
rect 21430 58046 21498 58102
rect 21554 58046 21622 58102
rect 21678 58046 21774 58102
rect 21154 57978 21774 58046
rect 21154 57922 21250 57978
rect 21306 57922 21374 57978
rect 21430 57922 21498 57978
rect 21554 57922 21622 57978
rect 21678 57922 21774 57978
rect 21154 40350 21774 57922
rect 21154 40294 21250 40350
rect 21306 40294 21374 40350
rect 21430 40294 21498 40350
rect 21554 40294 21622 40350
rect 21678 40294 21774 40350
rect 21154 40226 21774 40294
rect 21154 40170 21250 40226
rect 21306 40170 21374 40226
rect 21430 40170 21498 40226
rect 21554 40170 21622 40226
rect 21678 40170 21774 40226
rect 21154 40102 21774 40170
rect 21154 40046 21250 40102
rect 21306 40046 21374 40102
rect 21430 40046 21498 40102
rect 21554 40046 21622 40102
rect 21678 40046 21774 40102
rect 21154 39978 21774 40046
rect 21154 39922 21250 39978
rect 21306 39922 21374 39978
rect 21430 39922 21498 39978
rect 21554 39922 21622 39978
rect 21678 39922 21774 39978
rect 21154 22350 21774 39922
rect 21154 22294 21250 22350
rect 21306 22294 21374 22350
rect 21430 22294 21498 22350
rect 21554 22294 21622 22350
rect 21678 22294 21774 22350
rect 21154 22226 21774 22294
rect 21154 22170 21250 22226
rect 21306 22170 21374 22226
rect 21430 22170 21498 22226
rect 21554 22170 21622 22226
rect 21678 22170 21774 22226
rect 21154 22102 21774 22170
rect 21154 22046 21250 22102
rect 21306 22046 21374 22102
rect 21430 22046 21498 22102
rect 21554 22046 21622 22102
rect 21678 22046 21774 22102
rect 21154 21978 21774 22046
rect 21154 21922 21250 21978
rect 21306 21922 21374 21978
rect 21430 21922 21498 21978
rect 21554 21922 21622 21978
rect 21678 21922 21774 21978
rect 18172 12898 18228 12908
rect 16044 9986 16100 9996
rect 6874 9922 6970 9978
rect 7026 9922 7094 9978
rect 7150 9922 7218 9978
rect 7274 9922 7342 9978
rect 7398 9922 7494 9978
rect 6874 -1120 7494 9922
rect 6874 -1176 6970 -1120
rect 7026 -1176 7094 -1120
rect 7150 -1176 7218 -1120
rect 7274 -1176 7342 -1120
rect 7398 -1176 7494 -1120
rect 6874 -1244 7494 -1176
rect 6874 -1300 6970 -1244
rect 7026 -1300 7094 -1244
rect 7150 -1300 7218 -1244
rect 7274 -1300 7342 -1244
rect 7398 -1300 7494 -1244
rect 6874 -1368 7494 -1300
rect 6874 -1424 6970 -1368
rect 7026 -1424 7094 -1368
rect 7150 -1424 7218 -1368
rect 7274 -1424 7342 -1368
rect 7398 -1424 7494 -1368
rect 6874 -1492 7494 -1424
rect 6874 -1548 6970 -1492
rect 7026 -1548 7094 -1492
rect 7150 -1548 7218 -1492
rect 7274 -1548 7342 -1492
rect 7398 -1548 7494 -1492
rect 6874 -1644 7494 -1548
rect 21154 4350 21774 21922
rect 22652 21028 22708 78932
rect 22652 20962 22708 20972
rect 22764 18116 22820 82124
rect 24874 82170 24970 82226
rect 25026 82170 25094 82226
rect 25150 82170 25218 82226
rect 25274 82170 25342 82226
rect 25398 82170 25494 82226
rect 24874 82102 25494 82170
rect 24874 82046 24970 82102
rect 25026 82046 25094 82102
rect 25150 82046 25218 82102
rect 25274 82046 25342 82102
rect 25398 82046 25494 82102
rect 24874 81978 25494 82046
rect 24874 81922 24970 81978
rect 25026 81922 25094 81978
rect 25150 81922 25218 81978
rect 25274 81922 25342 81978
rect 25398 81922 25494 81978
rect 23324 70756 23380 70766
rect 22764 18050 22820 18060
rect 22876 70644 22932 70654
rect 22876 14532 22932 70588
rect 23100 70532 23156 70542
rect 23100 18228 23156 70476
rect 23324 19572 23380 70700
rect 23324 19506 23380 19516
rect 24874 64350 25494 81922
rect 39154 148350 39774 158858
rect 39154 148294 39250 148350
rect 39306 148294 39374 148350
rect 39430 148294 39498 148350
rect 39554 148294 39622 148350
rect 39678 148294 39774 148350
rect 39154 148226 39774 148294
rect 39154 148170 39250 148226
rect 39306 148170 39374 148226
rect 39430 148170 39498 148226
rect 39554 148170 39622 148226
rect 39678 148170 39774 148226
rect 39154 148102 39774 148170
rect 39154 148046 39250 148102
rect 39306 148046 39374 148102
rect 39430 148046 39498 148102
rect 39554 148046 39622 148102
rect 39678 148046 39774 148102
rect 39154 147978 39774 148046
rect 39154 147922 39250 147978
rect 39306 147922 39374 147978
rect 39430 147922 39498 147978
rect 39554 147922 39622 147978
rect 39678 147922 39774 147978
rect 39154 130350 39774 147922
rect 39154 130294 39250 130350
rect 39306 130294 39374 130350
rect 39430 130294 39498 130350
rect 39554 130294 39622 130350
rect 39678 130294 39774 130350
rect 39154 130226 39774 130294
rect 39154 130170 39250 130226
rect 39306 130170 39374 130226
rect 39430 130170 39498 130226
rect 39554 130170 39622 130226
rect 39678 130170 39774 130226
rect 39154 130102 39774 130170
rect 39154 130046 39250 130102
rect 39306 130046 39374 130102
rect 39430 130046 39498 130102
rect 39554 130046 39622 130102
rect 39678 130046 39774 130102
rect 39154 129978 39774 130046
rect 39154 129922 39250 129978
rect 39306 129922 39374 129978
rect 39430 129922 39498 129978
rect 39554 129922 39622 129978
rect 39678 129922 39774 129978
rect 39154 112350 39774 129922
rect 39154 112294 39250 112350
rect 39306 112294 39374 112350
rect 39430 112294 39498 112350
rect 39554 112294 39622 112350
rect 39678 112294 39774 112350
rect 39154 112226 39774 112294
rect 39154 112170 39250 112226
rect 39306 112170 39374 112226
rect 39430 112170 39498 112226
rect 39554 112170 39622 112226
rect 39678 112170 39774 112226
rect 39154 112102 39774 112170
rect 39154 112046 39250 112102
rect 39306 112046 39374 112102
rect 39430 112046 39498 112102
rect 39554 112046 39622 112102
rect 39678 112046 39774 112102
rect 39154 111978 39774 112046
rect 39154 111922 39250 111978
rect 39306 111922 39374 111978
rect 39430 111922 39498 111978
rect 39554 111922 39622 111978
rect 39678 111922 39774 111978
rect 39154 94350 39774 111922
rect 39154 94294 39250 94350
rect 39306 94294 39374 94350
rect 39430 94294 39498 94350
rect 39554 94294 39622 94350
rect 39678 94294 39774 94350
rect 39154 94226 39774 94294
rect 39154 94170 39250 94226
rect 39306 94170 39374 94226
rect 39430 94170 39498 94226
rect 39554 94170 39622 94226
rect 39678 94170 39774 94226
rect 39154 94102 39774 94170
rect 39154 94046 39250 94102
rect 39306 94046 39374 94102
rect 39430 94046 39498 94102
rect 39554 94046 39622 94102
rect 39678 94046 39774 94102
rect 39154 93978 39774 94046
rect 39154 93922 39250 93978
rect 39306 93922 39374 93978
rect 39430 93922 39498 93978
rect 39554 93922 39622 93978
rect 39678 93922 39774 93978
rect 39154 76350 39774 93922
rect 39154 76294 39250 76350
rect 39306 76294 39374 76350
rect 39430 76294 39498 76350
rect 39554 76294 39622 76350
rect 39678 76294 39774 76350
rect 39154 76226 39774 76294
rect 39154 76170 39250 76226
rect 39306 76170 39374 76226
rect 39430 76170 39498 76226
rect 39554 76170 39622 76226
rect 39678 76170 39774 76226
rect 39154 76102 39774 76170
rect 39154 76046 39250 76102
rect 39306 76046 39374 76102
rect 39430 76046 39498 76102
rect 39554 76046 39622 76102
rect 39678 76046 39774 76102
rect 39154 75978 39774 76046
rect 39154 75922 39250 75978
rect 39306 75922 39374 75978
rect 39430 75922 39498 75978
rect 39554 75922 39622 75978
rect 39678 75922 39774 75978
rect 36988 68628 37044 68638
rect 24874 64294 24970 64350
rect 25026 64294 25094 64350
rect 25150 64294 25218 64350
rect 25274 64294 25342 64350
rect 25398 64294 25494 64350
rect 24874 64226 25494 64294
rect 24874 64170 24970 64226
rect 25026 64170 25094 64226
rect 25150 64170 25218 64226
rect 25274 64170 25342 64226
rect 25398 64170 25494 64226
rect 24874 64102 25494 64170
rect 24874 64046 24970 64102
rect 25026 64046 25094 64102
rect 25150 64046 25218 64102
rect 25274 64046 25342 64102
rect 25398 64046 25494 64102
rect 24874 63978 25494 64046
rect 24874 63922 24970 63978
rect 25026 63922 25094 63978
rect 25150 63922 25218 63978
rect 25274 63922 25342 63978
rect 25398 63922 25494 63978
rect 24874 46350 25494 63922
rect 24874 46294 24970 46350
rect 25026 46294 25094 46350
rect 25150 46294 25218 46350
rect 25274 46294 25342 46350
rect 25398 46294 25494 46350
rect 24874 46226 25494 46294
rect 24874 46170 24970 46226
rect 25026 46170 25094 46226
rect 25150 46170 25218 46226
rect 25274 46170 25342 46226
rect 25398 46170 25494 46226
rect 24874 46102 25494 46170
rect 24874 46046 24970 46102
rect 25026 46046 25094 46102
rect 25150 46046 25218 46102
rect 25274 46046 25342 46102
rect 25398 46046 25494 46102
rect 24874 45978 25494 46046
rect 24874 45922 24970 45978
rect 25026 45922 25094 45978
rect 25150 45922 25218 45978
rect 25274 45922 25342 45978
rect 25398 45922 25494 45978
rect 24874 28350 25494 45922
rect 24874 28294 24970 28350
rect 25026 28294 25094 28350
rect 25150 28294 25218 28350
rect 25274 28294 25342 28350
rect 25398 28294 25494 28350
rect 24874 28226 25494 28294
rect 24874 28170 24970 28226
rect 25026 28170 25094 28226
rect 25150 28170 25218 28226
rect 25274 28170 25342 28226
rect 25398 28170 25494 28226
rect 24874 28102 25494 28170
rect 24874 28046 24970 28102
rect 25026 28046 25094 28102
rect 25150 28046 25218 28102
rect 25274 28046 25342 28102
rect 25398 28046 25494 28102
rect 24874 27978 25494 28046
rect 24874 27922 24970 27978
rect 25026 27922 25094 27978
rect 25150 27922 25218 27978
rect 25274 27922 25342 27978
rect 25398 27922 25494 27978
rect 23100 18162 23156 18172
rect 22876 14466 22932 14476
rect 21154 4294 21250 4350
rect 21306 4294 21374 4350
rect 21430 4294 21498 4350
rect 21554 4294 21622 4350
rect 21678 4294 21774 4350
rect 21154 4226 21774 4294
rect 21154 4170 21250 4226
rect 21306 4170 21374 4226
rect 21430 4170 21498 4226
rect 21554 4170 21622 4226
rect 21678 4170 21774 4226
rect 21154 4102 21774 4170
rect 21154 4046 21250 4102
rect 21306 4046 21374 4102
rect 21430 4046 21498 4102
rect 21554 4046 21622 4102
rect 21678 4046 21774 4102
rect 21154 3978 21774 4046
rect 21154 3922 21250 3978
rect 21306 3922 21374 3978
rect 21430 3922 21498 3978
rect 21554 3922 21622 3978
rect 21678 3922 21774 3978
rect 21154 -160 21774 3922
rect 21154 -216 21250 -160
rect 21306 -216 21374 -160
rect 21430 -216 21498 -160
rect 21554 -216 21622 -160
rect 21678 -216 21774 -160
rect 21154 -284 21774 -216
rect 21154 -340 21250 -284
rect 21306 -340 21374 -284
rect 21430 -340 21498 -284
rect 21554 -340 21622 -284
rect 21678 -340 21774 -284
rect 21154 -408 21774 -340
rect 21154 -464 21250 -408
rect 21306 -464 21374 -408
rect 21430 -464 21498 -408
rect 21554 -464 21622 -408
rect 21678 -464 21774 -408
rect 21154 -532 21774 -464
rect 21154 -588 21250 -532
rect 21306 -588 21374 -532
rect 21430 -588 21498 -532
rect 21554 -588 21622 -532
rect 21678 -588 21774 -532
rect 21154 -1644 21774 -588
rect 24874 10350 25494 27922
rect 25564 68404 25620 68414
rect 25564 20132 25620 68348
rect 25564 20066 25620 20076
rect 28588 68404 28644 68414
rect 24874 10294 24970 10350
rect 25026 10294 25094 10350
rect 25150 10294 25218 10350
rect 25274 10294 25342 10350
rect 25398 10294 25494 10350
rect 24874 10226 25494 10294
rect 24874 10170 24970 10226
rect 25026 10170 25094 10226
rect 25150 10170 25218 10226
rect 25274 10170 25342 10226
rect 25398 10170 25494 10226
rect 24874 10102 25494 10170
rect 24874 10046 24970 10102
rect 25026 10046 25094 10102
rect 25150 10046 25218 10102
rect 25274 10046 25342 10102
rect 25398 10046 25494 10102
rect 24874 9978 25494 10046
rect 24874 9922 24970 9978
rect 25026 9922 25094 9978
rect 25150 9922 25218 9978
rect 25274 9922 25342 9978
rect 25398 9922 25494 9978
rect 24874 -1120 25494 9922
rect 28588 6804 28644 68348
rect 36988 16212 37044 68572
rect 36988 16146 37044 16156
rect 39154 58350 39774 75922
rect 42874 154350 43494 158858
rect 42874 154294 42970 154350
rect 43026 154294 43094 154350
rect 43150 154294 43218 154350
rect 43274 154294 43342 154350
rect 43398 154294 43494 154350
rect 42874 154226 43494 154294
rect 42874 154170 42970 154226
rect 43026 154170 43094 154226
rect 43150 154170 43218 154226
rect 43274 154170 43342 154226
rect 43398 154170 43494 154226
rect 42874 154102 43494 154170
rect 42874 154046 42970 154102
rect 43026 154046 43094 154102
rect 43150 154046 43218 154102
rect 43274 154046 43342 154102
rect 43398 154046 43494 154102
rect 42874 153978 43494 154046
rect 42874 153922 42970 153978
rect 43026 153922 43094 153978
rect 43150 153922 43218 153978
rect 43274 153922 43342 153978
rect 43398 153922 43494 153978
rect 42874 136350 43494 153922
rect 42874 136294 42970 136350
rect 43026 136294 43094 136350
rect 43150 136294 43218 136350
rect 43274 136294 43342 136350
rect 43398 136294 43494 136350
rect 42874 136226 43494 136294
rect 42874 136170 42970 136226
rect 43026 136170 43094 136226
rect 43150 136170 43218 136226
rect 43274 136170 43342 136226
rect 43398 136170 43494 136226
rect 42874 136102 43494 136170
rect 42874 136046 42970 136102
rect 43026 136046 43094 136102
rect 43150 136046 43218 136102
rect 43274 136046 43342 136102
rect 43398 136046 43494 136102
rect 42874 135978 43494 136046
rect 42874 135922 42970 135978
rect 43026 135922 43094 135978
rect 43150 135922 43218 135978
rect 43274 135922 43342 135978
rect 43398 135922 43494 135978
rect 42874 118350 43494 135922
rect 42874 118294 42970 118350
rect 43026 118294 43094 118350
rect 43150 118294 43218 118350
rect 43274 118294 43342 118350
rect 43398 118294 43494 118350
rect 42874 118226 43494 118294
rect 42874 118170 42970 118226
rect 43026 118170 43094 118226
rect 43150 118170 43218 118226
rect 43274 118170 43342 118226
rect 43398 118170 43494 118226
rect 42874 118102 43494 118170
rect 42874 118046 42970 118102
rect 43026 118046 43094 118102
rect 43150 118046 43218 118102
rect 43274 118046 43342 118102
rect 43398 118046 43494 118102
rect 42874 117978 43494 118046
rect 42874 117922 42970 117978
rect 43026 117922 43094 117978
rect 43150 117922 43218 117978
rect 43274 117922 43342 117978
rect 43398 117922 43494 117978
rect 42874 100350 43494 117922
rect 57154 148350 57774 158858
rect 57154 148294 57250 148350
rect 57306 148294 57374 148350
rect 57430 148294 57498 148350
rect 57554 148294 57622 148350
rect 57678 148294 57774 148350
rect 57154 148226 57774 148294
rect 57154 148170 57250 148226
rect 57306 148170 57374 148226
rect 57430 148170 57498 148226
rect 57554 148170 57622 148226
rect 57678 148170 57774 148226
rect 57154 148102 57774 148170
rect 57154 148046 57250 148102
rect 57306 148046 57374 148102
rect 57430 148046 57498 148102
rect 57554 148046 57622 148102
rect 57678 148046 57774 148102
rect 57154 147978 57774 148046
rect 57154 147922 57250 147978
rect 57306 147922 57374 147978
rect 57430 147922 57498 147978
rect 57554 147922 57622 147978
rect 57678 147922 57774 147978
rect 57154 130350 57774 147922
rect 57154 130294 57250 130350
rect 57306 130294 57374 130350
rect 57430 130294 57498 130350
rect 57554 130294 57622 130350
rect 57678 130294 57774 130350
rect 57154 130226 57774 130294
rect 57154 130170 57250 130226
rect 57306 130170 57374 130226
rect 57430 130170 57498 130226
rect 57554 130170 57622 130226
rect 57678 130170 57774 130226
rect 57154 130102 57774 130170
rect 57154 130046 57250 130102
rect 57306 130046 57374 130102
rect 57430 130046 57498 130102
rect 57554 130046 57622 130102
rect 57678 130046 57774 130102
rect 57154 129978 57774 130046
rect 57154 129922 57250 129978
rect 57306 129922 57374 129978
rect 57430 129922 57498 129978
rect 57554 129922 57622 129978
rect 57678 129922 57774 129978
rect 57154 112350 57774 129922
rect 57154 112294 57250 112350
rect 57306 112294 57374 112350
rect 57430 112294 57498 112350
rect 57554 112294 57622 112350
rect 57678 112294 57774 112350
rect 57154 112226 57774 112294
rect 57154 112170 57250 112226
rect 57306 112170 57374 112226
rect 57430 112170 57498 112226
rect 57554 112170 57622 112226
rect 57678 112170 57774 112226
rect 57154 112102 57774 112170
rect 57154 112046 57250 112102
rect 57306 112046 57374 112102
rect 57430 112046 57498 112102
rect 57554 112046 57622 112102
rect 57678 112046 57774 112102
rect 57154 111978 57774 112046
rect 57154 111922 57250 111978
rect 57306 111922 57374 111978
rect 57430 111922 57498 111978
rect 57554 111922 57622 111978
rect 57678 111922 57774 111978
rect 57154 111238 57774 111922
rect 60874 154350 61494 158858
rect 60874 154294 60970 154350
rect 61026 154294 61094 154350
rect 61150 154294 61218 154350
rect 61274 154294 61342 154350
rect 61398 154294 61494 154350
rect 60874 154226 61494 154294
rect 60874 154170 60970 154226
rect 61026 154170 61094 154226
rect 61150 154170 61218 154226
rect 61274 154170 61342 154226
rect 61398 154170 61494 154226
rect 60874 154102 61494 154170
rect 60874 154046 60970 154102
rect 61026 154046 61094 154102
rect 61150 154046 61218 154102
rect 61274 154046 61342 154102
rect 61398 154046 61494 154102
rect 60874 153978 61494 154046
rect 60874 153922 60970 153978
rect 61026 153922 61094 153978
rect 61150 153922 61218 153978
rect 61274 153922 61342 153978
rect 61398 153922 61494 153978
rect 60874 136350 61494 153922
rect 60874 136294 60970 136350
rect 61026 136294 61094 136350
rect 61150 136294 61218 136350
rect 61274 136294 61342 136350
rect 61398 136294 61494 136350
rect 60874 136226 61494 136294
rect 60874 136170 60970 136226
rect 61026 136170 61094 136226
rect 61150 136170 61218 136226
rect 61274 136170 61342 136226
rect 61398 136170 61494 136226
rect 60874 136102 61494 136170
rect 60874 136046 60970 136102
rect 61026 136046 61094 136102
rect 61150 136046 61218 136102
rect 61274 136046 61342 136102
rect 61398 136046 61494 136102
rect 60874 135978 61494 136046
rect 60874 135922 60970 135978
rect 61026 135922 61094 135978
rect 61150 135922 61218 135978
rect 61274 135922 61342 135978
rect 61398 135922 61494 135978
rect 60874 118350 61494 135922
rect 60874 118294 60970 118350
rect 61026 118294 61094 118350
rect 61150 118294 61218 118350
rect 61274 118294 61342 118350
rect 61398 118294 61494 118350
rect 60874 118226 61494 118294
rect 60874 118170 60970 118226
rect 61026 118170 61094 118226
rect 61150 118170 61218 118226
rect 61274 118170 61342 118226
rect 61398 118170 61494 118226
rect 60874 118102 61494 118170
rect 60874 118046 60970 118102
rect 61026 118046 61094 118102
rect 61150 118046 61218 118102
rect 61274 118046 61342 118102
rect 61398 118046 61494 118102
rect 60874 117978 61494 118046
rect 60874 117922 60970 117978
rect 61026 117922 61094 117978
rect 61150 117922 61218 117978
rect 61274 117922 61342 117978
rect 61398 117922 61494 117978
rect 60874 111238 61494 117922
rect 75154 148350 75774 158858
rect 75154 148294 75250 148350
rect 75306 148294 75374 148350
rect 75430 148294 75498 148350
rect 75554 148294 75622 148350
rect 75678 148294 75774 148350
rect 75154 148226 75774 148294
rect 75154 148170 75250 148226
rect 75306 148170 75374 148226
rect 75430 148170 75498 148226
rect 75554 148170 75622 148226
rect 75678 148170 75774 148226
rect 75154 148102 75774 148170
rect 75154 148046 75250 148102
rect 75306 148046 75374 148102
rect 75430 148046 75498 148102
rect 75554 148046 75622 148102
rect 75678 148046 75774 148102
rect 75154 147978 75774 148046
rect 75154 147922 75250 147978
rect 75306 147922 75374 147978
rect 75430 147922 75498 147978
rect 75554 147922 75622 147978
rect 75678 147922 75774 147978
rect 75154 130350 75774 147922
rect 75154 130294 75250 130350
rect 75306 130294 75374 130350
rect 75430 130294 75498 130350
rect 75554 130294 75622 130350
rect 75678 130294 75774 130350
rect 75154 130226 75774 130294
rect 75154 130170 75250 130226
rect 75306 130170 75374 130226
rect 75430 130170 75498 130226
rect 75554 130170 75622 130226
rect 75678 130170 75774 130226
rect 75154 130102 75774 130170
rect 75154 130046 75250 130102
rect 75306 130046 75374 130102
rect 75430 130046 75498 130102
rect 75554 130046 75622 130102
rect 75678 130046 75774 130102
rect 75154 129978 75774 130046
rect 75154 129922 75250 129978
rect 75306 129922 75374 129978
rect 75430 129922 75498 129978
rect 75554 129922 75622 129978
rect 75678 129922 75774 129978
rect 75154 112350 75774 129922
rect 75154 112294 75250 112350
rect 75306 112294 75374 112350
rect 75430 112294 75498 112350
rect 75554 112294 75622 112350
rect 75678 112294 75774 112350
rect 75154 112226 75774 112294
rect 75154 112170 75250 112226
rect 75306 112170 75374 112226
rect 75430 112170 75498 112226
rect 75554 112170 75622 112226
rect 75678 112170 75774 112226
rect 75154 112102 75774 112170
rect 75154 112046 75250 112102
rect 75306 112046 75374 112102
rect 75430 112046 75498 112102
rect 75554 112046 75622 112102
rect 75678 112046 75774 112102
rect 75154 111978 75774 112046
rect 75154 111922 75250 111978
rect 75306 111922 75374 111978
rect 75430 111922 75498 111978
rect 75554 111922 75622 111978
rect 75678 111922 75774 111978
rect 75154 111238 75774 111922
rect 78874 154350 79494 158858
rect 78874 154294 78970 154350
rect 79026 154294 79094 154350
rect 79150 154294 79218 154350
rect 79274 154294 79342 154350
rect 79398 154294 79494 154350
rect 78874 154226 79494 154294
rect 78874 154170 78970 154226
rect 79026 154170 79094 154226
rect 79150 154170 79218 154226
rect 79274 154170 79342 154226
rect 79398 154170 79494 154226
rect 78874 154102 79494 154170
rect 78874 154046 78970 154102
rect 79026 154046 79094 154102
rect 79150 154046 79218 154102
rect 79274 154046 79342 154102
rect 79398 154046 79494 154102
rect 78874 153978 79494 154046
rect 78874 153922 78970 153978
rect 79026 153922 79094 153978
rect 79150 153922 79218 153978
rect 79274 153922 79342 153978
rect 79398 153922 79494 153978
rect 78874 136350 79494 153922
rect 78874 136294 78970 136350
rect 79026 136294 79094 136350
rect 79150 136294 79218 136350
rect 79274 136294 79342 136350
rect 79398 136294 79494 136350
rect 78874 136226 79494 136294
rect 78874 136170 78970 136226
rect 79026 136170 79094 136226
rect 79150 136170 79218 136226
rect 79274 136170 79342 136226
rect 79398 136170 79494 136226
rect 78874 136102 79494 136170
rect 78874 136046 78970 136102
rect 79026 136046 79094 136102
rect 79150 136046 79218 136102
rect 79274 136046 79342 136102
rect 79398 136046 79494 136102
rect 78874 135978 79494 136046
rect 78874 135922 78970 135978
rect 79026 135922 79094 135978
rect 79150 135922 79218 135978
rect 79274 135922 79342 135978
rect 79398 135922 79494 135978
rect 78874 118350 79494 135922
rect 78874 118294 78970 118350
rect 79026 118294 79094 118350
rect 79150 118294 79218 118350
rect 79274 118294 79342 118350
rect 79398 118294 79494 118350
rect 78874 118226 79494 118294
rect 78874 118170 78970 118226
rect 79026 118170 79094 118226
rect 79150 118170 79218 118226
rect 79274 118170 79342 118226
rect 79398 118170 79494 118226
rect 78874 118102 79494 118170
rect 78874 118046 78970 118102
rect 79026 118046 79094 118102
rect 79150 118046 79218 118102
rect 79274 118046 79342 118102
rect 79398 118046 79494 118102
rect 78874 117978 79494 118046
rect 78874 117922 78970 117978
rect 79026 117922 79094 117978
rect 79150 117922 79218 117978
rect 79274 117922 79342 117978
rect 79398 117922 79494 117978
rect 78874 111238 79494 117922
rect 93154 148350 93774 158858
rect 93154 148294 93250 148350
rect 93306 148294 93374 148350
rect 93430 148294 93498 148350
rect 93554 148294 93622 148350
rect 93678 148294 93774 148350
rect 93154 148226 93774 148294
rect 93154 148170 93250 148226
rect 93306 148170 93374 148226
rect 93430 148170 93498 148226
rect 93554 148170 93622 148226
rect 93678 148170 93774 148226
rect 93154 148102 93774 148170
rect 93154 148046 93250 148102
rect 93306 148046 93374 148102
rect 93430 148046 93498 148102
rect 93554 148046 93622 148102
rect 93678 148046 93774 148102
rect 93154 147978 93774 148046
rect 93154 147922 93250 147978
rect 93306 147922 93374 147978
rect 93430 147922 93498 147978
rect 93554 147922 93622 147978
rect 93678 147922 93774 147978
rect 93154 130350 93774 147922
rect 93154 130294 93250 130350
rect 93306 130294 93374 130350
rect 93430 130294 93498 130350
rect 93554 130294 93622 130350
rect 93678 130294 93774 130350
rect 93154 130226 93774 130294
rect 93154 130170 93250 130226
rect 93306 130170 93374 130226
rect 93430 130170 93498 130226
rect 93554 130170 93622 130226
rect 93678 130170 93774 130226
rect 93154 130102 93774 130170
rect 93154 130046 93250 130102
rect 93306 130046 93374 130102
rect 93430 130046 93498 130102
rect 93554 130046 93622 130102
rect 93678 130046 93774 130102
rect 93154 129978 93774 130046
rect 93154 129922 93250 129978
rect 93306 129922 93374 129978
rect 93430 129922 93498 129978
rect 93554 129922 93622 129978
rect 93678 129922 93774 129978
rect 93154 112350 93774 129922
rect 93154 112294 93250 112350
rect 93306 112294 93374 112350
rect 93430 112294 93498 112350
rect 93554 112294 93622 112350
rect 93678 112294 93774 112350
rect 93154 112226 93774 112294
rect 93154 112170 93250 112226
rect 93306 112170 93374 112226
rect 93430 112170 93498 112226
rect 93554 112170 93622 112226
rect 93678 112170 93774 112226
rect 93154 112102 93774 112170
rect 93154 112046 93250 112102
rect 93306 112046 93374 112102
rect 93430 112046 93498 112102
rect 93554 112046 93622 112102
rect 93678 112046 93774 112102
rect 93154 111978 93774 112046
rect 93154 111922 93250 111978
rect 93306 111922 93374 111978
rect 93430 111922 93498 111978
rect 93554 111922 93622 111978
rect 93678 111922 93774 111978
rect 93154 111238 93774 111922
rect 96874 154350 97494 158858
rect 96874 154294 96970 154350
rect 97026 154294 97094 154350
rect 97150 154294 97218 154350
rect 97274 154294 97342 154350
rect 97398 154294 97494 154350
rect 96874 154226 97494 154294
rect 96874 154170 96970 154226
rect 97026 154170 97094 154226
rect 97150 154170 97218 154226
rect 97274 154170 97342 154226
rect 97398 154170 97494 154226
rect 96874 154102 97494 154170
rect 96874 154046 96970 154102
rect 97026 154046 97094 154102
rect 97150 154046 97218 154102
rect 97274 154046 97342 154102
rect 97398 154046 97494 154102
rect 96874 153978 97494 154046
rect 96874 153922 96970 153978
rect 97026 153922 97094 153978
rect 97150 153922 97218 153978
rect 97274 153922 97342 153978
rect 97398 153922 97494 153978
rect 96874 136350 97494 153922
rect 96874 136294 96970 136350
rect 97026 136294 97094 136350
rect 97150 136294 97218 136350
rect 97274 136294 97342 136350
rect 97398 136294 97494 136350
rect 96874 136226 97494 136294
rect 96874 136170 96970 136226
rect 97026 136170 97094 136226
rect 97150 136170 97218 136226
rect 97274 136170 97342 136226
rect 97398 136170 97494 136226
rect 96874 136102 97494 136170
rect 96874 136046 96970 136102
rect 97026 136046 97094 136102
rect 97150 136046 97218 136102
rect 97274 136046 97342 136102
rect 97398 136046 97494 136102
rect 96874 135978 97494 136046
rect 96874 135922 96970 135978
rect 97026 135922 97094 135978
rect 97150 135922 97218 135978
rect 97274 135922 97342 135978
rect 97398 135922 97494 135978
rect 96874 118350 97494 135922
rect 96874 118294 96970 118350
rect 97026 118294 97094 118350
rect 97150 118294 97218 118350
rect 97274 118294 97342 118350
rect 97398 118294 97494 118350
rect 96874 118226 97494 118294
rect 96874 118170 96970 118226
rect 97026 118170 97094 118226
rect 97150 118170 97218 118226
rect 97274 118170 97342 118226
rect 97398 118170 97494 118226
rect 96874 118102 97494 118170
rect 96874 118046 96970 118102
rect 97026 118046 97094 118102
rect 97150 118046 97218 118102
rect 97274 118046 97342 118102
rect 97398 118046 97494 118102
rect 96874 117978 97494 118046
rect 96874 117922 96970 117978
rect 97026 117922 97094 117978
rect 97150 117922 97218 117978
rect 97274 117922 97342 117978
rect 97398 117922 97494 117978
rect 96874 111238 97494 117922
rect 111154 148350 111774 158858
rect 111154 148294 111250 148350
rect 111306 148294 111374 148350
rect 111430 148294 111498 148350
rect 111554 148294 111622 148350
rect 111678 148294 111774 148350
rect 111154 148226 111774 148294
rect 111154 148170 111250 148226
rect 111306 148170 111374 148226
rect 111430 148170 111498 148226
rect 111554 148170 111622 148226
rect 111678 148170 111774 148226
rect 111154 148102 111774 148170
rect 111154 148046 111250 148102
rect 111306 148046 111374 148102
rect 111430 148046 111498 148102
rect 111554 148046 111622 148102
rect 111678 148046 111774 148102
rect 111154 147978 111774 148046
rect 111154 147922 111250 147978
rect 111306 147922 111374 147978
rect 111430 147922 111498 147978
rect 111554 147922 111622 147978
rect 111678 147922 111774 147978
rect 111154 130350 111774 147922
rect 111154 130294 111250 130350
rect 111306 130294 111374 130350
rect 111430 130294 111498 130350
rect 111554 130294 111622 130350
rect 111678 130294 111774 130350
rect 111154 130226 111774 130294
rect 111154 130170 111250 130226
rect 111306 130170 111374 130226
rect 111430 130170 111498 130226
rect 111554 130170 111622 130226
rect 111678 130170 111774 130226
rect 111154 130102 111774 130170
rect 111154 130046 111250 130102
rect 111306 130046 111374 130102
rect 111430 130046 111498 130102
rect 111554 130046 111622 130102
rect 111678 130046 111774 130102
rect 111154 129978 111774 130046
rect 111154 129922 111250 129978
rect 111306 129922 111374 129978
rect 111430 129922 111498 129978
rect 111554 129922 111622 129978
rect 111678 129922 111774 129978
rect 111154 112350 111774 129922
rect 111154 112294 111250 112350
rect 111306 112294 111374 112350
rect 111430 112294 111498 112350
rect 111554 112294 111622 112350
rect 111678 112294 111774 112350
rect 111154 112226 111774 112294
rect 111154 112170 111250 112226
rect 111306 112170 111374 112226
rect 111430 112170 111498 112226
rect 111554 112170 111622 112226
rect 111678 112170 111774 112226
rect 111154 112102 111774 112170
rect 111154 112046 111250 112102
rect 111306 112046 111374 112102
rect 111430 112046 111498 112102
rect 111554 112046 111622 112102
rect 111678 112046 111774 112102
rect 111154 111978 111774 112046
rect 111154 111922 111250 111978
rect 111306 111922 111374 111978
rect 111430 111922 111498 111978
rect 111554 111922 111622 111978
rect 111678 111922 111774 111978
rect 111154 111238 111774 111922
rect 114874 154350 115494 158858
rect 114874 154294 114970 154350
rect 115026 154294 115094 154350
rect 115150 154294 115218 154350
rect 115274 154294 115342 154350
rect 115398 154294 115494 154350
rect 114874 154226 115494 154294
rect 114874 154170 114970 154226
rect 115026 154170 115094 154226
rect 115150 154170 115218 154226
rect 115274 154170 115342 154226
rect 115398 154170 115494 154226
rect 114874 154102 115494 154170
rect 114874 154046 114970 154102
rect 115026 154046 115094 154102
rect 115150 154046 115218 154102
rect 115274 154046 115342 154102
rect 115398 154046 115494 154102
rect 114874 153978 115494 154046
rect 114874 153922 114970 153978
rect 115026 153922 115094 153978
rect 115150 153922 115218 153978
rect 115274 153922 115342 153978
rect 115398 153922 115494 153978
rect 114874 136350 115494 153922
rect 114874 136294 114970 136350
rect 115026 136294 115094 136350
rect 115150 136294 115218 136350
rect 115274 136294 115342 136350
rect 115398 136294 115494 136350
rect 114874 136226 115494 136294
rect 114874 136170 114970 136226
rect 115026 136170 115094 136226
rect 115150 136170 115218 136226
rect 115274 136170 115342 136226
rect 115398 136170 115494 136226
rect 114874 136102 115494 136170
rect 114874 136046 114970 136102
rect 115026 136046 115094 136102
rect 115150 136046 115218 136102
rect 115274 136046 115342 136102
rect 115398 136046 115494 136102
rect 114874 135978 115494 136046
rect 114874 135922 114970 135978
rect 115026 135922 115094 135978
rect 115150 135922 115218 135978
rect 115274 135922 115342 135978
rect 115398 135922 115494 135978
rect 114874 118350 115494 135922
rect 114874 118294 114970 118350
rect 115026 118294 115094 118350
rect 115150 118294 115218 118350
rect 115274 118294 115342 118350
rect 115398 118294 115494 118350
rect 114874 118226 115494 118294
rect 114874 118170 114970 118226
rect 115026 118170 115094 118226
rect 115150 118170 115218 118226
rect 115274 118170 115342 118226
rect 115398 118170 115494 118226
rect 114874 118102 115494 118170
rect 114874 118046 114970 118102
rect 115026 118046 115094 118102
rect 115150 118046 115218 118102
rect 115274 118046 115342 118102
rect 115398 118046 115494 118102
rect 114874 117978 115494 118046
rect 114874 117922 114970 117978
rect 115026 117922 115094 117978
rect 115150 117922 115218 117978
rect 115274 117922 115342 117978
rect 115398 117922 115494 117978
rect 114874 111238 115494 117922
rect 129154 148350 129774 158858
rect 129154 148294 129250 148350
rect 129306 148294 129374 148350
rect 129430 148294 129498 148350
rect 129554 148294 129622 148350
rect 129678 148294 129774 148350
rect 129154 148226 129774 148294
rect 129154 148170 129250 148226
rect 129306 148170 129374 148226
rect 129430 148170 129498 148226
rect 129554 148170 129622 148226
rect 129678 148170 129774 148226
rect 129154 148102 129774 148170
rect 129154 148046 129250 148102
rect 129306 148046 129374 148102
rect 129430 148046 129498 148102
rect 129554 148046 129622 148102
rect 129678 148046 129774 148102
rect 129154 147978 129774 148046
rect 129154 147922 129250 147978
rect 129306 147922 129374 147978
rect 129430 147922 129498 147978
rect 129554 147922 129622 147978
rect 129678 147922 129774 147978
rect 129154 130350 129774 147922
rect 129154 130294 129250 130350
rect 129306 130294 129374 130350
rect 129430 130294 129498 130350
rect 129554 130294 129622 130350
rect 129678 130294 129774 130350
rect 129154 130226 129774 130294
rect 129154 130170 129250 130226
rect 129306 130170 129374 130226
rect 129430 130170 129498 130226
rect 129554 130170 129622 130226
rect 129678 130170 129774 130226
rect 129154 130102 129774 130170
rect 129154 130046 129250 130102
rect 129306 130046 129374 130102
rect 129430 130046 129498 130102
rect 129554 130046 129622 130102
rect 129678 130046 129774 130102
rect 129154 129978 129774 130046
rect 129154 129922 129250 129978
rect 129306 129922 129374 129978
rect 129430 129922 129498 129978
rect 129554 129922 129622 129978
rect 129678 129922 129774 129978
rect 129154 112350 129774 129922
rect 129154 112294 129250 112350
rect 129306 112294 129374 112350
rect 129430 112294 129498 112350
rect 129554 112294 129622 112350
rect 129678 112294 129774 112350
rect 129154 112226 129774 112294
rect 129154 112170 129250 112226
rect 129306 112170 129374 112226
rect 129430 112170 129498 112226
rect 129554 112170 129622 112226
rect 129678 112170 129774 112226
rect 129154 112102 129774 112170
rect 129154 112046 129250 112102
rect 129306 112046 129374 112102
rect 129430 112046 129498 112102
rect 129554 112046 129622 112102
rect 129678 112046 129774 112102
rect 129154 111978 129774 112046
rect 129154 111922 129250 111978
rect 129306 111922 129374 111978
rect 129430 111922 129498 111978
rect 129554 111922 129622 111978
rect 129678 111922 129774 111978
rect 129154 111238 129774 111922
rect 132874 154350 133494 158858
rect 132874 154294 132970 154350
rect 133026 154294 133094 154350
rect 133150 154294 133218 154350
rect 133274 154294 133342 154350
rect 133398 154294 133494 154350
rect 132874 154226 133494 154294
rect 132874 154170 132970 154226
rect 133026 154170 133094 154226
rect 133150 154170 133218 154226
rect 133274 154170 133342 154226
rect 133398 154170 133494 154226
rect 132874 154102 133494 154170
rect 132874 154046 132970 154102
rect 133026 154046 133094 154102
rect 133150 154046 133218 154102
rect 133274 154046 133342 154102
rect 133398 154046 133494 154102
rect 132874 153978 133494 154046
rect 132874 153922 132970 153978
rect 133026 153922 133094 153978
rect 133150 153922 133218 153978
rect 133274 153922 133342 153978
rect 133398 153922 133494 153978
rect 132874 136350 133494 153922
rect 132874 136294 132970 136350
rect 133026 136294 133094 136350
rect 133150 136294 133218 136350
rect 133274 136294 133342 136350
rect 133398 136294 133494 136350
rect 132874 136226 133494 136294
rect 132874 136170 132970 136226
rect 133026 136170 133094 136226
rect 133150 136170 133218 136226
rect 133274 136170 133342 136226
rect 133398 136170 133494 136226
rect 132874 136102 133494 136170
rect 132874 136046 132970 136102
rect 133026 136046 133094 136102
rect 133150 136046 133218 136102
rect 133274 136046 133342 136102
rect 133398 136046 133494 136102
rect 132874 135978 133494 136046
rect 132874 135922 132970 135978
rect 133026 135922 133094 135978
rect 133150 135922 133218 135978
rect 133274 135922 133342 135978
rect 133398 135922 133494 135978
rect 132874 118350 133494 135922
rect 132874 118294 132970 118350
rect 133026 118294 133094 118350
rect 133150 118294 133218 118350
rect 133274 118294 133342 118350
rect 133398 118294 133494 118350
rect 132874 118226 133494 118294
rect 132874 118170 132970 118226
rect 133026 118170 133094 118226
rect 133150 118170 133218 118226
rect 133274 118170 133342 118226
rect 133398 118170 133494 118226
rect 132874 118102 133494 118170
rect 132874 118046 132970 118102
rect 133026 118046 133094 118102
rect 133150 118046 133218 118102
rect 133274 118046 133342 118102
rect 133398 118046 133494 118102
rect 132874 117978 133494 118046
rect 132874 117922 132970 117978
rect 133026 117922 133094 117978
rect 133150 117922 133218 117978
rect 133274 117922 133342 117978
rect 133398 117922 133494 117978
rect 132874 111238 133494 117922
rect 147154 148350 147774 158858
rect 147154 148294 147250 148350
rect 147306 148294 147374 148350
rect 147430 148294 147498 148350
rect 147554 148294 147622 148350
rect 147678 148294 147774 148350
rect 147154 148226 147774 148294
rect 147154 148170 147250 148226
rect 147306 148170 147374 148226
rect 147430 148170 147498 148226
rect 147554 148170 147622 148226
rect 147678 148170 147774 148226
rect 147154 148102 147774 148170
rect 147154 148046 147250 148102
rect 147306 148046 147374 148102
rect 147430 148046 147498 148102
rect 147554 148046 147622 148102
rect 147678 148046 147774 148102
rect 147154 147978 147774 148046
rect 147154 147922 147250 147978
rect 147306 147922 147374 147978
rect 147430 147922 147498 147978
rect 147554 147922 147622 147978
rect 147678 147922 147774 147978
rect 147154 130350 147774 147922
rect 147154 130294 147250 130350
rect 147306 130294 147374 130350
rect 147430 130294 147498 130350
rect 147554 130294 147622 130350
rect 147678 130294 147774 130350
rect 147154 130226 147774 130294
rect 147154 130170 147250 130226
rect 147306 130170 147374 130226
rect 147430 130170 147498 130226
rect 147554 130170 147622 130226
rect 147678 130170 147774 130226
rect 147154 130102 147774 130170
rect 147154 130046 147250 130102
rect 147306 130046 147374 130102
rect 147430 130046 147498 130102
rect 147554 130046 147622 130102
rect 147678 130046 147774 130102
rect 147154 129978 147774 130046
rect 147154 129922 147250 129978
rect 147306 129922 147374 129978
rect 147430 129922 147498 129978
rect 147554 129922 147622 129978
rect 147678 129922 147774 129978
rect 147154 112350 147774 129922
rect 147154 112294 147250 112350
rect 147306 112294 147374 112350
rect 147430 112294 147498 112350
rect 147554 112294 147622 112350
rect 147678 112294 147774 112350
rect 147154 112226 147774 112294
rect 147154 112170 147250 112226
rect 147306 112170 147374 112226
rect 147430 112170 147498 112226
rect 147554 112170 147622 112226
rect 147678 112170 147774 112226
rect 147154 112102 147774 112170
rect 147154 112046 147250 112102
rect 147306 112046 147374 112102
rect 147430 112046 147498 112102
rect 147554 112046 147622 112102
rect 147678 112046 147774 112102
rect 147154 111978 147774 112046
rect 147154 111922 147250 111978
rect 147306 111922 147374 111978
rect 147430 111922 147498 111978
rect 147554 111922 147622 111978
rect 147678 111922 147774 111978
rect 147154 111238 147774 111922
rect 150874 154350 151494 158858
rect 150874 154294 150970 154350
rect 151026 154294 151094 154350
rect 151150 154294 151218 154350
rect 151274 154294 151342 154350
rect 151398 154294 151494 154350
rect 150874 154226 151494 154294
rect 150874 154170 150970 154226
rect 151026 154170 151094 154226
rect 151150 154170 151218 154226
rect 151274 154170 151342 154226
rect 151398 154170 151494 154226
rect 150874 154102 151494 154170
rect 150874 154046 150970 154102
rect 151026 154046 151094 154102
rect 151150 154046 151218 154102
rect 151274 154046 151342 154102
rect 151398 154046 151494 154102
rect 150874 153978 151494 154046
rect 150874 153922 150970 153978
rect 151026 153922 151094 153978
rect 151150 153922 151218 153978
rect 151274 153922 151342 153978
rect 151398 153922 151494 153978
rect 150874 136350 151494 153922
rect 150874 136294 150970 136350
rect 151026 136294 151094 136350
rect 151150 136294 151218 136350
rect 151274 136294 151342 136350
rect 151398 136294 151494 136350
rect 150874 136226 151494 136294
rect 150874 136170 150970 136226
rect 151026 136170 151094 136226
rect 151150 136170 151218 136226
rect 151274 136170 151342 136226
rect 151398 136170 151494 136226
rect 150874 136102 151494 136170
rect 150874 136046 150970 136102
rect 151026 136046 151094 136102
rect 151150 136046 151218 136102
rect 151274 136046 151342 136102
rect 151398 136046 151494 136102
rect 150874 135978 151494 136046
rect 150874 135922 150970 135978
rect 151026 135922 151094 135978
rect 151150 135922 151218 135978
rect 151274 135922 151342 135978
rect 151398 135922 151494 135978
rect 150874 118350 151494 135922
rect 150874 118294 150970 118350
rect 151026 118294 151094 118350
rect 151150 118294 151218 118350
rect 151274 118294 151342 118350
rect 151398 118294 151494 118350
rect 150874 118226 151494 118294
rect 150874 118170 150970 118226
rect 151026 118170 151094 118226
rect 151150 118170 151218 118226
rect 151274 118170 151342 118226
rect 151398 118170 151494 118226
rect 150874 118102 151494 118170
rect 150874 118046 150970 118102
rect 151026 118046 151094 118102
rect 151150 118046 151218 118102
rect 151274 118046 151342 118102
rect 151398 118046 151494 118102
rect 150874 117978 151494 118046
rect 150874 117922 150970 117978
rect 151026 117922 151094 117978
rect 151150 117922 151218 117978
rect 151274 117922 151342 117978
rect 151398 117922 151494 117978
rect 150874 111238 151494 117922
rect 165154 148350 165774 158858
rect 165154 148294 165250 148350
rect 165306 148294 165374 148350
rect 165430 148294 165498 148350
rect 165554 148294 165622 148350
rect 165678 148294 165774 148350
rect 165154 148226 165774 148294
rect 165154 148170 165250 148226
rect 165306 148170 165374 148226
rect 165430 148170 165498 148226
rect 165554 148170 165622 148226
rect 165678 148170 165774 148226
rect 165154 148102 165774 148170
rect 165154 148046 165250 148102
rect 165306 148046 165374 148102
rect 165430 148046 165498 148102
rect 165554 148046 165622 148102
rect 165678 148046 165774 148102
rect 165154 147978 165774 148046
rect 165154 147922 165250 147978
rect 165306 147922 165374 147978
rect 165430 147922 165498 147978
rect 165554 147922 165622 147978
rect 165678 147922 165774 147978
rect 165154 130350 165774 147922
rect 165154 130294 165250 130350
rect 165306 130294 165374 130350
rect 165430 130294 165498 130350
rect 165554 130294 165622 130350
rect 165678 130294 165774 130350
rect 165154 130226 165774 130294
rect 165154 130170 165250 130226
rect 165306 130170 165374 130226
rect 165430 130170 165498 130226
rect 165554 130170 165622 130226
rect 165678 130170 165774 130226
rect 165154 130102 165774 130170
rect 165154 130046 165250 130102
rect 165306 130046 165374 130102
rect 165430 130046 165498 130102
rect 165554 130046 165622 130102
rect 165678 130046 165774 130102
rect 165154 129978 165774 130046
rect 165154 129922 165250 129978
rect 165306 129922 165374 129978
rect 165430 129922 165498 129978
rect 165554 129922 165622 129978
rect 165678 129922 165774 129978
rect 165154 112350 165774 129922
rect 165154 112294 165250 112350
rect 165306 112294 165374 112350
rect 165430 112294 165498 112350
rect 165554 112294 165622 112350
rect 165678 112294 165774 112350
rect 165154 112226 165774 112294
rect 165154 112170 165250 112226
rect 165306 112170 165374 112226
rect 165430 112170 165498 112226
rect 165554 112170 165622 112226
rect 165678 112170 165774 112226
rect 165154 112102 165774 112170
rect 165154 112046 165250 112102
rect 165306 112046 165374 112102
rect 165430 112046 165498 112102
rect 165554 112046 165622 112102
rect 165678 112046 165774 112102
rect 165154 111978 165774 112046
rect 165154 111922 165250 111978
rect 165306 111922 165374 111978
rect 165430 111922 165498 111978
rect 165554 111922 165622 111978
rect 165678 111922 165774 111978
rect 165154 111238 165774 111922
rect 168874 154350 169494 158858
rect 168874 154294 168970 154350
rect 169026 154294 169094 154350
rect 169150 154294 169218 154350
rect 169274 154294 169342 154350
rect 169398 154294 169494 154350
rect 168874 154226 169494 154294
rect 168874 154170 168970 154226
rect 169026 154170 169094 154226
rect 169150 154170 169218 154226
rect 169274 154170 169342 154226
rect 169398 154170 169494 154226
rect 168874 154102 169494 154170
rect 168874 154046 168970 154102
rect 169026 154046 169094 154102
rect 169150 154046 169218 154102
rect 169274 154046 169342 154102
rect 169398 154046 169494 154102
rect 168874 153978 169494 154046
rect 168874 153922 168970 153978
rect 169026 153922 169094 153978
rect 169150 153922 169218 153978
rect 169274 153922 169342 153978
rect 169398 153922 169494 153978
rect 168874 136350 169494 153922
rect 168874 136294 168970 136350
rect 169026 136294 169094 136350
rect 169150 136294 169218 136350
rect 169274 136294 169342 136350
rect 169398 136294 169494 136350
rect 168874 136226 169494 136294
rect 168874 136170 168970 136226
rect 169026 136170 169094 136226
rect 169150 136170 169218 136226
rect 169274 136170 169342 136226
rect 169398 136170 169494 136226
rect 168874 136102 169494 136170
rect 168874 136046 168970 136102
rect 169026 136046 169094 136102
rect 169150 136046 169218 136102
rect 169274 136046 169342 136102
rect 169398 136046 169494 136102
rect 168874 135978 169494 136046
rect 168874 135922 168970 135978
rect 169026 135922 169094 135978
rect 169150 135922 169218 135978
rect 169274 135922 169342 135978
rect 169398 135922 169494 135978
rect 168874 118350 169494 135922
rect 168874 118294 168970 118350
rect 169026 118294 169094 118350
rect 169150 118294 169218 118350
rect 169274 118294 169342 118350
rect 169398 118294 169494 118350
rect 168874 118226 169494 118294
rect 168874 118170 168970 118226
rect 169026 118170 169094 118226
rect 169150 118170 169218 118226
rect 169274 118170 169342 118226
rect 169398 118170 169494 118226
rect 168874 118102 169494 118170
rect 168874 118046 168970 118102
rect 169026 118046 169094 118102
rect 169150 118046 169218 118102
rect 169274 118046 169342 118102
rect 169398 118046 169494 118102
rect 168874 117978 169494 118046
rect 168874 117922 168970 117978
rect 169026 117922 169094 117978
rect 169150 117922 169218 117978
rect 169274 117922 169342 117978
rect 169398 117922 169494 117978
rect 168874 111238 169494 117922
rect 183154 148350 183774 158858
rect 183154 148294 183250 148350
rect 183306 148294 183374 148350
rect 183430 148294 183498 148350
rect 183554 148294 183622 148350
rect 183678 148294 183774 148350
rect 183154 148226 183774 148294
rect 183154 148170 183250 148226
rect 183306 148170 183374 148226
rect 183430 148170 183498 148226
rect 183554 148170 183622 148226
rect 183678 148170 183774 148226
rect 183154 148102 183774 148170
rect 183154 148046 183250 148102
rect 183306 148046 183374 148102
rect 183430 148046 183498 148102
rect 183554 148046 183622 148102
rect 183678 148046 183774 148102
rect 183154 147978 183774 148046
rect 183154 147922 183250 147978
rect 183306 147922 183374 147978
rect 183430 147922 183498 147978
rect 183554 147922 183622 147978
rect 183678 147922 183774 147978
rect 183154 130350 183774 147922
rect 183154 130294 183250 130350
rect 183306 130294 183374 130350
rect 183430 130294 183498 130350
rect 183554 130294 183622 130350
rect 183678 130294 183774 130350
rect 183154 130226 183774 130294
rect 183154 130170 183250 130226
rect 183306 130170 183374 130226
rect 183430 130170 183498 130226
rect 183554 130170 183622 130226
rect 183678 130170 183774 130226
rect 183154 130102 183774 130170
rect 183154 130046 183250 130102
rect 183306 130046 183374 130102
rect 183430 130046 183498 130102
rect 183554 130046 183622 130102
rect 183678 130046 183774 130102
rect 183154 129978 183774 130046
rect 183154 129922 183250 129978
rect 183306 129922 183374 129978
rect 183430 129922 183498 129978
rect 183554 129922 183622 129978
rect 183678 129922 183774 129978
rect 183154 112350 183774 129922
rect 183154 112294 183250 112350
rect 183306 112294 183374 112350
rect 183430 112294 183498 112350
rect 183554 112294 183622 112350
rect 183678 112294 183774 112350
rect 183154 112226 183774 112294
rect 183154 112170 183250 112226
rect 183306 112170 183374 112226
rect 183430 112170 183498 112226
rect 183554 112170 183622 112226
rect 183678 112170 183774 112226
rect 183154 112102 183774 112170
rect 183154 112046 183250 112102
rect 183306 112046 183374 112102
rect 183430 112046 183498 112102
rect 183554 112046 183622 112102
rect 183678 112046 183774 112102
rect 183154 111978 183774 112046
rect 183154 111922 183250 111978
rect 183306 111922 183374 111978
rect 183430 111922 183498 111978
rect 183554 111922 183622 111978
rect 183678 111922 183774 111978
rect 42874 100294 42970 100350
rect 43026 100294 43094 100350
rect 43150 100294 43218 100350
rect 43274 100294 43342 100350
rect 43398 100294 43494 100350
rect 42874 100226 43494 100294
rect 42874 100170 42970 100226
rect 43026 100170 43094 100226
rect 43150 100170 43218 100226
rect 43274 100170 43342 100226
rect 43398 100170 43494 100226
rect 42874 100102 43494 100170
rect 42874 100046 42970 100102
rect 43026 100046 43094 100102
rect 43150 100046 43218 100102
rect 43274 100046 43342 100102
rect 43398 100046 43494 100102
rect 42874 99978 43494 100046
rect 42874 99922 42970 99978
rect 43026 99922 43094 99978
rect 43150 99922 43218 99978
rect 43274 99922 43342 99978
rect 43398 99922 43494 99978
rect 42874 82350 43494 99922
rect 42874 82294 42970 82350
rect 43026 82294 43094 82350
rect 43150 82294 43218 82350
rect 43274 82294 43342 82350
rect 43398 82294 43494 82350
rect 42874 82226 43494 82294
rect 42874 82170 42970 82226
rect 43026 82170 43094 82226
rect 43150 82170 43218 82226
rect 43274 82170 43342 82226
rect 43398 82170 43494 82226
rect 42874 82102 43494 82170
rect 42874 82046 42970 82102
rect 43026 82046 43094 82102
rect 43150 82046 43218 82102
rect 43274 82046 43342 82102
rect 43398 82046 43494 82102
rect 42874 81978 43494 82046
rect 42874 81922 42970 81978
rect 43026 81922 43094 81978
rect 43150 81922 43218 81978
rect 43274 81922 43342 81978
rect 43398 81922 43494 81978
rect 39154 58294 39250 58350
rect 39306 58294 39374 58350
rect 39430 58294 39498 58350
rect 39554 58294 39622 58350
rect 39678 58294 39774 58350
rect 39154 58226 39774 58294
rect 39154 58170 39250 58226
rect 39306 58170 39374 58226
rect 39430 58170 39498 58226
rect 39554 58170 39622 58226
rect 39678 58170 39774 58226
rect 39154 58102 39774 58170
rect 39154 58046 39250 58102
rect 39306 58046 39374 58102
rect 39430 58046 39498 58102
rect 39554 58046 39622 58102
rect 39678 58046 39774 58102
rect 39154 57978 39774 58046
rect 39154 57922 39250 57978
rect 39306 57922 39374 57978
rect 39430 57922 39498 57978
rect 39554 57922 39622 57978
rect 39678 57922 39774 57978
rect 39154 40350 39774 57922
rect 39154 40294 39250 40350
rect 39306 40294 39374 40350
rect 39430 40294 39498 40350
rect 39554 40294 39622 40350
rect 39678 40294 39774 40350
rect 39154 40226 39774 40294
rect 39154 40170 39250 40226
rect 39306 40170 39374 40226
rect 39430 40170 39498 40226
rect 39554 40170 39622 40226
rect 39678 40170 39774 40226
rect 39154 40102 39774 40170
rect 39154 40046 39250 40102
rect 39306 40046 39374 40102
rect 39430 40046 39498 40102
rect 39554 40046 39622 40102
rect 39678 40046 39774 40102
rect 39154 39978 39774 40046
rect 39154 39922 39250 39978
rect 39306 39922 39374 39978
rect 39430 39922 39498 39978
rect 39554 39922 39622 39978
rect 39678 39922 39774 39978
rect 39154 22350 39774 39922
rect 39154 22294 39250 22350
rect 39306 22294 39374 22350
rect 39430 22294 39498 22350
rect 39554 22294 39622 22350
rect 39678 22294 39774 22350
rect 39154 22226 39774 22294
rect 39154 22170 39250 22226
rect 39306 22170 39374 22226
rect 39430 22170 39498 22226
rect 39554 22170 39622 22226
rect 39678 22170 39774 22226
rect 39154 22102 39774 22170
rect 39154 22046 39250 22102
rect 39306 22046 39374 22102
rect 39430 22046 39498 22102
rect 39554 22046 39622 22102
rect 39678 22046 39774 22102
rect 39154 21978 39774 22046
rect 39154 21922 39250 21978
rect 39306 21922 39374 21978
rect 39430 21922 39498 21978
rect 39554 21922 39622 21978
rect 39678 21922 39774 21978
rect 28588 6738 28644 6748
rect 24874 -1176 24970 -1120
rect 25026 -1176 25094 -1120
rect 25150 -1176 25218 -1120
rect 25274 -1176 25342 -1120
rect 25398 -1176 25494 -1120
rect 24874 -1244 25494 -1176
rect 24874 -1300 24970 -1244
rect 25026 -1300 25094 -1244
rect 25150 -1300 25218 -1244
rect 25274 -1300 25342 -1244
rect 25398 -1300 25494 -1244
rect 24874 -1368 25494 -1300
rect 24874 -1424 24970 -1368
rect 25026 -1424 25094 -1368
rect 25150 -1424 25218 -1368
rect 25274 -1424 25342 -1368
rect 25398 -1424 25494 -1368
rect 24874 -1492 25494 -1424
rect 24874 -1548 24970 -1492
rect 25026 -1548 25094 -1492
rect 25150 -1548 25218 -1492
rect 25274 -1548 25342 -1492
rect 25398 -1548 25494 -1492
rect 24874 -1644 25494 -1548
rect 39154 4350 39774 21922
rect 42028 68628 42084 68638
rect 42028 18004 42084 68572
rect 42028 17938 42084 17948
rect 42874 64350 43494 81922
rect 183154 94350 183774 111922
rect 183154 94294 183250 94350
rect 183306 94294 183374 94350
rect 183430 94294 183498 94350
rect 183554 94294 183622 94350
rect 183678 94294 183774 94350
rect 183154 94226 183774 94294
rect 183154 94170 183250 94226
rect 183306 94170 183374 94226
rect 183430 94170 183498 94226
rect 183554 94170 183622 94226
rect 183678 94170 183774 94226
rect 183154 94102 183774 94170
rect 183154 94046 183250 94102
rect 183306 94046 183374 94102
rect 183430 94046 183498 94102
rect 183554 94046 183622 94102
rect 183678 94046 183774 94102
rect 183154 93978 183774 94046
rect 183154 93922 183250 93978
rect 183306 93922 183374 93978
rect 183430 93922 183498 93978
rect 183554 93922 183622 93978
rect 183678 93922 183774 93978
rect 57154 76350 57774 77594
rect 57154 76294 57250 76350
rect 57306 76294 57374 76350
rect 57430 76294 57498 76350
rect 57554 76294 57622 76350
rect 57678 76294 57774 76350
rect 57154 76226 57774 76294
rect 57154 76170 57250 76226
rect 57306 76170 57374 76226
rect 57430 76170 57498 76226
rect 57554 76170 57622 76226
rect 57678 76170 57774 76226
rect 57154 76102 57774 76170
rect 57154 76046 57250 76102
rect 57306 76046 57374 76102
rect 57430 76046 57498 76102
rect 57554 76046 57622 76102
rect 57678 76046 57774 76102
rect 57154 75978 57774 76046
rect 57154 75922 57250 75978
rect 57306 75922 57374 75978
rect 57430 75922 57498 75978
rect 57554 75922 57622 75978
rect 57678 75922 57774 75978
rect 42874 64294 42970 64350
rect 43026 64294 43094 64350
rect 43150 64294 43218 64350
rect 43274 64294 43342 64350
rect 43398 64294 43494 64350
rect 42874 64226 43494 64294
rect 42874 64170 42970 64226
rect 43026 64170 43094 64226
rect 43150 64170 43218 64226
rect 43274 64170 43342 64226
rect 43398 64170 43494 64226
rect 42874 64102 43494 64170
rect 42874 64046 42970 64102
rect 43026 64046 43094 64102
rect 43150 64046 43218 64102
rect 43274 64046 43342 64102
rect 43398 64046 43494 64102
rect 42874 63978 43494 64046
rect 42874 63922 42970 63978
rect 43026 63922 43094 63978
rect 43150 63922 43218 63978
rect 43274 63922 43342 63978
rect 43398 63922 43494 63978
rect 42874 46350 43494 63922
rect 42874 46294 42970 46350
rect 43026 46294 43094 46350
rect 43150 46294 43218 46350
rect 43274 46294 43342 46350
rect 43398 46294 43494 46350
rect 42874 46226 43494 46294
rect 42874 46170 42970 46226
rect 43026 46170 43094 46226
rect 43150 46170 43218 46226
rect 43274 46170 43342 46226
rect 43398 46170 43494 46226
rect 42874 46102 43494 46170
rect 42874 46046 42970 46102
rect 43026 46046 43094 46102
rect 43150 46046 43218 46102
rect 43274 46046 43342 46102
rect 43398 46046 43494 46102
rect 42874 45978 43494 46046
rect 42874 45922 42970 45978
rect 43026 45922 43094 45978
rect 43150 45922 43218 45978
rect 43274 45922 43342 45978
rect 43398 45922 43494 45978
rect 42874 28350 43494 45922
rect 42874 28294 42970 28350
rect 43026 28294 43094 28350
rect 43150 28294 43218 28350
rect 43274 28294 43342 28350
rect 43398 28294 43494 28350
rect 42874 28226 43494 28294
rect 42874 28170 42970 28226
rect 43026 28170 43094 28226
rect 43150 28170 43218 28226
rect 43274 28170 43342 28226
rect 43398 28170 43494 28226
rect 42874 28102 43494 28170
rect 42874 28046 42970 28102
rect 43026 28046 43094 28102
rect 43150 28046 43218 28102
rect 43274 28046 43342 28102
rect 43398 28046 43494 28102
rect 42874 27978 43494 28046
rect 42874 27922 42970 27978
rect 43026 27922 43094 27978
rect 43150 27922 43218 27978
rect 43274 27922 43342 27978
rect 43398 27922 43494 27978
rect 39154 4294 39250 4350
rect 39306 4294 39374 4350
rect 39430 4294 39498 4350
rect 39554 4294 39622 4350
rect 39678 4294 39774 4350
rect 39154 4226 39774 4294
rect 39154 4170 39250 4226
rect 39306 4170 39374 4226
rect 39430 4170 39498 4226
rect 39554 4170 39622 4226
rect 39678 4170 39774 4226
rect 39154 4102 39774 4170
rect 39154 4046 39250 4102
rect 39306 4046 39374 4102
rect 39430 4046 39498 4102
rect 39554 4046 39622 4102
rect 39678 4046 39774 4102
rect 39154 3978 39774 4046
rect 39154 3922 39250 3978
rect 39306 3922 39374 3978
rect 39430 3922 39498 3978
rect 39554 3922 39622 3978
rect 39678 3922 39774 3978
rect 39154 -160 39774 3922
rect 39154 -216 39250 -160
rect 39306 -216 39374 -160
rect 39430 -216 39498 -160
rect 39554 -216 39622 -160
rect 39678 -216 39774 -160
rect 39154 -284 39774 -216
rect 39154 -340 39250 -284
rect 39306 -340 39374 -284
rect 39430 -340 39498 -284
rect 39554 -340 39622 -284
rect 39678 -340 39774 -284
rect 39154 -408 39774 -340
rect 39154 -464 39250 -408
rect 39306 -464 39374 -408
rect 39430 -464 39498 -408
rect 39554 -464 39622 -408
rect 39678 -464 39774 -408
rect 39154 -532 39774 -464
rect 39154 -588 39250 -532
rect 39306 -588 39374 -532
rect 39430 -588 39498 -532
rect 39554 -588 39622 -532
rect 39678 -588 39774 -532
rect 39154 -1644 39774 -588
rect 42874 10350 43494 27922
rect 48748 68628 48804 68638
rect 48748 12852 48804 68572
rect 52108 68628 52164 68638
rect 52108 16548 52164 68572
rect 53788 68628 53844 68638
rect 53788 19796 53844 68572
rect 53788 19730 53844 19740
rect 55468 68628 55524 68638
rect 55468 16772 55524 68572
rect 55468 16706 55524 16716
rect 57154 58350 57774 75922
rect 57154 58294 57250 58350
rect 57306 58294 57374 58350
rect 57430 58294 57498 58350
rect 57554 58294 57622 58350
rect 57678 58294 57774 58350
rect 57154 58226 57774 58294
rect 57154 58170 57250 58226
rect 57306 58170 57374 58226
rect 57430 58170 57498 58226
rect 57554 58170 57622 58226
rect 57678 58170 57774 58226
rect 57154 58102 57774 58170
rect 57154 58046 57250 58102
rect 57306 58046 57374 58102
rect 57430 58046 57498 58102
rect 57554 58046 57622 58102
rect 57678 58046 57774 58102
rect 57154 57978 57774 58046
rect 57154 57922 57250 57978
rect 57306 57922 57374 57978
rect 57430 57922 57498 57978
rect 57554 57922 57622 57978
rect 57678 57922 57774 57978
rect 57154 40350 57774 57922
rect 57154 40294 57250 40350
rect 57306 40294 57374 40350
rect 57430 40294 57498 40350
rect 57554 40294 57622 40350
rect 57678 40294 57774 40350
rect 57154 40226 57774 40294
rect 57154 40170 57250 40226
rect 57306 40170 57374 40226
rect 57430 40170 57498 40226
rect 57554 40170 57622 40226
rect 57678 40170 57774 40226
rect 57154 40102 57774 40170
rect 57154 40046 57250 40102
rect 57306 40046 57374 40102
rect 57430 40046 57498 40102
rect 57554 40046 57622 40102
rect 57678 40046 57774 40102
rect 57154 39978 57774 40046
rect 57154 39922 57250 39978
rect 57306 39922 57374 39978
rect 57430 39922 57498 39978
rect 57554 39922 57622 39978
rect 57678 39922 57774 39978
rect 57154 22350 57774 39922
rect 57154 22294 57250 22350
rect 57306 22294 57374 22350
rect 57430 22294 57498 22350
rect 57554 22294 57622 22350
rect 57678 22294 57774 22350
rect 57154 22226 57774 22294
rect 57154 22170 57250 22226
rect 57306 22170 57374 22226
rect 57430 22170 57498 22226
rect 57554 22170 57622 22226
rect 57678 22170 57774 22226
rect 57154 22102 57774 22170
rect 57154 22046 57250 22102
rect 57306 22046 57374 22102
rect 57430 22046 57498 22102
rect 57554 22046 57622 22102
rect 57678 22046 57774 22102
rect 57154 21978 57774 22046
rect 57154 21922 57250 21978
rect 57306 21922 57374 21978
rect 57430 21922 57498 21978
rect 57554 21922 57622 21978
rect 57678 21922 57774 21978
rect 52108 16482 52164 16492
rect 48748 12786 48804 12796
rect 42874 10294 42970 10350
rect 43026 10294 43094 10350
rect 43150 10294 43218 10350
rect 43274 10294 43342 10350
rect 43398 10294 43494 10350
rect 42874 10226 43494 10294
rect 42874 10170 42970 10226
rect 43026 10170 43094 10226
rect 43150 10170 43218 10226
rect 43274 10170 43342 10226
rect 43398 10170 43494 10226
rect 42874 10102 43494 10170
rect 42874 10046 42970 10102
rect 43026 10046 43094 10102
rect 43150 10046 43218 10102
rect 43274 10046 43342 10102
rect 43398 10046 43494 10102
rect 42874 9978 43494 10046
rect 42874 9922 42970 9978
rect 43026 9922 43094 9978
rect 43150 9922 43218 9978
rect 43274 9922 43342 9978
rect 43398 9922 43494 9978
rect 42874 -1120 43494 9922
rect 42874 -1176 42970 -1120
rect 43026 -1176 43094 -1120
rect 43150 -1176 43218 -1120
rect 43274 -1176 43342 -1120
rect 43398 -1176 43494 -1120
rect 42874 -1244 43494 -1176
rect 42874 -1300 42970 -1244
rect 43026 -1300 43094 -1244
rect 43150 -1300 43218 -1244
rect 43274 -1300 43342 -1244
rect 43398 -1300 43494 -1244
rect 42874 -1368 43494 -1300
rect 42874 -1424 42970 -1368
rect 43026 -1424 43094 -1368
rect 43150 -1424 43218 -1368
rect 43274 -1424 43342 -1368
rect 43398 -1424 43494 -1368
rect 42874 -1492 43494 -1424
rect 42874 -1548 42970 -1492
rect 43026 -1548 43094 -1492
rect 43150 -1548 43218 -1492
rect 43274 -1548 43342 -1492
rect 43398 -1548 43494 -1492
rect 42874 -1644 43494 -1548
rect 57154 4350 57774 21922
rect 58828 68516 58884 68526
rect 58828 18452 58884 68460
rect 60732 68516 60788 68526
rect 60732 21140 60788 68460
rect 60732 21074 60788 21084
rect 60874 64350 61494 77594
rect 60874 64294 60970 64350
rect 61026 64294 61094 64350
rect 61150 64294 61218 64350
rect 61274 64294 61342 64350
rect 61398 64294 61494 64350
rect 60874 64226 61494 64294
rect 60874 64170 60970 64226
rect 61026 64170 61094 64226
rect 61150 64170 61218 64226
rect 61274 64170 61342 64226
rect 61398 64170 61494 64226
rect 60874 64102 61494 64170
rect 60874 64046 60970 64102
rect 61026 64046 61094 64102
rect 61150 64046 61218 64102
rect 61274 64046 61342 64102
rect 61398 64046 61494 64102
rect 60874 63978 61494 64046
rect 60874 63922 60970 63978
rect 61026 63922 61094 63978
rect 61150 63922 61218 63978
rect 61274 63922 61342 63978
rect 61398 63922 61494 63978
rect 60874 46350 61494 63922
rect 75154 76350 75774 77594
rect 75154 76294 75250 76350
rect 75306 76294 75374 76350
rect 75430 76294 75498 76350
rect 75554 76294 75622 76350
rect 75678 76294 75774 76350
rect 75154 76226 75774 76294
rect 75154 76170 75250 76226
rect 75306 76170 75374 76226
rect 75430 76170 75498 76226
rect 75554 76170 75622 76226
rect 75678 76170 75774 76226
rect 75154 76102 75774 76170
rect 75154 76046 75250 76102
rect 75306 76046 75374 76102
rect 75430 76046 75498 76102
rect 75554 76046 75622 76102
rect 75678 76046 75774 76102
rect 75154 75978 75774 76046
rect 75154 75922 75250 75978
rect 75306 75922 75374 75978
rect 75430 75922 75498 75978
rect 75554 75922 75622 75978
rect 75678 75922 75774 75978
rect 75154 58350 75774 75922
rect 75154 58294 75250 58350
rect 75306 58294 75374 58350
rect 75430 58294 75498 58350
rect 75554 58294 75622 58350
rect 75678 58294 75774 58350
rect 75154 58226 75774 58294
rect 75154 58170 75250 58226
rect 75306 58170 75374 58226
rect 75430 58170 75498 58226
rect 75554 58170 75622 58226
rect 75678 58170 75774 58226
rect 75154 58102 75774 58170
rect 75154 58046 75250 58102
rect 75306 58046 75374 58102
rect 75430 58046 75498 58102
rect 75554 58046 75622 58102
rect 75678 58046 75774 58102
rect 75154 57978 75774 58046
rect 75154 57922 75250 57978
rect 75306 57922 75374 57978
rect 75430 57922 75498 57978
rect 75554 57922 75622 57978
rect 75678 57922 75774 57978
rect 64540 53732 64596 53742
rect 60874 46294 60970 46350
rect 61026 46294 61094 46350
rect 61150 46294 61218 46350
rect 61274 46294 61342 46350
rect 61398 46294 61494 46350
rect 60874 46226 61494 46294
rect 60874 46170 60970 46226
rect 61026 46170 61094 46226
rect 61150 46170 61218 46226
rect 61274 46170 61342 46226
rect 61398 46170 61494 46226
rect 60874 46102 61494 46170
rect 60874 46046 60970 46102
rect 61026 46046 61094 46102
rect 61150 46046 61218 46102
rect 61274 46046 61342 46102
rect 61398 46046 61494 46102
rect 60874 45978 61494 46046
rect 60874 45922 60970 45978
rect 61026 45922 61094 45978
rect 61150 45922 61218 45978
rect 61274 45922 61342 45978
rect 61398 45922 61494 45978
rect 60874 28350 61494 45922
rect 64316 46452 64372 46462
rect 61964 35588 62020 35598
rect 60874 28294 60970 28350
rect 61026 28294 61094 28350
rect 61150 28294 61218 28350
rect 61274 28294 61342 28350
rect 61398 28294 61494 28350
rect 60874 28226 61494 28294
rect 60874 28170 60970 28226
rect 61026 28170 61094 28226
rect 61150 28170 61218 28226
rect 61274 28170 61342 28226
rect 61398 28170 61494 28226
rect 60874 28102 61494 28170
rect 60874 28046 60970 28102
rect 61026 28046 61094 28102
rect 61150 28046 61218 28102
rect 61274 28046 61342 28102
rect 61398 28046 61494 28102
rect 60874 27978 61494 28046
rect 60874 27922 60970 27978
rect 61026 27922 61094 27978
rect 61150 27922 61218 27978
rect 61274 27922 61342 27978
rect 61398 27922 61494 27978
rect 60620 20916 60676 20926
rect 60620 19684 60676 20860
rect 60620 19618 60676 19628
rect 58828 18386 58884 18396
rect 57154 4294 57250 4350
rect 57306 4294 57374 4350
rect 57430 4294 57498 4350
rect 57554 4294 57622 4350
rect 57678 4294 57774 4350
rect 57154 4226 57774 4294
rect 57154 4170 57250 4226
rect 57306 4170 57374 4226
rect 57430 4170 57498 4226
rect 57554 4170 57622 4226
rect 57678 4170 57774 4226
rect 57154 4102 57774 4170
rect 57154 4046 57250 4102
rect 57306 4046 57374 4102
rect 57430 4046 57498 4102
rect 57554 4046 57622 4102
rect 57678 4046 57774 4102
rect 57154 3978 57774 4046
rect 57154 3922 57250 3978
rect 57306 3922 57374 3978
rect 57430 3922 57498 3978
rect 57554 3922 57622 3978
rect 57678 3922 57774 3978
rect 57154 -160 57774 3922
rect 57154 -216 57250 -160
rect 57306 -216 57374 -160
rect 57430 -216 57498 -160
rect 57554 -216 57622 -160
rect 57678 -216 57774 -160
rect 57154 -284 57774 -216
rect 57154 -340 57250 -284
rect 57306 -340 57374 -284
rect 57430 -340 57498 -284
rect 57554 -340 57622 -284
rect 57678 -340 57774 -284
rect 57154 -408 57774 -340
rect 57154 -464 57250 -408
rect 57306 -464 57374 -408
rect 57430 -464 57498 -408
rect 57554 -464 57622 -408
rect 57678 -464 57774 -408
rect 57154 -532 57774 -464
rect 57154 -588 57250 -532
rect 57306 -588 57374 -532
rect 57430 -588 57498 -532
rect 57554 -588 57622 -532
rect 57678 -588 57774 -532
rect 57154 -1644 57774 -588
rect 60874 10350 61494 27922
rect 61740 34804 61796 34814
rect 61628 23940 61684 23950
rect 61628 21364 61684 23884
rect 61628 21298 61684 21308
rect 61628 20916 61684 20926
rect 61740 20916 61796 34748
rect 61964 27188 62020 35532
rect 64092 33348 64148 33358
rect 61964 27122 62020 27132
rect 63868 30436 63924 30446
rect 61684 20860 61796 20916
rect 61852 21700 61908 21710
rect 61628 20850 61684 20860
rect 61852 20244 61908 21644
rect 63868 21476 63924 30380
rect 63868 21410 63924 21420
rect 63980 27524 64036 27534
rect 61852 20178 61908 20188
rect 63980 19460 64036 27468
rect 63980 19394 64036 19404
rect 64092 18116 64148 33292
rect 64204 28980 64260 28990
rect 64204 19908 64260 28924
rect 64204 19842 64260 19852
rect 64316 18340 64372 46396
rect 64316 18274 64372 18284
rect 64092 18050 64148 18060
rect 64540 14756 64596 53676
rect 64540 14690 64596 14700
rect 75154 40350 75774 57922
rect 75154 40294 75250 40350
rect 75306 40294 75374 40350
rect 75430 40294 75498 40350
rect 75554 40294 75622 40350
rect 75678 40294 75774 40350
rect 75154 40226 75774 40294
rect 75154 40170 75250 40226
rect 75306 40170 75374 40226
rect 75430 40170 75498 40226
rect 75554 40170 75622 40226
rect 75678 40170 75774 40226
rect 75154 40102 75774 40170
rect 75154 40046 75250 40102
rect 75306 40046 75374 40102
rect 75430 40046 75498 40102
rect 75554 40046 75622 40102
rect 75678 40046 75774 40102
rect 75154 39978 75774 40046
rect 75154 39922 75250 39978
rect 75306 39922 75374 39978
rect 75430 39922 75498 39978
rect 75554 39922 75622 39978
rect 75678 39922 75774 39978
rect 75154 22350 75774 39922
rect 75154 22294 75250 22350
rect 75306 22294 75374 22350
rect 75430 22294 75498 22350
rect 75554 22294 75622 22350
rect 75678 22294 75774 22350
rect 75154 22226 75774 22294
rect 75154 22170 75250 22226
rect 75306 22170 75374 22226
rect 75430 22170 75498 22226
rect 75554 22170 75622 22226
rect 75678 22170 75774 22226
rect 75154 22102 75774 22170
rect 75154 22046 75250 22102
rect 75306 22046 75374 22102
rect 75430 22046 75498 22102
rect 75554 22046 75622 22102
rect 75678 22046 75774 22102
rect 75154 21978 75774 22046
rect 75154 21922 75250 21978
rect 75306 21922 75374 21978
rect 75430 21922 75498 21978
rect 75554 21922 75622 21978
rect 75678 21922 75774 21978
rect 60874 10294 60970 10350
rect 61026 10294 61094 10350
rect 61150 10294 61218 10350
rect 61274 10294 61342 10350
rect 61398 10294 61494 10350
rect 60874 10226 61494 10294
rect 60874 10170 60970 10226
rect 61026 10170 61094 10226
rect 61150 10170 61218 10226
rect 61274 10170 61342 10226
rect 61398 10170 61494 10226
rect 60874 10102 61494 10170
rect 60874 10046 60970 10102
rect 61026 10046 61094 10102
rect 61150 10046 61218 10102
rect 61274 10046 61342 10102
rect 61398 10046 61494 10102
rect 60874 9978 61494 10046
rect 60874 9922 60970 9978
rect 61026 9922 61094 9978
rect 61150 9922 61218 9978
rect 61274 9922 61342 9978
rect 61398 9922 61494 9978
rect 60874 -1120 61494 9922
rect 60874 -1176 60970 -1120
rect 61026 -1176 61094 -1120
rect 61150 -1176 61218 -1120
rect 61274 -1176 61342 -1120
rect 61398 -1176 61494 -1120
rect 60874 -1244 61494 -1176
rect 60874 -1300 60970 -1244
rect 61026 -1300 61094 -1244
rect 61150 -1300 61218 -1244
rect 61274 -1300 61342 -1244
rect 61398 -1300 61494 -1244
rect 60874 -1368 61494 -1300
rect 60874 -1424 60970 -1368
rect 61026 -1424 61094 -1368
rect 61150 -1424 61218 -1368
rect 61274 -1424 61342 -1368
rect 61398 -1424 61494 -1368
rect 60874 -1492 61494 -1424
rect 60874 -1548 60970 -1492
rect 61026 -1548 61094 -1492
rect 61150 -1548 61218 -1492
rect 61274 -1548 61342 -1492
rect 61398 -1548 61494 -1492
rect 60874 -1644 61494 -1548
rect 75154 4350 75774 21922
rect 75154 4294 75250 4350
rect 75306 4294 75374 4350
rect 75430 4294 75498 4350
rect 75554 4294 75622 4350
rect 75678 4294 75774 4350
rect 75154 4226 75774 4294
rect 75154 4170 75250 4226
rect 75306 4170 75374 4226
rect 75430 4170 75498 4226
rect 75554 4170 75622 4226
rect 75678 4170 75774 4226
rect 75154 4102 75774 4170
rect 75154 4046 75250 4102
rect 75306 4046 75374 4102
rect 75430 4046 75498 4102
rect 75554 4046 75622 4102
rect 75678 4046 75774 4102
rect 75154 3978 75774 4046
rect 75154 3922 75250 3978
rect 75306 3922 75374 3978
rect 75430 3922 75498 3978
rect 75554 3922 75622 3978
rect 75678 3922 75774 3978
rect 75154 -160 75774 3922
rect 75154 -216 75250 -160
rect 75306 -216 75374 -160
rect 75430 -216 75498 -160
rect 75554 -216 75622 -160
rect 75678 -216 75774 -160
rect 75154 -284 75774 -216
rect 75154 -340 75250 -284
rect 75306 -340 75374 -284
rect 75430 -340 75498 -284
rect 75554 -340 75622 -284
rect 75678 -340 75774 -284
rect 75154 -408 75774 -340
rect 75154 -464 75250 -408
rect 75306 -464 75374 -408
rect 75430 -464 75498 -408
rect 75554 -464 75622 -408
rect 75678 -464 75774 -408
rect 75154 -532 75774 -464
rect 75154 -588 75250 -532
rect 75306 -588 75374 -532
rect 75430 -588 75498 -532
rect 75554 -588 75622 -532
rect 75678 -588 75774 -532
rect 75154 -1644 75774 -588
rect 78874 64350 79494 77594
rect 78874 64294 78970 64350
rect 79026 64294 79094 64350
rect 79150 64294 79218 64350
rect 79274 64294 79342 64350
rect 79398 64294 79494 64350
rect 78874 64226 79494 64294
rect 78874 64170 78970 64226
rect 79026 64170 79094 64226
rect 79150 64170 79218 64226
rect 79274 64170 79342 64226
rect 79398 64170 79494 64226
rect 78874 64102 79494 64170
rect 78874 64046 78970 64102
rect 79026 64046 79094 64102
rect 79150 64046 79218 64102
rect 79274 64046 79342 64102
rect 79398 64046 79494 64102
rect 78874 63978 79494 64046
rect 78874 63922 78970 63978
rect 79026 63922 79094 63978
rect 79150 63922 79218 63978
rect 79274 63922 79342 63978
rect 79398 63922 79494 63978
rect 78874 46350 79494 63922
rect 78874 46294 78970 46350
rect 79026 46294 79094 46350
rect 79150 46294 79218 46350
rect 79274 46294 79342 46350
rect 79398 46294 79494 46350
rect 78874 46226 79494 46294
rect 78874 46170 78970 46226
rect 79026 46170 79094 46226
rect 79150 46170 79218 46226
rect 79274 46170 79342 46226
rect 79398 46170 79494 46226
rect 78874 46102 79494 46170
rect 78874 46046 78970 46102
rect 79026 46046 79094 46102
rect 79150 46046 79218 46102
rect 79274 46046 79342 46102
rect 79398 46046 79494 46102
rect 78874 45978 79494 46046
rect 78874 45922 78970 45978
rect 79026 45922 79094 45978
rect 79150 45922 79218 45978
rect 79274 45922 79342 45978
rect 79398 45922 79494 45978
rect 78874 28350 79494 45922
rect 78874 28294 78970 28350
rect 79026 28294 79094 28350
rect 79150 28294 79218 28350
rect 79274 28294 79342 28350
rect 79398 28294 79494 28350
rect 78874 28226 79494 28294
rect 78874 28170 78970 28226
rect 79026 28170 79094 28226
rect 79150 28170 79218 28226
rect 79274 28170 79342 28226
rect 79398 28170 79494 28226
rect 78874 28102 79494 28170
rect 78874 28046 78970 28102
rect 79026 28046 79094 28102
rect 79150 28046 79218 28102
rect 79274 28046 79342 28102
rect 79398 28046 79494 28102
rect 78874 27978 79494 28046
rect 78874 27922 78970 27978
rect 79026 27922 79094 27978
rect 79150 27922 79218 27978
rect 79274 27922 79342 27978
rect 79398 27922 79494 27978
rect 78874 10350 79494 27922
rect 78874 10294 78970 10350
rect 79026 10294 79094 10350
rect 79150 10294 79218 10350
rect 79274 10294 79342 10350
rect 79398 10294 79494 10350
rect 78874 10226 79494 10294
rect 78874 10170 78970 10226
rect 79026 10170 79094 10226
rect 79150 10170 79218 10226
rect 79274 10170 79342 10226
rect 79398 10170 79494 10226
rect 78874 10102 79494 10170
rect 78874 10046 78970 10102
rect 79026 10046 79094 10102
rect 79150 10046 79218 10102
rect 79274 10046 79342 10102
rect 79398 10046 79494 10102
rect 78874 9978 79494 10046
rect 78874 9922 78970 9978
rect 79026 9922 79094 9978
rect 79150 9922 79218 9978
rect 79274 9922 79342 9978
rect 79398 9922 79494 9978
rect 78874 -1120 79494 9922
rect 78874 -1176 78970 -1120
rect 79026 -1176 79094 -1120
rect 79150 -1176 79218 -1120
rect 79274 -1176 79342 -1120
rect 79398 -1176 79494 -1120
rect 78874 -1244 79494 -1176
rect 78874 -1300 78970 -1244
rect 79026 -1300 79094 -1244
rect 79150 -1300 79218 -1244
rect 79274 -1300 79342 -1244
rect 79398 -1300 79494 -1244
rect 78874 -1368 79494 -1300
rect 78874 -1424 78970 -1368
rect 79026 -1424 79094 -1368
rect 79150 -1424 79218 -1368
rect 79274 -1424 79342 -1368
rect 79398 -1424 79494 -1368
rect 78874 -1492 79494 -1424
rect 78874 -1548 78970 -1492
rect 79026 -1548 79094 -1492
rect 79150 -1548 79218 -1492
rect 79274 -1548 79342 -1492
rect 79398 -1548 79494 -1492
rect 78874 -1644 79494 -1548
rect 93154 76350 93774 77594
rect 93154 76294 93250 76350
rect 93306 76294 93374 76350
rect 93430 76294 93498 76350
rect 93554 76294 93622 76350
rect 93678 76294 93774 76350
rect 93154 76226 93774 76294
rect 93154 76170 93250 76226
rect 93306 76170 93374 76226
rect 93430 76170 93498 76226
rect 93554 76170 93622 76226
rect 93678 76170 93774 76226
rect 93154 76102 93774 76170
rect 93154 76046 93250 76102
rect 93306 76046 93374 76102
rect 93430 76046 93498 76102
rect 93554 76046 93622 76102
rect 93678 76046 93774 76102
rect 93154 75978 93774 76046
rect 93154 75922 93250 75978
rect 93306 75922 93374 75978
rect 93430 75922 93498 75978
rect 93554 75922 93622 75978
rect 93678 75922 93774 75978
rect 93154 58350 93774 75922
rect 93154 58294 93250 58350
rect 93306 58294 93374 58350
rect 93430 58294 93498 58350
rect 93554 58294 93622 58350
rect 93678 58294 93774 58350
rect 93154 58226 93774 58294
rect 93154 58170 93250 58226
rect 93306 58170 93374 58226
rect 93430 58170 93498 58226
rect 93554 58170 93622 58226
rect 93678 58170 93774 58226
rect 93154 58102 93774 58170
rect 93154 58046 93250 58102
rect 93306 58046 93374 58102
rect 93430 58046 93498 58102
rect 93554 58046 93622 58102
rect 93678 58046 93774 58102
rect 93154 57978 93774 58046
rect 93154 57922 93250 57978
rect 93306 57922 93374 57978
rect 93430 57922 93498 57978
rect 93554 57922 93622 57978
rect 93678 57922 93774 57978
rect 93154 40350 93774 57922
rect 93154 40294 93250 40350
rect 93306 40294 93374 40350
rect 93430 40294 93498 40350
rect 93554 40294 93622 40350
rect 93678 40294 93774 40350
rect 93154 40226 93774 40294
rect 93154 40170 93250 40226
rect 93306 40170 93374 40226
rect 93430 40170 93498 40226
rect 93554 40170 93622 40226
rect 93678 40170 93774 40226
rect 93154 40102 93774 40170
rect 93154 40046 93250 40102
rect 93306 40046 93374 40102
rect 93430 40046 93498 40102
rect 93554 40046 93622 40102
rect 93678 40046 93774 40102
rect 93154 39978 93774 40046
rect 93154 39922 93250 39978
rect 93306 39922 93374 39978
rect 93430 39922 93498 39978
rect 93554 39922 93622 39978
rect 93678 39922 93774 39978
rect 93154 22350 93774 39922
rect 93154 22294 93250 22350
rect 93306 22294 93374 22350
rect 93430 22294 93498 22350
rect 93554 22294 93622 22350
rect 93678 22294 93774 22350
rect 93154 22226 93774 22294
rect 93154 22170 93250 22226
rect 93306 22170 93374 22226
rect 93430 22170 93498 22226
rect 93554 22170 93622 22226
rect 93678 22170 93774 22226
rect 93154 22102 93774 22170
rect 93154 22046 93250 22102
rect 93306 22046 93374 22102
rect 93430 22046 93498 22102
rect 93554 22046 93622 22102
rect 93678 22046 93774 22102
rect 93154 21978 93774 22046
rect 93154 21922 93250 21978
rect 93306 21922 93374 21978
rect 93430 21922 93498 21978
rect 93554 21922 93622 21978
rect 93678 21922 93774 21978
rect 93154 4350 93774 21922
rect 93154 4294 93250 4350
rect 93306 4294 93374 4350
rect 93430 4294 93498 4350
rect 93554 4294 93622 4350
rect 93678 4294 93774 4350
rect 93154 4226 93774 4294
rect 93154 4170 93250 4226
rect 93306 4170 93374 4226
rect 93430 4170 93498 4226
rect 93554 4170 93622 4226
rect 93678 4170 93774 4226
rect 93154 4102 93774 4170
rect 93154 4046 93250 4102
rect 93306 4046 93374 4102
rect 93430 4046 93498 4102
rect 93554 4046 93622 4102
rect 93678 4046 93774 4102
rect 93154 3978 93774 4046
rect 93154 3922 93250 3978
rect 93306 3922 93374 3978
rect 93430 3922 93498 3978
rect 93554 3922 93622 3978
rect 93678 3922 93774 3978
rect 93154 -160 93774 3922
rect 93154 -216 93250 -160
rect 93306 -216 93374 -160
rect 93430 -216 93498 -160
rect 93554 -216 93622 -160
rect 93678 -216 93774 -160
rect 93154 -284 93774 -216
rect 93154 -340 93250 -284
rect 93306 -340 93374 -284
rect 93430 -340 93498 -284
rect 93554 -340 93622 -284
rect 93678 -340 93774 -284
rect 93154 -408 93774 -340
rect 93154 -464 93250 -408
rect 93306 -464 93374 -408
rect 93430 -464 93498 -408
rect 93554 -464 93622 -408
rect 93678 -464 93774 -408
rect 93154 -532 93774 -464
rect 93154 -588 93250 -532
rect 93306 -588 93374 -532
rect 93430 -588 93498 -532
rect 93554 -588 93622 -532
rect 93678 -588 93774 -532
rect 93154 -1644 93774 -588
rect 96874 64350 97494 77594
rect 96874 64294 96970 64350
rect 97026 64294 97094 64350
rect 97150 64294 97218 64350
rect 97274 64294 97342 64350
rect 97398 64294 97494 64350
rect 96874 64226 97494 64294
rect 96874 64170 96970 64226
rect 97026 64170 97094 64226
rect 97150 64170 97218 64226
rect 97274 64170 97342 64226
rect 97398 64170 97494 64226
rect 96874 64102 97494 64170
rect 96874 64046 96970 64102
rect 97026 64046 97094 64102
rect 97150 64046 97218 64102
rect 97274 64046 97342 64102
rect 97398 64046 97494 64102
rect 96874 63978 97494 64046
rect 96874 63922 96970 63978
rect 97026 63922 97094 63978
rect 97150 63922 97218 63978
rect 97274 63922 97342 63978
rect 97398 63922 97494 63978
rect 96874 46350 97494 63922
rect 96874 46294 96970 46350
rect 97026 46294 97094 46350
rect 97150 46294 97218 46350
rect 97274 46294 97342 46350
rect 97398 46294 97494 46350
rect 96874 46226 97494 46294
rect 96874 46170 96970 46226
rect 97026 46170 97094 46226
rect 97150 46170 97218 46226
rect 97274 46170 97342 46226
rect 97398 46170 97494 46226
rect 96874 46102 97494 46170
rect 96874 46046 96970 46102
rect 97026 46046 97094 46102
rect 97150 46046 97218 46102
rect 97274 46046 97342 46102
rect 97398 46046 97494 46102
rect 96874 45978 97494 46046
rect 96874 45922 96970 45978
rect 97026 45922 97094 45978
rect 97150 45922 97218 45978
rect 97274 45922 97342 45978
rect 97398 45922 97494 45978
rect 96874 28350 97494 45922
rect 96874 28294 96970 28350
rect 97026 28294 97094 28350
rect 97150 28294 97218 28350
rect 97274 28294 97342 28350
rect 97398 28294 97494 28350
rect 96874 28226 97494 28294
rect 96874 28170 96970 28226
rect 97026 28170 97094 28226
rect 97150 28170 97218 28226
rect 97274 28170 97342 28226
rect 97398 28170 97494 28226
rect 96874 28102 97494 28170
rect 96874 28046 96970 28102
rect 97026 28046 97094 28102
rect 97150 28046 97218 28102
rect 97274 28046 97342 28102
rect 97398 28046 97494 28102
rect 96874 27978 97494 28046
rect 96874 27922 96970 27978
rect 97026 27922 97094 27978
rect 97150 27922 97218 27978
rect 97274 27922 97342 27978
rect 97398 27922 97494 27978
rect 96874 10350 97494 27922
rect 96874 10294 96970 10350
rect 97026 10294 97094 10350
rect 97150 10294 97218 10350
rect 97274 10294 97342 10350
rect 97398 10294 97494 10350
rect 96874 10226 97494 10294
rect 96874 10170 96970 10226
rect 97026 10170 97094 10226
rect 97150 10170 97218 10226
rect 97274 10170 97342 10226
rect 97398 10170 97494 10226
rect 96874 10102 97494 10170
rect 96874 10046 96970 10102
rect 97026 10046 97094 10102
rect 97150 10046 97218 10102
rect 97274 10046 97342 10102
rect 97398 10046 97494 10102
rect 96874 9978 97494 10046
rect 96874 9922 96970 9978
rect 97026 9922 97094 9978
rect 97150 9922 97218 9978
rect 97274 9922 97342 9978
rect 97398 9922 97494 9978
rect 96874 -1120 97494 9922
rect 96874 -1176 96970 -1120
rect 97026 -1176 97094 -1120
rect 97150 -1176 97218 -1120
rect 97274 -1176 97342 -1120
rect 97398 -1176 97494 -1120
rect 96874 -1244 97494 -1176
rect 96874 -1300 96970 -1244
rect 97026 -1300 97094 -1244
rect 97150 -1300 97218 -1244
rect 97274 -1300 97342 -1244
rect 97398 -1300 97494 -1244
rect 96874 -1368 97494 -1300
rect 96874 -1424 96970 -1368
rect 97026 -1424 97094 -1368
rect 97150 -1424 97218 -1368
rect 97274 -1424 97342 -1368
rect 97398 -1424 97494 -1368
rect 96874 -1492 97494 -1424
rect 96874 -1548 96970 -1492
rect 97026 -1548 97094 -1492
rect 97150 -1548 97218 -1492
rect 97274 -1548 97342 -1492
rect 97398 -1548 97494 -1492
rect 96874 -1644 97494 -1548
rect 111154 76350 111774 77594
rect 111154 76294 111250 76350
rect 111306 76294 111374 76350
rect 111430 76294 111498 76350
rect 111554 76294 111622 76350
rect 111678 76294 111774 76350
rect 111154 76226 111774 76294
rect 111154 76170 111250 76226
rect 111306 76170 111374 76226
rect 111430 76170 111498 76226
rect 111554 76170 111622 76226
rect 111678 76170 111774 76226
rect 111154 76102 111774 76170
rect 111154 76046 111250 76102
rect 111306 76046 111374 76102
rect 111430 76046 111498 76102
rect 111554 76046 111622 76102
rect 111678 76046 111774 76102
rect 111154 75978 111774 76046
rect 111154 75922 111250 75978
rect 111306 75922 111374 75978
rect 111430 75922 111498 75978
rect 111554 75922 111622 75978
rect 111678 75922 111774 75978
rect 111154 58350 111774 75922
rect 111154 58294 111250 58350
rect 111306 58294 111374 58350
rect 111430 58294 111498 58350
rect 111554 58294 111622 58350
rect 111678 58294 111774 58350
rect 111154 58226 111774 58294
rect 111154 58170 111250 58226
rect 111306 58170 111374 58226
rect 111430 58170 111498 58226
rect 111554 58170 111622 58226
rect 111678 58170 111774 58226
rect 111154 58102 111774 58170
rect 111154 58046 111250 58102
rect 111306 58046 111374 58102
rect 111430 58046 111498 58102
rect 111554 58046 111622 58102
rect 111678 58046 111774 58102
rect 111154 57978 111774 58046
rect 111154 57922 111250 57978
rect 111306 57922 111374 57978
rect 111430 57922 111498 57978
rect 111554 57922 111622 57978
rect 111678 57922 111774 57978
rect 111154 40350 111774 57922
rect 111154 40294 111250 40350
rect 111306 40294 111374 40350
rect 111430 40294 111498 40350
rect 111554 40294 111622 40350
rect 111678 40294 111774 40350
rect 111154 40226 111774 40294
rect 111154 40170 111250 40226
rect 111306 40170 111374 40226
rect 111430 40170 111498 40226
rect 111554 40170 111622 40226
rect 111678 40170 111774 40226
rect 111154 40102 111774 40170
rect 111154 40046 111250 40102
rect 111306 40046 111374 40102
rect 111430 40046 111498 40102
rect 111554 40046 111622 40102
rect 111678 40046 111774 40102
rect 111154 39978 111774 40046
rect 111154 39922 111250 39978
rect 111306 39922 111374 39978
rect 111430 39922 111498 39978
rect 111554 39922 111622 39978
rect 111678 39922 111774 39978
rect 111154 22350 111774 39922
rect 111154 22294 111250 22350
rect 111306 22294 111374 22350
rect 111430 22294 111498 22350
rect 111554 22294 111622 22350
rect 111678 22294 111774 22350
rect 111154 22226 111774 22294
rect 111154 22170 111250 22226
rect 111306 22170 111374 22226
rect 111430 22170 111498 22226
rect 111554 22170 111622 22226
rect 111678 22170 111774 22226
rect 111154 22102 111774 22170
rect 111154 22046 111250 22102
rect 111306 22046 111374 22102
rect 111430 22046 111498 22102
rect 111554 22046 111622 22102
rect 111678 22046 111774 22102
rect 111154 21978 111774 22046
rect 111154 21922 111250 21978
rect 111306 21922 111374 21978
rect 111430 21922 111498 21978
rect 111554 21922 111622 21978
rect 111678 21922 111774 21978
rect 111154 4350 111774 21922
rect 111154 4294 111250 4350
rect 111306 4294 111374 4350
rect 111430 4294 111498 4350
rect 111554 4294 111622 4350
rect 111678 4294 111774 4350
rect 111154 4226 111774 4294
rect 111154 4170 111250 4226
rect 111306 4170 111374 4226
rect 111430 4170 111498 4226
rect 111554 4170 111622 4226
rect 111678 4170 111774 4226
rect 111154 4102 111774 4170
rect 111154 4046 111250 4102
rect 111306 4046 111374 4102
rect 111430 4046 111498 4102
rect 111554 4046 111622 4102
rect 111678 4046 111774 4102
rect 111154 3978 111774 4046
rect 111154 3922 111250 3978
rect 111306 3922 111374 3978
rect 111430 3922 111498 3978
rect 111554 3922 111622 3978
rect 111678 3922 111774 3978
rect 111154 -160 111774 3922
rect 111154 -216 111250 -160
rect 111306 -216 111374 -160
rect 111430 -216 111498 -160
rect 111554 -216 111622 -160
rect 111678 -216 111774 -160
rect 111154 -284 111774 -216
rect 111154 -340 111250 -284
rect 111306 -340 111374 -284
rect 111430 -340 111498 -284
rect 111554 -340 111622 -284
rect 111678 -340 111774 -284
rect 111154 -408 111774 -340
rect 111154 -464 111250 -408
rect 111306 -464 111374 -408
rect 111430 -464 111498 -408
rect 111554 -464 111622 -408
rect 111678 -464 111774 -408
rect 111154 -532 111774 -464
rect 111154 -588 111250 -532
rect 111306 -588 111374 -532
rect 111430 -588 111498 -532
rect 111554 -588 111622 -532
rect 111678 -588 111774 -532
rect 111154 -1644 111774 -588
rect 114874 64350 115494 77594
rect 114874 64294 114970 64350
rect 115026 64294 115094 64350
rect 115150 64294 115218 64350
rect 115274 64294 115342 64350
rect 115398 64294 115494 64350
rect 114874 64226 115494 64294
rect 114874 64170 114970 64226
rect 115026 64170 115094 64226
rect 115150 64170 115218 64226
rect 115274 64170 115342 64226
rect 115398 64170 115494 64226
rect 114874 64102 115494 64170
rect 114874 64046 114970 64102
rect 115026 64046 115094 64102
rect 115150 64046 115218 64102
rect 115274 64046 115342 64102
rect 115398 64046 115494 64102
rect 114874 63978 115494 64046
rect 114874 63922 114970 63978
rect 115026 63922 115094 63978
rect 115150 63922 115218 63978
rect 115274 63922 115342 63978
rect 115398 63922 115494 63978
rect 114874 46350 115494 63922
rect 114874 46294 114970 46350
rect 115026 46294 115094 46350
rect 115150 46294 115218 46350
rect 115274 46294 115342 46350
rect 115398 46294 115494 46350
rect 114874 46226 115494 46294
rect 114874 46170 114970 46226
rect 115026 46170 115094 46226
rect 115150 46170 115218 46226
rect 115274 46170 115342 46226
rect 115398 46170 115494 46226
rect 114874 46102 115494 46170
rect 114874 46046 114970 46102
rect 115026 46046 115094 46102
rect 115150 46046 115218 46102
rect 115274 46046 115342 46102
rect 115398 46046 115494 46102
rect 114874 45978 115494 46046
rect 114874 45922 114970 45978
rect 115026 45922 115094 45978
rect 115150 45922 115218 45978
rect 115274 45922 115342 45978
rect 115398 45922 115494 45978
rect 114874 28350 115494 45922
rect 114874 28294 114970 28350
rect 115026 28294 115094 28350
rect 115150 28294 115218 28350
rect 115274 28294 115342 28350
rect 115398 28294 115494 28350
rect 114874 28226 115494 28294
rect 114874 28170 114970 28226
rect 115026 28170 115094 28226
rect 115150 28170 115218 28226
rect 115274 28170 115342 28226
rect 115398 28170 115494 28226
rect 114874 28102 115494 28170
rect 114874 28046 114970 28102
rect 115026 28046 115094 28102
rect 115150 28046 115218 28102
rect 115274 28046 115342 28102
rect 115398 28046 115494 28102
rect 114874 27978 115494 28046
rect 114874 27922 114970 27978
rect 115026 27922 115094 27978
rect 115150 27922 115218 27978
rect 115274 27922 115342 27978
rect 115398 27922 115494 27978
rect 114874 10350 115494 27922
rect 114874 10294 114970 10350
rect 115026 10294 115094 10350
rect 115150 10294 115218 10350
rect 115274 10294 115342 10350
rect 115398 10294 115494 10350
rect 114874 10226 115494 10294
rect 114874 10170 114970 10226
rect 115026 10170 115094 10226
rect 115150 10170 115218 10226
rect 115274 10170 115342 10226
rect 115398 10170 115494 10226
rect 114874 10102 115494 10170
rect 114874 10046 114970 10102
rect 115026 10046 115094 10102
rect 115150 10046 115218 10102
rect 115274 10046 115342 10102
rect 115398 10046 115494 10102
rect 114874 9978 115494 10046
rect 114874 9922 114970 9978
rect 115026 9922 115094 9978
rect 115150 9922 115218 9978
rect 115274 9922 115342 9978
rect 115398 9922 115494 9978
rect 114874 -1120 115494 9922
rect 114874 -1176 114970 -1120
rect 115026 -1176 115094 -1120
rect 115150 -1176 115218 -1120
rect 115274 -1176 115342 -1120
rect 115398 -1176 115494 -1120
rect 114874 -1244 115494 -1176
rect 114874 -1300 114970 -1244
rect 115026 -1300 115094 -1244
rect 115150 -1300 115218 -1244
rect 115274 -1300 115342 -1244
rect 115398 -1300 115494 -1244
rect 114874 -1368 115494 -1300
rect 114874 -1424 114970 -1368
rect 115026 -1424 115094 -1368
rect 115150 -1424 115218 -1368
rect 115274 -1424 115342 -1368
rect 115398 -1424 115494 -1368
rect 114874 -1492 115494 -1424
rect 114874 -1548 114970 -1492
rect 115026 -1548 115094 -1492
rect 115150 -1548 115218 -1492
rect 115274 -1548 115342 -1492
rect 115398 -1548 115494 -1492
rect 114874 -1644 115494 -1548
rect 129154 76350 129774 77594
rect 129154 76294 129250 76350
rect 129306 76294 129374 76350
rect 129430 76294 129498 76350
rect 129554 76294 129622 76350
rect 129678 76294 129774 76350
rect 129154 76226 129774 76294
rect 129154 76170 129250 76226
rect 129306 76170 129374 76226
rect 129430 76170 129498 76226
rect 129554 76170 129622 76226
rect 129678 76170 129774 76226
rect 129154 76102 129774 76170
rect 129154 76046 129250 76102
rect 129306 76046 129374 76102
rect 129430 76046 129498 76102
rect 129554 76046 129622 76102
rect 129678 76046 129774 76102
rect 129154 75978 129774 76046
rect 129154 75922 129250 75978
rect 129306 75922 129374 75978
rect 129430 75922 129498 75978
rect 129554 75922 129622 75978
rect 129678 75922 129774 75978
rect 129154 58350 129774 75922
rect 129154 58294 129250 58350
rect 129306 58294 129374 58350
rect 129430 58294 129498 58350
rect 129554 58294 129622 58350
rect 129678 58294 129774 58350
rect 129154 58226 129774 58294
rect 129154 58170 129250 58226
rect 129306 58170 129374 58226
rect 129430 58170 129498 58226
rect 129554 58170 129622 58226
rect 129678 58170 129774 58226
rect 129154 58102 129774 58170
rect 129154 58046 129250 58102
rect 129306 58046 129374 58102
rect 129430 58046 129498 58102
rect 129554 58046 129622 58102
rect 129678 58046 129774 58102
rect 129154 57978 129774 58046
rect 129154 57922 129250 57978
rect 129306 57922 129374 57978
rect 129430 57922 129498 57978
rect 129554 57922 129622 57978
rect 129678 57922 129774 57978
rect 129154 40350 129774 57922
rect 129154 40294 129250 40350
rect 129306 40294 129374 40350
rect 129430 40294 129498 40350
rect 129554 40294 129622 40350
rect 129678 40294 129774 40350
rect 129154 40226 129774 40294
rect 129154 40170 129250 40226
rect 129306 40170 129374 40226
rect 129430 40170 129498 40226
rect 129554 40170 129622 40226
rect 129678 40170 129774 40226
rect 129154 40102 129774 40170
rect 129154 40046 129250 40102
rect 129306 40046 129374 40102
rect 129430 40046 129498 40102
rect 129554 40046 129622 40102
rect 129678 40046 129774 40102
rect 129154 39978 129774 40046
rect 129154 39922 129250 39978
rect 129306 39922 129374 39978
rect 129430 39922 129498 39978
rect 129554 39922 129622 39978
rect 129678 39922 129774 39978
rect 129154 22350 129774 39922
rect 129154 22294 129250 22350
rect 129306 22294 129374 22350
rect 129430 22294 129498 22350
rect 129554 22294 129622 22350
rect 129678 22294 129774 22350
rect 129154 22226 129774 22294
rect 129154 22170 129250 22226
rect 129306 22170 129374 22226
rect 129430 22170 129498 22226
rect 129554 22170 129622 22226
rect 129678 22170 129774 22226
rect 129154 22102 129774 22170
rect 129154 22046 129250 22102
rect 129306 22046 129374 22102
rect 129430 22046 129498 22102
rect 129554 22046 129622 22102
rect 129678 22046 129774 22102
rect 129154 21978 129774 22046
rect 129154 21922 129250 21978
rect 129306 21922 129374 21978
rect 129430 21922 129498 21978
rect 129554 21922 129622 21978
rect 129678 21922 129774 21978
rect 129154 4350 129774 21922
rect 129154 4294 129250 4350
rect 129306 4294 129374 4350
rect 129430 4294 129498 4350
rect 129554 4294 129622 4350
rect 129678 4294 129774 4350
rect 129154 4226 129774 4294
rect 129154 4170 129250 4226
rect 129306 4170 129374 4226
rect 129430 4170 129498 4226
rect 129554 4170 129622 4226
rect 129678 4170 129774 4226
rect 129154 4102 129774 4170
rect 129154 4046 129250 4102
rect 129306 4046 129374 4102
rect 129430 4046 129498 4102
rect 129554 4046 129622 4102
rect 129678 4046 129774 4102
rect 129154 3978 129774 4046
rect 129154 3922 129250 3978
rect 129306 3922 129374 3978
rect 129430 3922 129498 3978
rect 129554 3922 129622 3978
rect 129678 3922 129774 3978
rect 129154 -160 129774 3922
rect 129154 -216 129250 -160
rect 129306 -216 129374 -160
rect 129430 -216 129498 -160
rect 129554 -216 129622 -160
rect 129678 -216 129774 -160
rect 129154 -284 129774 -216
rect 129154 -340 129250 -284
rect 129306 -340 129374 -284
rect 129430 -340 129498 -284
rect 129554 -340 129622 -284
rect 129678 -340 129774 -284
rect 129154 -408 129774 -340
rect 129154 -464 129250 -408
rect 129306 -464 129374 -408
rect 129430 -464 129498 -408
rect 129554 -464 129622 -408
rect 129678 -464 129774 -408
rect 129154 -532 129774 -464
rect 129154 -588 129250 -532
rect 129306 -588 129374 -532
rect 129430 -588 129498 -532
rect 129554 -588 129622 -532
rect 129678 -588 129774 -532
rect 129154 -1644 129774 -588
rect 132874 64350 133494 77594
rect 132874 64294 132970 64350
rect 133026 64294 133094 64350
rect 133150 64294 133218 64350
rect 133274 64294 133342 64350
rect 133398 64294 133494 64350
rect 132874 64226 133494 64294
rect 132874 64170 132970 64226
rect 133026 64170 133094 64226
rect 133150 64170 133218 64226
rect 133274 64170 133342 64226
rect 133398 64170 133494 64226
rect 132874 64102 133494 64170
rect 132874 64046 132970 64102
rect 133026 64046 133094 64102
rect 133150 64046 133218 64102
rect 133274 64046 133342 64102
rect 133398 64046 133494 64102
rect 132874 63978 133494 64046
rect 132874 63922 132970 63978
rect 133026 63922 133094 63978
rect 133150 63922 133218 63978
rect 133274 63922 133342 63978
rect 133398 63922 133494 63978
rect 132874 46350 133494 63922
rect 132874 46294 132970 46350
rect 133026 46294 133094 46350
rect 133150 46294 133218 46350
rect 133274 46294 133342 46350
rect 133398 46294 133494 46350
rect 132874 46226 133494 46294
rect 132874 46170 132970 46226
rect 133026 46170 133094 46226
rect 133150 46170 133218 46226
rect 133274 46170 133342 46226
rect 133398 46170 133494 46226
rect 132874 46102 133494 46170
rect 132874 46046 132970 46102
rect 133026 46046 133094 46102
rect 133150 46046 133218 46102
rect 133274 46046 133342 46102
rect 133398 46046 133494 46102
rect 132874 45978 133494 46046
rect 132874 45922 132970 45978
rect 133026 45922 133094 45978
rect 133150 45922 133218 45978
rect 133274 45922 133342 45978
rect 133398 45922 133494 45978
rect 132874 28350 133494 45922
rect 132874 28294 132970 28350
rect 133026 28294 133094 28350
rect 133150 28294 133218 28350
rect 133274 28294 133342 28350
rect 133398 28294 133494 28350
rect 132874 28226 133494 28294
rect 132874 28170 132970 28226
rect 133026 28170 133094 28226
rect 133150 28170 133218 28226
rect 133274 28170 133342 28226
rect 133398 28170 133494 28226
rect 132874 28102 133494 28170
rect 132874 28046 132970 28102
rect 133026 28046 133094 28102
rect 133150 28046 133218 28102
rect 133274 28046 133342 28102
rect 133398 28046 133494 28102
rect 132874 27978 133494 28046
rect 132874 27922 132970 27978
rect 133026 27922 133094 27978
rect 133150 27922 133218 27978
rect 133274 27922 133342 27978
rect 133398 27922 133494 27978
rect 132874 10350 133494 27922
rect 132874 10294 132970 10350
rect 133026 10294 133094 10350
rect 133150 10294 133218 10350
rect 133274 10294 133342 10350
rect 133398 10294 133494 10350
rect 132874 10226 133494 10294
rect 132874 10170 132970 10226
rect 133026 10170 133094 10226
rect 133150 10170 133218 10226
rect 133274 10170 133342 10226
rect 133398 10170 133494 10226
rect 132874 10102 133494 10170
rect 132874 10046 132970 10102
rect 133026 10046 133094 10102
rect 133150 10046 133218 10102
rect 133274 10046 133342 10102
rect 133398 10046 133494 10102
rect 132874 9978 133494 10046
rect 132874 9922 132970 9978
rect 133026 9922 133094 9978
rect 133150 9922 133218 9978
rect 133274 9922 133342 9978
rect 133398 9922 133494 9978
rect 132874 -1120 133494 9922
rect 132874 -1176 132970 -1120
rect 133026 -1176 133094 -1120
rect 133150 -1176 133218 -1120
rect 133274 -1176 133342 -1120
rect 133398 -1176 133494 -1120
rect 132874 -1244 133494 -1176
rect 132874 -1300 132970 -1244
rect 133026 -1300 133094 -1244
rect 133150 -1300 133218 -1244
rect 133274 -1300 133342 -1244
rect 133398 -1300 133494 -1244
rect 132874 -1368 133494 -1300
rect 132874 -1424 132970 -1368
rect 133026 -1424 133094 -1368
rect 133150 -1424 133218 -1368
rect 133274 -1424 133342 -1368
rect 133398 -1424 133494 -1368
rect 132874 -1492 133494 -1424
rect 132874 -1548 132970 -1492
rect 133026 -1548 133094 -1492
rect 133150 -1548 133218 -1492
rect 133274 -1548 133342 -1492
rect 133398 -1548 133494 -1492
rect 132874 -1644 133494 -1548
rect 147154 76350 147774 77594
rect 147154 76294 147250 76350
rect 147306 76294 147374 76350
rect 147430 76294 147498 76350
rect 147554 76294 147622 76350
rect 147678 76294 147774 76350
rect 147154 76226 147774 76294
rect 147154 76170 147250 76226
rect 147306 76170 147374 76226
rect 147430 76170 147498 76226
rect 147554 76170 147622 76226
rect 147678 76170 147774 76226
rect 147154 76102 147774 76170
rect 147154 76046 147250 76102
rect 147306 76046 147374 76102
rect 147430 76046 147498 76102
rect 147554 76046 147622 76102
rect 147678 76046 147774 76102
rect 147154 75978 147774 76046
rect 147154 75922 147250 75978
rect 147306 75922 147374 75978
rect 147430 75922 147498 75978
rect 147554 75922 147622 75978
rect 147678 75922 147774 75978
rect 147154 58350 147774 75922
rect 147154 58294 147250 58350
rect 147306 58294 147374 58350
rect 147430 58294 147498 58350
rect 147554 58294 147622 58350
rect 147678 58294 147774 58350
rect 147154 58226 147774 58294
rect 147154 58170 147250 58226
rect 147306 58170 147374 58226
rect 147430 58170 147498 58226
rect 147554 58170 147622 58226
rect 147678 58170 147774 58226
rect 147154 58102 147774 58170
rect 147154 58046 147250 58102
rect 147306 58046 147374 58102
rect 147430 58046 147498 58102
rect 147554 58046 147622 58102
rect 147678 58046 147774 58102
rect 147154 57978 147774 58046
rect 147154 57922 147250 57978
rect 147306 57922 147374 57978
rect 147430 57922 147498 57978
rect 147554 57922 147622 57978
rect 147678 57922 147774 57978
rect 147154 40350 147774 57922
rect 147154 40294 147250 40350
rect 147306 40294 147374 40350
rect 147430 40294 147498 40350
rect 147554 40294 147622 40350
rect 147678 40294 147774 40350
rect 147154 40226 147774 40294
rect 147154 40170 147250 40226
rect 147306 40170 147374 40226
rect 147430 40170 147498 40226
rect 147554 40170 147622 40226
rect 147678 40170 147774 40226
rect 147154 40102 147774 40170
rect 147154 40046 147250 40102
rect 147306 40046 147374 40102
rect 147430 40046 147498 40102
rect 147554 40046 147622 40102
rect 147678 40046 147774 40102
rect 147154 39978 147774 40046
rect 147154 39922 147250 39978
rect 147306 39922 147374 39978
rect 147430 39922 147498 39978
rect 147554 39922 147622 39978
rect 147678 39922 147774 39978
rect 147154 22350 147774 39922
rect 147154 22294 147250 22350
rect 147306 22294 147374 22350
rect 147430 22294 147498 22350
rect 147554 22294 147622 22350
rect 147678 22294 147774 22350
rect 147154 22226 147774 22294
rect 147154 22170 147250 22226
rect 147306 22170 147374 22226
rect 147430 22170 147498 22226
rect 147554 22170 147622 22226
rect 147678 22170 147774 22226
rect 147154 22102 147774 22170
rect 147154 22046 147250 22102
rect 147306 22046 147374 22102
rect 147430 22046 147498 22102
rect 147554 22046 147622 22102
rect 147678 22046 147774 22102
rect 147154 21978 147774 22046
rect 147154 21922 147250 21978
rect 147306 21922 147374 21978
rect 147430 21922 147498 21978
rect 147554 21922 147622 21978
rect 147678 21922 147774 21978
rect 147154 4350 147774 21922
rect 147154 4294 147250 4350
rect 147306 4294 147374 4350
rect 147430 4294 147498 4350
rect 147554 4294 147622 4350
rect 147678 4294 147774 4350
rect 147154 4226 147774 4294
rect 147154 4170 147250 4226
rect 147306 4170 147374 4226
rect 147430 4170 147498 4226
rect 147554 4170 147622 4226
rect 147678 4170 147774 4226
rect 147154 4102 147774 4170
rect 147154 4046 147250 4102
rect 147306 4046 147374 4102
rect 147430 4046 147498 4102
rect 147554 4046 147622 4102
rect 147678 4046 147774 4102
rect 147154 3978 147774 4046
rect 147154 3922 147250 3978
rect 147306 3922 147374 3978
rect 147430 3922 147498 3978
rect 147554 3922 147622 3978
rect 147678 3922 147774 3978
rect 147154 -160 147774 3922
rect 147154 -216 147250 -160
rect 147306 -216 147374 -160
rect 147430 -216 147498 -160
rect 147554 -216 147622 -160
rect 147678 -216 147774 -160
rect 147154 -284 147774 -216
rect 147154 -340 147250 -284
rect 147306 -340 147374 -284
rect 147430 -340 147498 -284
rect 147554 -340 147622 -284
rect 147678 -340 147774 -284
rect 147154 -408 147774 -340
rect 147154 -464 147250 -408
rect 147306 -464 147374 -408
rect 147430 -464 147498 -408
rect 147554 -464 147622 -408
rect 147678 -464 147774 -408
rect 147154 -532 147774 -464
rect 147154 -588 147250 -532
rect 147306 -588 147374 -532
rect 147430 -588 147498 -532
rect 147554 -588 147622 -532
rect 147678 -588 147774 -532
rect 147154 -1644 147774 -588
rect 150874 64350 151494 77594
rect 150874 64294 150970 64350
rect 151026 64294 151094 64350
rect 151150 64294 151218 64350
rect 151274 64294 151342 64350
rect 151398 64294 151494 64350
rect 150874 64226 151494 64294
rect 150874 64170 150970 64226
rect 151026 64170 151094 64226
rect 151150 64170 151218 64226
rect 151274 64170 151342 64226
rect 151398 64170 151494 64226
rect 150874 64102 151494 64170
rect 150874 64046 150970 64102
rect 151026 64046 151094 64102
rect 151150 64046 151218 64102
rect 151274 64046 151342 64102
rect 151398 64046 151494 64102
rect 150874 63978 151494 64046
rect 150874 63922 150970 63978
rect 151026 63922 151094 63978
rect 151150 63922 151218 63978
rect 151274 63922 151342 63978
rect 151398 63922 151494 63978
rect 150874 46350 151494 63922
rect 150874 46294 150970 46350
rect 151026 46294 151094 46350
rect 151150 46294 151218 46350
rect 151274 46294 151342 46350
rect 151398 46294 151494 46350
rect 150874 46226 151494 46294
rect 150874 46170 150970 46226
rect 151026 46170 151094 46226
rect 151150 46170 151218 46226
rect 151274 46170 151342 46226
rect 151398 46170 151494 46226
rect 150874 46102 151494 46170
rect 150874 46046 150970 46102
rect 151026 46046 151094 46102
rect 151150 46046 151218 46102
rect 151274 46046 151342 46102
rect 151398 46046 151494 46102
rect 150874 45978 151494 46046
rect 150874 45922 150970 45978
rect 151026 45922 151094 45978
rect 151150 45922 151218 45978
rect 151274 45922 151342 45978
rect 151398 45922 151494 45978
rect 150874 28350 151494 45922
rect 150874 28294 150970 28350
rect 151026 28294 151094 28350
rect 151150 28294 151218 28350
rect 151274 28294 151342 28350
rect 151398 28294 151494 28350
rect 150874 28226 151494 28294
rect 150874 28170 150970 28226
rect 151026 28170 151094 28226
rect 151150 28170 151218 28226
rect 151274 28170 151342 28226
rect 151398 28170 151494 28226
rect 150874 28102 151494 28170
rect 150874 28046 150970 28102
rect 151026 28046 151094 28102
rect 151150 28046 151218 28102
rect 151274 28046 151342 28102
rect 151398 28046 151494 28102
rect 150874 27978 151494 28046
rect 150874 27922 150970 27978
rect 151026 27922 151094 27978
rect 151150 27922 151218 27978
rect 151274 27922 151342 27978
rect 151398 27922 151494 27978
rect 150874 10350 151494 27922
rect 150874 10294 150970 10350
rect 151026 10294 151094 10350
rect 151150 10294 151218 10350
rect 151274 10294 151342 10350
rect 151398 10294 151494 10350
rect 150874 10226 151494 10294
rect 150874 10170 150970 10226
rect 151026 10170 151094 10226
rect 151150 10170 151218 10226
rect 151274 10170 151342 10226
rect 151398 10170 151494 10226
rect 150874 10102 151494 10170
rect 150874 10046 150970 10102
rect 151026 10046 151094 10102
rect 151150 10046 151218 10102
rect 151274 10046 151342 10102
rect 151398 10046 151494 10102
rect 150874 9978 151494 10046
rect 150874 9922 150970 9978
rect 151026 9922 151094 9978
rect 151150 9922 151218 9978
rect 151274 9922 151342 9978
rect 151398 9922 151494 9978
rect 150874 -1120 151494 9922
rect 150874 -1176 150970 -1120
rect 151026 -1176 151094 -1120
rect 151150 -1176 151218 -1120
rect 151274 -1176 151342 -1120
rect 151398 -1176 151494 -1120
rect 150874 -1244 151494 -1176
rect 150874 -1300 150970 -1244
rect 151026 -1300 151094 -1244
rect 151150 -1300 151218 -1244
rect 151274 -1300 151342 -1244
rect 151398 -1300 151494 -1244
rect 150874 -1368 151494 -1300
rect 150874 -1424 150970 -1368
rect 151026 -1424 151094 -1368
rect 151150 -1424 151218 -1368
rect 151274 -1424 151342 -1368
rect 151398 -1424 151494 -1368
rect 150874 -1492 151494 -1424
rect 150874 -1548 150970 -1492
rect 151026 -1548 151094 -1492
rect 151150 -1548 151218 -1492
rect 151274 -1548 151342 -1492
rect 151398 -1548 151494 -1492
rect 150874 -1644 151494 -1548
rect 165154 76350 165774 77594
rect 165154 76294 165250 76350
rect 165306 76294 165374 76350
rect 165430 76294 165498 76350
rect 165554 76294 165622 76350
rect 165678 76294 165774 76350
rect 165154 76226 165774 76294
rect 165154 76170 165250 76226
rect 165306 76170 165374 76226
rect 165430 76170 165498 76226
rect 165554 76170 165622 76226
rect 165678 76170 165774 76226
rect 165154 76102 165774 76170
rect 165154 76046 165250 76102
rect 165306 76046 165374 76102
rect 165430 76046 165498 76102
rect 165554 76046 165622 76102
rect 165678 76046 165774 76102
rect 165154 75978 165774 76046
rect 165154 75922 165250 75978
rect 165306 75922 165374 75978
rect 165430 75922 165498 75978
rect 165554 75922 165622 75978
rect 165678 75922 165774 75978
rect 165154 58350 165774 75922
rect 165154 58294 165250 58350
rect 165306 58294 165374 58350
rect 165430 58294 165498 58350
rect 165554 58294 165622 58350
rect 165678 58294 165774 58350
rect 165154 58226 165774 58294
rect 165154 58170 165250 58226
rect 165306 58170 165374 58226
rect 165430 58170 165498 58226
rect 165554 58170 165622 58226
rect 165678 58170 165774 58226
rect 165154 58102 165774 58170
rect 165154 58046 165250 58102
rect 165306 58046 165374 58102
rect 165430 58046 165498 58102
rect 165554 58046 165622 58102
rect 165678 58046 165774 58102
rect 165154 57978 165774 58046
rect 165154 57922 165250 57978
rect 165306 57922 165374 57978
rect 165430 57922 165498 57978
rect 165554 57922 165622 57978
rect 165678 57922 165774 57978
rect 165154 40350 165774 57922
rect 165154 40294 165250 40350
rect 165306 40294 165374 40350
rect 165430 40294 165498 40350
rect 165554 40294 165622 40350
rect 165678 40294 165774 40350
rect 165154 40226 165774 40294
rect 165154 40170 165250 40226
rect 165306 40170 165374 40226
rect 165430 40170 165498 40226
rect 165554 40170 165622 40226
rect 165678 40170 165774 40226
rect 165154 40102 165774 40170
rect 165154 40046 165250 40102
rect 165306 40046 165374 40102
rect 165430 40046 165498 40102
rect 165554 40046 165622 40102
rect 165678 40046 165774 40102
rect 165154 39978 165774 40046
rect 165154 39922 165250 39978
rect 165306 39922 165374 39978
rect 165430 39922 165498 39978
rect 165554 39922 165622 39978
rect 165678 39922 165774 39978
rect 165154 22350 165774 39922
rect 165154 22294 165250 22350
rect 165306 22294 165374 22350
rect 165430 22294 165498 22350
rect 165554 22294 165622 22350
rect 165678 22294 165774 22350
rect 165154 22226 165774 22294
rect 165154 22170 165250 22226
rect 165306 22170 165374 22226
rect 165430 22170 165498 22226
rect 165554 22170 165622 22226
rect 165678 22170 165774 22226
rect 165154 22102 165774 22170
rect 165154 22046 165250 22102
rect 165306 22046 165374 22102
rect 165430 22046 165498 22102
rect 165554 22046 165622 22102
rect 165678 22046 165774 22102
rect 165154 21978 165774 22046
rect 165154 21922 165250 21978
rect 165306 21922 165374 21978
rect 165430 21922 165498 21978
rect 165554 21922 165622 21978
rect 165678 21922 165774 21978
rect 165154 4350 165774 21922
rect 165154 4294 165250 4350
rect 165306 4294 165374 4350
rect 165430 4294 165498 4350
rect 165554 4294 165622 4350
rect 165678 4294 165774 4350
rect 165154 4226 165774 4294
rect 165154 4170 165250 4226
rect 165306 4170 165374 4226
rect 165430 4170 165498 4226
rect 165554 4170 165622 4226
rect 165678 4170 165774 4226
rect 165154 4102 165774 4170
rect 165154 4046 165250 4102
rect 165306 4046 165374 4102
rect 165430 4046 165498 4102
rect 165554 4046 165622 4102
rect 165678 4046 165774 4102
rect 165154 3978 165774 4046
rect 165154 3922 165250 3978
rect 165306 3922 165374 3978
rect 165430 3922 165498 3978
rect 165554 3922 165622 3978
rect 165678 3922 165774 3978
rect 165154 -160 165774 3922
rect 165154 -216 165250 -160
rect 165306 -216 165374 -160
rect 165430 -216 165498 -160
rect 165554 -216 165622 -160
rect 165678 -216 165774 -160
rect 165154 -284 165774 -216
rect 165154 -340 165250 -284
rect 165306 -340 165374 -284
rect 165430 -340 165498 -284
rect 165554 -340 165622 -284
rect 165678 -340 165774 -284
rect 165154 -408 165774 -340
rect 165154 -464 165250 -408
rect 165306 -464 165374 -408
rect 165430 -464 165498 -408
rect 165554 -464 165622 -408
rect 165678 -464 165774 -408
rect 165154 -532 165774 -464
rect 165154 -588 165250 -532
rect 165306 -588 165374 -532
rect 165430 -588 165498 -532
rect 165554 -588 165622 -532
rect 165678 -588 165774 -532
rect 165154 -1644 165774 -588
rect 168874 64350 169494 77594
rect 168874 64294 168970 64350
rect 169026 64294 169094 64350
rect 169150 64294 169218 64350
rect 169274 64294 169342 64350
rect 169398 64294 169494 64350
rect 168874 64226 169494 64294
rect 168874 64170 168970 64226
rect 169026 64170 169094 64226
rect 169150 64170 169218 64226
rect 169274 64170 169342 64226
rect 169398 64170 169494 64226
rect 168874 64102 169494 64170
rect 168874 64046 168970 64102
rect 169026 64046 169094 64102
rect 169150 64046 169218 64102
rect 169274 64046 169342 64102
rect 169398 64046 169494 64102
rect 168874 63978 169494 64046
rect 168874 63922 168970 63978
rect 169026 63922 169094 63978
rect 169150 63922 169218 63978
rect 169274 63922 169342 63978
rect 169398 63922 169494 63978
rect 168874 46350 169494 63922
rect 168874 46294 168970 46350
rect 169026 46294 169094 46350
rect 169150 46294 169218 46350
rect 169274 46294 169342 46350
rect 169398 46294 169494 46350
rect 168874 46226 169494 46294
rect 168874 46170 168970 46226
rect 169026 46170 169094 46226
rect 169150 46170 169218 46226
rect 169274 46170 169342 46226
rect 169398 46170 169494 46226
rect 168874 46102 169494 46170
rect 168874 46046 168970 46102
rect 169026 46046 169094 46102
rect 169150 46046 169218 46102
rect 169274 46046 169342 46102
rect 169398 46046 169494 46102
rect 168874 45978 169494 46046
rect 168874 45922 168970 45978
rect 169026 45922 169094 45978
rect 169150 45922 169218 45978
rect 169274 45922 169342 45978
rect 169398 45922 169494 45978
rect 168874 28350 169494 45922
rect 168874 28294 168970 28350
rect 169026 28294 169094 28350
rect 169150 28294 169218 28350
rect 169274 28294 169342 28350
rect 169398 28294 169494 28350
rect 168874 28226 169494 28294
rect 168874 28170 168970 28226
rect 169026 28170 169094 28226
rect 169150 28170 169218 28226
rect 169274 28170 169342 28226
rect 169398 28170 169494 28226
rect 168874 28102 169494 28170
rect 168874 28046 168970 28102
rect 169026 28046 169094 28102
rect 169150 28046 169218 28102
rect 169274 28046 169342 28102
rect 169398 28046 169494 28102
rect 168874 27978 169494 28046
rect 168874 27922 168970 27978
rect 169026 27922 169094 27978
rect 169150 27922 169218 27978
rect 169274 27922 169342 27978
rect 169398 27922 169494 27978
rect 168874 10350 169494 27922
rect 168874 10294 168970 10350
rect 169026 10294 169094 10350
rect 169150 10294 169218 10350
rect 169274 10294 169342 10350
rect 169398 10294 169494 10350
rect 168874 10226 169494 10294
rect 168874 10170 168970 10226
rect 169026 10170 169094 10226
rect 169150 10170 169218 10226
rect 169274 10170 169342 10226
rect 169398 10170 169494 10226
rect 168874 10102 169494 10170
rect 168874 10046 168970 10102
rect 169026 10046 169094 10102
rect 169150 10046 169218 10102
rect 169274 10046 169342 10102
rect 169398 10046 169494 10102
rect 168874 9978 169494 10046
rect 168874 9922 168970 9978
rect 169026 9922 169094 9978
rect 169150 9922 169218 9978
rect 169274 9922 169342 9978
rect 169398 9922 169494 9978
rect 168874 -1120 169494 9922
rect 168874 -1176 168970 -1120
rect 169026 -1176 169094 -1120
rect 169150 -1176 169218 -1120
rect 169274 -1176 169342 -1120
rect 169398 -1176 169494 -1120
rect 168874 -1244 169494 -1176
rect 168874 -1300 168970 -1244
rect 169026 -1300 169094 -1244
rect 169150 -1300 169218 -1244
rect 169274 -1300 169342 -1244
rect 169398 -1300 169494 -1244
rect 168874 -1368 169494 -1300
rect 168874 -1424 168970 -1368
rect 169026 -1424 169094 -1368
rect 169150 -1424 169218 -1368
rect 169274 -1424 169342 -1368
rect 169398 -1424 169494 -1368
rect 168874 -1492 169494 -1424
rect 168874 -1548 168970 -1492
rect 169026 -1548 169094 -1492
rect 169150 -1548 169218 -1492
rect 169274 -1548 169342 -1492
rect 169398 -1548 169494 -1492
rect 168874 -1644 169494 -1548
rect 183154 76350 183774 93922
rect 183154 76294 183250 76350
rect 183306 76294 183374 76350
rect 183430 76294 183498 76350
rect 183554 76294 183622 76350
rect 183678 76294 183774 76350
rect 183154 76226 183774 76294
rect 183154 76170 183250 76226
rect 183306 76170 183374 76226
rect 183430 76170 183498 76226
rect 183554 76170 183622 76226
rect 183678 76170 183774 76226
rect 183154 76102 183774 76170
rect 183154 76046 183250 76102
rect 183306 76046 183374 76102
rect 183430 76046 183498 76102
rect 183554 76046 183622 76102
rect 183678 76046 183774 76102
rect 183154 75978 183774 76046
rect 183154 75922 183250 75978
rect 183306 75922 183374 75978
rect 183430 75922 183498 75978
rect 183554 75922 183622 75978
rect 183678 75922 183774 75978
rect 183154 58350 183774 75922
rect 183154 58294 183250 58350
rect 183306 58294 183374 58350
rect 183430 58294 183498 58350
rect 183554 58294 183622 58350
rect 183678 58294 183774 58350
rect 183154 58226 183774 58294
rect 183154 58170 183250 58226
rect 183306 58170 183374 58226
rect 183430 58170 183498 58226
rect 183554 58170 183622 58226
rect 183678 58170 183774 58226
rect 183154 58102 183774 58170
rect 183154 58046 183250 58102
rect 183306 58046 183374 58102
rect 183430 58046 183498 58102
rect 183554 58046 183622 58102
rect 183678 58046 183774 58102
rect 183154 57978 183774 58046
rect 183154 57922 183250 57978
rect 183306 57922 183374 57978
rect 183430 57922 183498 57978
rect 183554 57922 183622 57978
rect 183678 57922 183774 57978
rect 183154 40350 183774 57922
rect 183154 40294 183250 40350
rect 183306 40294 183374 40350
rect 183430 40294 183498 40350
rect 183554 40294 183622 40350
rect 183678 40294 183774 40350
rect 183154 40226 183774 40294
rect 183154 40170 183250 40226
rect 183306 40170 183374 40226
rect 183430 40170 183498 40226
rect 183554 40170 183622 40226
rect 183678 40170 183774 40226
rect 183154 40102 183774 40170
rect 183154 40046 183250 40102
rect 183306 40046 183374 40102
rect 183430 40046 183498 40102
rect 183554 40046 183622 40102
rect 183678 40046 183774 40102
rect 183154 39978 183774 40046
rect 183154 39922 183250 39978
rect 183306 39922 183374 39978
rect 183430 39922 183498 39978
rect 183554 39922 183622 39978
rect 183678 39922 183774 39978
rect 183154 22350 183774 39922
rect 183154 22294 183250 22350
rect 183306 22294 183374 22350
rect 183430 22294 183498 22350
rect 183554 22294 183622 22350
rect 183678 22294 183774 22350
rect 183154 22226 183774 22294
rect 183154 22170 183250 22226
rect 183306 22170 183374 22226
rect 183430 22170 183498 22226
rect 183554 22170 183622 22226
rect 183678 22170 183774 22226
rect 183154 22102 183774 22170
rect 183154 22046 183250 22102
rect 183306 22046 183374 22102
rect 183430 22046 183498 22102
rect 183554 22046 183622 22102
rect 183678 22046 183774 22102
rect 183154 21978 183774 22046
rect 183154 21922 183250 21978
rect 183306 21922 183374 21978
rect 183430 21922 183498 21978
rect 183554 21922 183622 21978
rect 183678 21922 183774 21978
rect 183154 4350 183774 21922
rect 183154 4294 183250 4350
rect 183306 4294 183374 4350
rect 183430 4294 183498 4350
rect 183554 4294 183622 4350
rect 183678 4294 183774 4350
rect 183154 4226 183774 4294
rect 183154 4170 183250 4226
rect 183306 4170 183374 4226
rect 183430 4170 183498 4226
rect 183554 4170 183622 4226
rect 183678 4170 183774 4226
rect 183154 4102 183774 4170
rect 183154 4046 183250 4102
rect 183306 4046 183374 4102
rect 183430 4046 183498 4102
rect 183554 4046 183622 4102
rect 183678 4046 183774 4102
rect 183154 3978 183774 4046
rect 183154 3922 183250 3978
rect 183306 3922 183374 3978
rect 183430 3922 183498 3978
rect 183554 3922 183622 3978
rect 183678 3922 183774 3978
rect 183154 -160 183774 3922
rect 183154 -216 183250 -160
rect 183306 -216 183374 -160
rect 183430 -216 183498 -160
rect 183554 -216 183622 -160
rect 183678 -216 183774 -160
rect 183154 -284 183774 -216
rect 183154 -340 183250 -284
rect 183306 -340 183374 -284
rect 183430 -340 183498 -284
rect 183554 -340 183622 -284
rect 183678 -340 183774 -284
rect 183154 -408 183774 -340
rect 183154 -464 183250 -408
rect 183306 -464 183374 -408
rect 183430 -464 183498 -408
rect 183554 -464 183622 -408
rect 183678 -464 183774 -408
rect 183154 -532 183774 -464
rect 183154 -588 183250 -532
rect 183306 -588 183374 -532
rect 183430 -588 183498 -532
rect 183554 -588 183622 -532
rect 183678 -588 183774 -532
rect 183154 -1644 183774 -588
rect 186874 154350 187494 158858
rect 186874 154294 186970 154350
rect 187026 154294 187094 154350
rect 187150 154294 187218 154350
rect 187274 154294 187342 154350
rect 187398 154294 187494 154350
rect 186874 154226 187494 154294
rect 186874 154170 186970 154226
rect 187026 154170 187094 154226
rect 187150 154170 187218 154226
rect 187274 154170 187342 154226
rect 187398 154170 187494 154226
rect 186874 154102 187494 154170
rect 186874 154046 186970 154102
rect 187026 154046 187094 154102
rect 187150 154046 187218 154102
rect 187274 154046 187342 154102
rect 187398 154046 187494 154102
rect 186874 153978 187494 154046
rect 186874 153922 186970 153978
rect 187026 153922 187094 153978
rect 187150 153922 187218 153978
rect 187274 153922 187342 153978
rect 187398 153922 187494 153978
rect 186874 136350 187494 153922
rect 186874 136294 186970 136350
rect 187026 136294 187094 136350
rect 187150 136294 187218 136350
rect 187274 136294 187342 136350
rect 187398 136294 187494 136350
rect 186874 136226 187494 136294
rect 186874 136170 186970 136226
rect 187026 136170 187094 136226
rect 187150 136170 187218 136226
rect 187274 136170 187342 136226
rect 187398 136170 187494 136226
rect 186874 136102 187494 136170
rect 186874 136046 186970 136102
rect 187026 136046 187094 136102
rect 187150 136046 187218 136102
rect 187274 136046 187342 136102
rect 187398 136046 187494 136102
rect 186874 135978 187494 136046
rect 186874 135922 186970 135978
rect 187026 135922 187094 135978
rect 187150 135922 187218 135978
rect 187274 135922 187342 135978
rect 187398 135922 187494 135978
rect 186874 118350 187494 135922
rect 186874 118294 186970 118350
rect 187026 118294 187094 118350
rect 187150 118294 187218 118350
rect 187274 118294 187342 118350
rect 187398 118294 187494 118350
rect 186874 118226 187494 118294
rect 186874 118170 186970 118226
rect 187026 118170 187094 118226
rect 187150 118170 187218 118226
rect 187274 118170 187342 118226
rect 187398 118170 187494 118226
rect 186874 118102 187494 118170
rect 186874 118046 186970 118102
rect 187026 118046 187094 118102
rect 187150 118046 187218 118102
rect 187274 118046 187342 118102
rect 187398 118046 187494 118102
rect 186874 117978 187494 118046
rect 186874 117922 186970 117978
rect 187026 117922 187094 117978
rect 187150 117922 187218 117978
rect 187274 117922 187342 117978
rect 187398 117922 187494 117978
rect 186874 100350 187494 117922
rect 186874 100294 186970 100350
rect 187026 100294 187094 100350
rect 187150 100294 187218 100350
rect 187274 100294 187342 100350
rect 187398 100294 187494 100350
rect 186874 100226 187494 100294
rect 186874 100170 186970 100226
rect 187026 100170 187094 100226
rect 187150 100170 187218 100226
rect 187274 100170 187342 100226
rect 187398 100170 187494 100226
rect 186874 100102 187494 100170
rect 186874 100046 186970 100102
rect 187026 100046 187094 100102
rect 187150 100046 187218 100102
rect 187274 100046 187342 100102
rect 187398 100046 187494 100102
rect 186874 99978 187494 100046
rect 186874 99922 186970 99978
rect 187026 99922 187094 99978
rect 187150 99922 187218 99978
rect 187274 99922 187342 99978
rect 187398 99922 187494 99978
rect 186874 82350 187494 99922
rect 186874 82294 186970 82350
rect 187026 82294 187094 82350
rect 187150 82294 187218 82350
rect 187274 82294 187342 82350
rect 187398 82294 187494 82350
rect 186874 82226 187494 82294
rect 186874 82170 186970 82226
rect 187026 82170 187094 82226
rect 187150 82170 187218 82226
rect 187274 82170 187342 82226
rect 187398 82170 187494 82226
rect 186874 82102 187494 82170
rect 186874 82046 186970 82102
rect 187026 82046 187094 82102
rect 187150 82046 187218 82102
rect 187274 82046 187342 82102
rect 187398 82046 187494 82102
rect 186874 81978 187494 82046
rect 186874 81922 186970 81978
rect 187026 81922 187094 81978
rect 187150 81922 187218 81978
rect 187274 81922 187342 81978
rect 187398 81922 187494 81978
rect 186874 64350 187494 81922
rect 188972 66836 189028 306572
rect 189084 118580 189140 308252
rect 189196 140308 189252 316764
rect 189420 316708 189476 316718
rect 189420 305284 189476 316652
rect 189420 152628 189476 305228
rect 189420 149548 189476 152572
rect 189420 149492 189812 149548
rect 189196 140242 189252 140252
rect 189756 125972 189812 149492
rect 189756 124404 189812 125916
rect 189756 124338 189812 124348
rect 189084 118514 189140 118524
rect 190652 68964 190708 587468
rect 197372 587300 197428 587310
rect 194012 587188 194068 587198
rect 190876 539364 190932 539374
rect 190764 316708 190820 316718
rect 190764 145572 190820 316652
rect 190764 145506 190820 145516
rect 190876 69188 190932 539308
rect 190876 69122 190932 69132
rect 190652 68898 190708 68908
rect 188972 66770 189028 66780
rect 194012 65492 194068 587132
rect 195692 304948 195748 304958
rect 195692 118804 195748 304892
rect 197260 168084 197316 168094
rect 197260 155988 197316 168028
rect 197260 155922 197316 155932
rect 195804 155764 195860 155774
rect 195804 137060 195860 155708
rect 197036 153748 197092 153758
rect 196252 153412 196308 153422
rect 196252 138628 196308 153356
rect 196252 138562 196308 138572
rect 195804 136994 195860 137004
rect 197036 133588 197092 153692
rect 197036 133522 197092 133532
rect 195692 118738 195748 118748
rect 195916 116340 195972 116350
rect 194012 65426 194068 65436
rect 195692 116004 195748 116014
rect 186874 64294 186970 64350
rect 187026 64294 187094 64350
rect 187150 64294 187218 64350
rect 187274 64294 187342 64350
rect 187398 64294 187494 64350
rect 186874 64226 187494 64294
rect 186874 64170 186970 64226
rect 187026 64170 187094 64226
rect 187150 64170 187218 64226
rect 187274 64170 187342 64226
rect 187398 64170 187494 64226
rect 186874 64102 187494 64170
rect 186874 64046 186970 64102
rect 187026 64046 187094 64102
rect 187150 64046 187218 64102
rect 187274 64046 187342 64102
rect 187398 64046 187494 64102
rect 186874 63978 187494 64046
rect 186874 63922 186970 63978
rect 187026 63922 187094 63978
rect 187150 63922 187218 63978
rect 187274 63922 187342 63978
rect 187398 63922 187494 63978
rect 186874 46350 187494 63922
rect 186874 46294 186970 46350
rect 187026 46294 187094 46350
rect 187150 46294 187218 46350
rect 187274 46294 187342 46350
rect 187398 46294 187494 46350
rect 186874 46226 187494 46294
rect 186874 46170 186970 46226
rect 187026 46170 187094 46226
rect 187150 46170 187218 46226
rect 187274 46170 187342 46226
rect 187398 46170 187494 46226
rect 186874 46102 187494 46170
rect 186874 46046 186970 46102
rect 187026 46046 187094 46102
rect 187150 46046 187218 46102
rect 187274 46046 187342 46102
rect 187398 46046 187494 46102
rect 186874 45978 187494 46046
rect 186874 45922 186970 45978
rect 187026 45922 187094 45978
rect 187150 45922 187218 45978
rect 187274 45922 187342 45978
rect 187398 45922 187494 45978
rect 186874 28350 187494 45922
rect 186874 28294 186970 28350
rect 187026 28294 187094 28350
rect 187150 28294 187218 28350
rect 187274 28294 187342 28350
rect 187398 28294 187494 28350
rect 186874 28226 187494 28294
rect 186874 28170 186970 28226
rect 187026 28170 187094 28226
rect 187150 28170 187218 28226
rect 187274 28170 187342 28226
rect 187398 28170 187494 28226
rect 186874 28102 187494 28170
rect 186874 28046 186970 28102
rect 187026 28046 187094 28102
rect 187150 28046 187218 28102
rect 187274 28046 187342 28102
rect 187398 28046 187494 28102
rect 186874 27978 187494 28046
rect 186874 27922 186970 27978
rect 187026 27922 187094 27978
rect 187150 27922 187218 27978
rect 187274 27922 187342 27978
rect 187398 27922 187494 27978
rect 186874 10350 187494 27922
rect 186874 10294 186970 10350
rect 187026 10294 187094 10350
rect 187150 10294 187218 10350
rect 187274 10294 187342 10350
rect 187398 10294 187494 10350
rect 186874 10226 187494 10294
rect 186874 10170 186970 10226
rect 187026 10170 187094 10226
rect 187150 10170 187218 10226
rect 187274 10170 187342 10226
rect 187398 10170 187494 10226
rect 186874 10102 187494 10170
rect 186874 10046 186970 10102
rect 187026 10046 187094 10102
rect 187150 10046 187218 10102
rect 187274 10046 187342 10102
rect 187398 10046 187494 10102
rect 186874 9978 187494 10046
rect 186874 9922 186970 9978
rect 187026 9922 187094 9978
rect 187150 9922 187218 9978
rect 187274 9922 187342 9978
rect 187398 9922 187494 9978
rect 186874 -1120 187494 9922
rect 195692 6692 195748 115948
rect 195692 6626 195748 6636
rect 195916 4004 195972 116284
rect 196252 116116 196308 116126
rect 196252 10388 196308 116060
rect 197372 68852 197428 587244
rect 201154 580350 201774 596784
rect 201154 580294 201250 580350
rect 201306 580294 201374 580350
rect 201430 580294 201498 580350
rect 201554 580294 201622 580350
rect 201678 580294 201774 580350
rect 201154 580226 201774 580294
rect 201154 580170 201250 580226
rect 201306 580170 201374 580226
rect 201430 580170 201498 580226
rect 201554 580170 201622 580226
rect 201678 580170 201774 580226
rect 201154 580102 201774 580170
rect 201154 580046 201250 580102
rect 201306 580046 201374 580102
rect 201430 580046 201498 580102
rect 201554 580046 201622 580102
rect 201678 580046 201774 580102
rect 201154 579978 201774 580046
rect 201154 579922 201250 579978
rect 201306 579922 201374 579978
rect 201430 579922 201498 579978
rect 201554 579922 201622 579978
rect 201678 579922 201774 579978
rect 201154 562350 201774 579922
rect 201154 562294 201250 562350
rect 201306 562294 201374 562350
rect 201430 562294 201498 562350
rect 201554 562294 201622 562350
rect 201678 562294 201774 562350
rect 201154 562226 201774 562294
rect 201154 562170 201250 562226
rect 201306 562170 201374 562226
rect 201430 562170 201498 562226
rect 201554 562170 201622 562226
rect 201678 562170 201774 562226
rect 201154 562102 201774 562170
rect 201154 562046 201250 562102
rect 201306 562046 201374 562102
rect 201430 562046 201498 562102
rect 201554 562046 201622 562102
rect 201678 562046 201774 562102
rect 201154 561978 201774 562046
rect 201154 561922 201250 561978
rect 201306 561922 201374 561978
rect 201430 561922 201498 561978
rect 201554 561922 201622 561978
rect 201678 561922 201774 561978
rect 201154 544350 201774 561922
rect 201154 544294 201250 544350
rect 201306 544294 201374 544350
rect 201430 544294 201498 544350
rect 201554 544294 201622 544350
rect 201678 544294 201774 544350
rect 201154 544226 201774 544294
rect 201154 544170 201250 544226
rect 201306 544170 201374 544226
rect 201430 544170 201498 544226
rect 201554 544170 201622 544226
rect 201678 544170 201774 544226
rect 201154 544102 201774 544170
rect 201154 544046 201250 544102
rect 201306 544046 201374 544102
rect 201430 544046 201498 544102
rect 201554 544046 201622 544102
rect 201678 544046 201774 544102
rect 201154 543978 201774 544046
rect 201154 543922 201250 543978
rect 201306 543922 201374 543978
rect 201430 543922 201498 543978
rect 201554 543922 201622 543978
rect 201678 543922 201774 543978
rect 201154 526350 201774 543922
rect 201154 526294 201250 526350
rect 201306 526294 201374 526350
rect 201430 526294 201498 526350
rect 201554 526294 201622 526350
rect 201678 526294 201774 526350
rect 201154 526226 201774 526294
rect 201154 526170 201250 526226
rect 201306 526170 201374 526226
rect 201430 526170 201498 526226
rect 201554 526170 201622 526226
rect 201678 526170 201774 526226
rect 201154 526102 201774 526170
rect 201154 526046 201250 526102
rect 201306 526046 201374 526102
rect 201430 526046 201498 526102
rect 201554 526046 201622 526102
rect 201678 526046 201774 526102
rect 201154 525978 201774 526046
rect 201154 525922 201250 525978
rect 201306 525922 201374 525978
rect 201430 525922 201498 525978
rect 201554 525922 201622 525978
rect 201678 525922 201774 525978
rect 201154 508350 201774 525922
rect 201154 508294 201250 508350
rect 201306 508294 201374 508350
rect 201430 508294 201498 508350
rect 201554 508294 201622 508350
rect 201678 508294 201774 508350
rect 201154 508226 201774 508294
rect 201154 508170 201250 508226
rect 201306 508170 201374 508226
rect 201430 508170 201498 508226
rect 201554 508170 201622 508226
rect 201678 508170 201774 508226
rect 201154 508102 201774 508170
rect 201154 508046 201250 508102
rect 201306 508046 201374 508102
rect 201430 508046 201498 508102
rect 201554 508046 201622 508102
rect 201678 508046 201774 508102
rect 201154 507978 201774 508046
rect 201154 507922 201250 507978
rect 201306 507922 201374 507978
rect 201430 507922 201498 507978
rect 201554 507922 201622 507978
rect 201678 507922 201774 507978
rect 197596 494004 197652 494014
rect 197484 316932 197540 316942
rect 197484 142100 197540 316876
rect 197484 142034 197540 142044
rect 197372 68786 197428 68796
rect 197484 126084 197540 126094
rect 196252 10322 196308 10332
rect 197484 7364 197540 126028
rect 197596 68740 197652 493948
rect 201154 490350 201774 507922
rect 201154 490294 201250 490350
rect 201306 490294 201374 490350
rect 201430 490294 201498 490350
rect 201554 490294 201622 490350
rect 201678 490294 201774 490350
rect 201154 490226 201774 490294
rect 201154 490170 201250 490226
rect 201306 490170 201374 490226
rect 201430 490170 201498 490226
rect 201554 490170 201622 490226
rect 201678 490170 201774 490226
rect 201154 490102 201774 490170
rect 201154 490046 201250 490102
rect 201306 490046 201374 490102
rect 201430 490046 201498 490102
rect 201554 490046 201622 490102
rect 201678 490046 201774 490102
rect 201154 489978 201774 490046
rect 201154 489922 201250 489978
rect 201306 489922 201374 489978
rect 201430 489922 201498 489978
rect 201554 489922 201622 489978
rect 201678 489922 201774 489978
rect 201154 472350 201774 489922
rect 201154 472294 201250 472350
rect 201306 472294 201374 472350
rect 201430 472294 201498 472350
rect 201554 472294 201622 472350
rect 201678 472294 201774 472350
rect 201154 472226 201774 472294
rect 201154 472170 201250 472226
rect 201306 472170 201374 472226
rect 201430 472170 201498 472226
rect 201554 472170 201622 472226
rect 201678 472170 201774 472226
rect 201154 472102 201774 472170
rect 201154 472046 201250 472102
rect 201306 472046 201374 472102
rect 201430 472046 201498 472102
rect 201554 472046 201622 472102
rect 201678 472046 201774 472102
rect 201154 471978 201774 472046
rect 201154 471922 201250 471978
rect 201306 471922 201374 471978
rect 201430 471922 201498 471978
rect 201554 471922 201622 471978
rect 201678 471922 201774 471978
rect 201154 454350 201774 471922
rect 201154 454294 201250 454350
rect 201306 454294 201374 454350
rect 201430 454294 201498 454350
rect 201554 454294 201622 454350
rect 201678 454294 201774 454350
rect 201154 454226 201774 454294
rect 201154 454170 201250 454226
rect 201306 454170 201374 454226
rect 201430 454170 201498 454226
rect 201554 454170 201622 454226
rect 201678 454170 201774 454226
rect 201154 454102 201774 454170
rect 201154 454046 201250 454102
rect 201306 454046 201374 454102
rect 201430 454046 201498 454102
rect 201554 454046 201622 454102
rect 201678 454046 201774 454102
rect 201154 453978 201774 454046
rect 201154 453922 201250 453978
rect 201306 453922 201374 453978
rect 201430 453922 201498 453978
rect 201554 453922 201622 453978
rect 201678 453922 201774 453978
rect 201154 436350 201774 453922
rect 201154 436294 201250 436350
rect 201306 436294 201374 436350
rect 201430 436294 201498 436350
rect 201554 436294 201622 436350
rect 201678 436294 201774 436350
rect 201154 436226 201774 436294
rect 201154 436170 201250 436226
rect 201306 436170 201374 436226
rect 201430 436170 201498 436226
rect 201554 436170 201622 436226
rect 201678 436170 201774 436226
rect 201154 436102 201774 436170
rect 201154 436046 201250 436102
rect 201306 436046 201374 436102
rect 201430 436046 201498 436102
rect 201554 436046 201622 436102
rect 201678 436046 201774 436102
rect 201154 435978 201774 436046
rect 201154 435922 201250 435978
rect 201306 435922 201374 435978
rect 201430 435922 201498 435978
rect 201554 435922 201622 435978
rect 201678 435922 201774 435978
rect 201154 418350 201774 435922
rect 201154 418294 201250 418350
rect 201306 418294 201374 418350
rect 201430 418294 201498 418350
rect 201554 418294 201622 418350
rect 201678 418294 201774 418350
rect 201154 418226 201774 418294
rect 201154 418170 201250 418226
rect 201306 418170 201374 418226
rect 201430 418170 201498 418226
rect 201554 418170 201622 418226
rect 201678 418170 201774 418226
rect 201154 418102 201774 418170
rect 201154 418046 201250 418102
rect 201306 418046 201374 418102
rect 201430 418046 201498 418102
rect 201554 418046 201622 418102
rect 201678 418046 201774 418102
rect 201154 417978 201774 418046
rect 201154 417922 201250 417978
rect 201306 417922 201374 417978
rect 201430 417922 201498 417978
rect 201554 417922 201622 417978
rect 201678 417922 201774 417978
rect 201154 400350 201774 417922
rect 201154 400294 201250 400350
rect 201306 400294 201374 400350
rect 201430 400294 201498 400350
rect 201554 400294 201622 400350
rect 201678 400294 201774 400350
rect 201154 400226 201774 400294
rect 201154 400170 201250 400226
rect 201306 400170 201374 400226
rect 201430 400170 201498 400226
rect 201554 400170 201622 400226
rect 201678 400170 201774 400226
rect 201154 400102 201774 400170
rect 201154 400046 201250 400102
rect 201306 400046 201374 400102
rect 201430 400046 201498 400102
rect 201554 400046 201622 400102
rect 201678 400046 201774 400102
rect 201154 399978 201774 400046
rect 201154 399922 201250 399978
rect 201306 399922 201374 399978
rect 201430 399922 201498 399978
rect 201554 399922 201622 399978
rect 201678 399922 201774 399978
rect 201154 382350 201774 399922
rect 201154 382294 201250 382350
rect 201306 382294 201374 382350
rect 201430 382294 201498 382350
rect 201554 382294 201622 382350
rect 201678 382294 201774 382350
rect 201154 382226 201774 382294
rect 201154 382170 201250 382226
rect 201306 382170 201374 382226
rect 201430 382170 201498 382226
rect 201554 382170 201622 382226
rect 201678 382170 201774 382226
rect 201154 382102 201774 382170
rect 201154 382046 201250 382102
rect 201306 382046 201374 382102
rect 201430 382046 201498 382102
rect 201554 382046 201622 382102
rect 201678 382046 201774 382102
rect 201154 381978 201774 382046
rect 201154 381922 201250 381978
rect 201306 381922 201374 381978
rect 201430 381922 201498 381978
rect 201554 381922 201622 381978
rect 201678 381922 201774 381978
rect 201154 364350 201774 381922
rect 201154 364294 201250 364350
rect 201306 364294 201374 364350
rect 201430 364294 201498 364350
rect 201554 364294 201622 364350
rect 201678 364294 201774 364350
rect 201154 364226 201774 364294
rect 201154 364170 201250 364226
rect 201306 364170 201374 364226
rect 201430 364170 201498 364226
rect 201554 364170 201622 364226
rect 201678 364170 201774 364226
rect 201154 364102 201774 364170
rect 201154 364046 201250 364102
rect 201306 364046 201374 364102
rect 201430 364046 201498 364102
rect 201554 364046 201622 364102
rect 201678 364046 201774 364102
rect 201154 363978 201774 364046
rect 201154 363922 201250 363978
rect 201306 363922 201374 363978
rect 201430 363922 201498 363978
rect 201554 363922 201622 363978
rect 201678 363922 201774 363978
rect 201154 346350 201774 363922
rect 201154 346294 201250 346350
rect 201306 346294 201374 346350
rect 201430 346294 201498 346350
rect 201554 346294 201622 346350
rect 201678 346294 201774 346350
rect 201154 346226 201774 346294
rect 201154 346170 201250 346226
rect 201306 346170 201374 346226
rect 201430 346170 201498 346226
rect 201554 346170 201622 346226
rect 201678 346170 201774 346226
rect 201154 346102 201774 346170
rect 201154 346046 201250 346102
rect 201306 346046 201374 346102
rect 201430 346046 201498 346102
rect 201554 346046 201622 346102
rect 201678 346046 201774 346102
rect 201154 345978 201774 346046
rect 201154 345922 201250 345978
rect 201306 345922 201374 345978
rect 201430 345922 201498 345978
rect 201554 345922 201622 345978
rect 201678 345922 201774 345978
rect 201154 328350 201774 345922
rect 201154 328294 201250 328350
rect 201306 328294 201374 328350
rect 201430 328294 201498 328350
rect 201554 328294 201622 328350
rect 201678 328294 201774 328350
rect 201154 328226 201774 328294
rect 201154 328170 201250 328226
rect 201306 328170 201374 328226
rect 201430 328170 201498 328226
rect 201554 328170 201622 328226
rect 201678 328170 201774 328226
rect 201154 328102 201774 328170
rect 201154 328046 201250 328102
rect 201306 328046 201374 328102
rect 201430 328046 201498 328102
rect 201554 328046 201622 328102
rect 201678 328046 201774 328102
rect 201154 327978 201774 328046
rect 201154 327922 201250 327978
rect 201306 327922 201374 327978
rect 201430 327922 201498 327978
rect 201554 327922 201622 327978
rect 201678 327922 201774 327978
rect 198156 315140 198212 315150
rect 198044 310100 198100 310110
rect 197708 300804 197764 300814
rect 197708 158900 197764 300748
rect 198044 168644 198100 310044
rect 198156 305844 198212 315084
rect 198156 305778 198212 305788
rect 199612 313348 199668 313358
rect 198044 168578 198100 168588
rect 199052 305172 199108 305182
rect 198268 159684 198324 159694
rect 197708 158834 197764 158844
rect 197932 158900 197988 158910
rect 197932 148708 197988 158844
rect 198156 154644 198212 154654
rect 197932 148642 197988 148652
rect 198044 154308 198100 154318
rect 198044 150948 198100 154252
rect 198156 152404 198212 154588
rect 198156 152338 198212 152348
rect 197596 68674 197652 68684
rect 197484 7298 197540 7308
rect 195916 3938 195972 3948
rect 198044 980 198100 150892
rect 198268 144676 198324 159628
rect 198828 158004 198884 158014
rect 198828 145348 198884 157948
rect 198828 145282 198884 145292
rect 198268 144610 198324 144620
rect 198268 129332 198324 129342
rect 198268 104132 198324 129276
rect 199052 129332 199108 305116
rect 199612 173068 199668 313292
rect 199388 173012 199668 173068
rect 201154 310350 201774 327922
rect 201154 310294 201250 310350
rect 201306 310294 201374 310350
rect 201430 310294 201498 310350
rect 201554 310294 201622 310350
rect 201678 310294 201774 310350
rect 201154 310226 201774 310294
rect 201154 310170 201250 310226
rect 201306 310170 201374 310226
rect 201430 310170 201498 310226
rect 201554 310170 201622 310226
rect 201678 310170 201774 310226
rect 201154 310102 201774 310170
rect 201154 310046 201250 310102
rect 201306 310046 201374 310102
rect 201430 310046 201498 310102
rect 201554 310046 201622 310102
rect 201678 310046 201774 310102
rect 201154 309978 201774 310046
rect 201154 309922 201250 309978
rect 201306 309922 201374 309978
rect 201430 309922 201498 309978
rect 201554 309922 201622 309978
rect 201678 309922 201774 309978
rect 201154 292350 201774 309922
rect 201154 292294 201250 292350
rect 201306 292294 201374 292350
rect 201430 292294 201498 292350
rect 201554 292294 201622 292350
rect 201678 292294 201774 292350
rect 201154 292226 201774 292294
rect 201154 292170 201250 292226
rect 201306 292170 201374 292226
rect 201430 292170 201498 292226
rect 201554 292170 201622 292226
rect 201678 292170 201774 292226
rect 201154 292102 201774 292170
rect 201154 292046 201250 292102
rect 201306 292046 201374 292102
rect 201430 292046 201498 292102
rect 201554 292046 201622 292102
rect 201678 292046 201774 292102
rect 201154 291978 201774 292046
rect 201154 291922 201250 291978
rect 201306 291922 201374 291978
rect 201430 291922 201498 291978
rect 201554 291922 201622 291978
rect 201678 291922 201774 291978
rect 201154 274350 201774 291922
rect 201154 274294 201250 274350
rect 201306 274294 201374 274350
rect 201430 274294 201498 274350
rect 201554 274294 201622 274350
rect 201678 274294 201774 274350
rect 201154 274226 201774 274294
rect 201154 274170 201250 274226
rect 201306 274170 201374 274226
rect 201430 274170 201498 274226
rect 201554 274170 201622 274226
rect 201678 274170 201774 274226
rect 201154 274102 201774 274170
rect 201154 274046 201250 274102
rect 201306 274046 201374 274102
rect 201430 274046 201498 274102
rect 201554 274046 201622 274102
rect 201678 274046 201774 274102
rect 201154 273978 201774 274046
rect 201154 273922 201250 273978
rect 201306 273922 201374 273978
rect 201430 273922 201498 273978
rect 201554 273922 201622 273978
rect 201678 273922 201774 273978
rect 201154 256350 201774 273922
rect 201154 256294 201250 256350
rect 201306 256294 201374 256350
rect 201430 256294 201498 256350
rect 201554 256294 201622 256350
rect 201678 256294 201774 256350
rect 201154 256226 201774 256294
rect 201154 256170 201250 256226
rect 201306 256170 201374 256226
rect 201430 256170 201498 256226
rect 201554 256170 201622 256226
rect 201678 256170 201774 256226
rect 201154 256102 201774 256170
rect 201154 256046 201250 256102
rect 201306 256046 201374 256102
rect 201430 256046 201498 256102
rect 201554 256046 201622 256102
rect 201678 256046 201774 256102
rect 201154 255978 201774 256046
rect 201154 255922 201250 255978
rect 201306 255922 201374 255978
rect 201430 255922 201498 255978
rect 201554 255922 201622 255978
rect 201678 255922 201774 255978
rect 201154 238350 201774 255922
rect 201154 238294 201250 238350
rect 201306 238294 201374 238350
rect 201430 238294 201498 238350
rect 201554 238294 201622 238350
rect 201678 238294 201774 238350
rect 201154 238226 201774 238294
rect 201154 238170 201250 238226
rect 201306 238170 201374 238226
rect 201430 238170 201498 238226
rect 201554 238170 201622 238226
rect 201678 238170 201774 238226
rect 201154 238102 201774 238170
rect 201154 238046 201250 238102
rect 201306 238046 201374 238102
rect 201430 238046 201498 238102
rect 201554 238046 201622 238102
rect 201678 238046 201774 238102
rect 201154 237978 201774 238046
rect 201154 237922 201250 237978
rect 201306 237922 201374 237978
rect 201430 237922 201498 237978
rect 201554 237922 201622 237978
rect 201678 237922 201774 237978
rect 201154 220350 201774 237922
rect 201154 220294 201250 220350
rect 201306 220294 201374 220350
rect 201430 220294 201498 220350
rect 201554 220294 201622 220350
rect 201678 220294 201774 220350
rect 201154 220226 201774 220294
rect 201154 220170 201250 220226
rect 201306 220170 201374 220226
rect 201430 220170 201498 220226
rect 201554 220170 201622 220226
rect 201678 220170 201774 220226
rect 201154 220102 201774 220170
rect 201154 220046 201250 220102
rect 201306 220046 201374 220102
rect 201430 220046 201498 220102
rect 201554 220046 201622 220102
rect 201678 220046 201774 220102
rect 201154 219978 201774 220046
rect 201154 219922 201250 219978
rect 201306 219922 201374 219978
rect 201430 219922 201498 219978
rect 201554 219922 201622 219978
rect 201678 219922 201774 219978
rect 201154 202350 201774 219922
rect 201154 202294 201250 202350
rect 201306 202294 201374 202350
rect 201430 202294 201498 202350
rect 201554 202294 201622 202350
rect 201678 202294 201774 202350
rect 201154 202226 201774 202294
rect 201154 202170 201250 202226
rect 201306 202170 201374 202226
rect 201430 202170 201498 202226
rect 201554 202170 201622 202226
rect 201678 202170 201774 202226
rect 201154 202102 201774 202170
rect 201154 202046 201250 202102
rect 201306 202046 201374 202102
rect 201430 202046 201498 202102
rect 201554 202046 201622 202102
rect 201678 202046 201774 202102
rect 201154 201978 201774 202046
rect 201154 201922 201250 201978
rect 201306 201922 201374 201978
rect 201430 201922 201498 201978
rect 201554 201922 201622 201978
rect 201678 201922 201774 201978
rect 201154 184350 201774 201922
rect 201154 184294 201250 184350
rect 201306 184294 201374 184350
rect 201430 184294 201498 184350
rect 201554 184294 201622 184350
rect 201678 184294 201774 184350
rect 201154 184226 201774 184294
rect 201154 184170 201250 184226
rect 201306 184170 201374 184226
rect 201430 184170 201498 184226
rect 201554 184170 201622 184226
rect 201678 184170 201774 184226
rect 201154 184102 201774 184170
rect 201154 184046 201250 184102
rect 201306 184046 201374 184102
rect 201430 184046 201498 184102
rect 201554 184046 201622 184102
rect 201678 184046 201774 184102
rect 201154 183978 201774 184046
rect 201154 183922 201250 183978
rect 201306 183922 201374 183978
rect 201430 183922 201498 183978
rect 201554 183922 201622 183978
rect 201678 183922 201774 183978
rect 199388 169092 199444 173012
rect 199388 169026 199444 169036
rect 201154 166350 201774 183922
rect 201154 166294 201250 166350
rect 201306 166294 201374 166350
rect 201430 166294 201498 166350
rect 201554 166294 201622 166350
rect 201678 166294 201774 166350
rect 201154 166226 201774 166294
rect 201154 166170 201250 166226
rect 201306 166170 201374 166226
rect 201430 166170 201498 166226
rect 201554 166170 201622 166226
rect 201678 166170 201774 166226
rect 201154 166102 201774 166170
rect 201154 166046 201250 166102
rect 201306 166046 201374 166102
rect 201430 166046 201498 166102
rect 201554 166046 201622 166102
rect 201678 166046 201774 166102
rect 201154 165978 201774 166046
rect 201154 165922 201250 165978
rect 201306 165922 201374 165978
rect 201430 165922 201498 165978
rect 201554 165922 201622 165978
rect 201678 165922 201774 165978
rect 199612 157108 199668 157118
rect 199052 129266 199108 129276
rect 199164 144676 199220 144686
rect 198268 104066 198324 104076
rect 199052 117796 199108 117806
rect 198940 4340 198996 4350
rect 198940 3780 198996 4284
rect 198940 3714 198996 3724
rect 199052 3332 199108 117740
rect 199164 6356 199220 144620
rect 199388 138740 199444 138750
rect 199612 138740 199668 157052
rect 199836 155988 199892 155998
rect 199444 138684 199668 138740
rect 199724 152516 199780 152526
rect 199388 138674 199444 138684
rect 199276 131124 199332 131134
rect 199276 10052 199332 131068
rect 199388 121044 199444 121054
rect 199444 120988 199556 121044
rect 199388 120978 199444 120988
rect 199276 9986 199332 9996
rect 199500 9604 199556 120988
rect 199500 9538 199556 9548
rect 199164 6290 199220 6300
rect 199724 6020 199780 152460
rect 199724 5954 199780 5964
rect 199836 4900 199892 155932
rect 199836 4834 199892 4844
rect 201154 148350 201774 165922
rect 201154 148294 201250 148350
rect 201306 148294 201374 148350
rect 201430 148294 201498 148350
rect 201554 148294 201622 148350
rect 201678 148294 201774 148350
rect 201154 148226 201774 148294
rect 201154 148170 201250 148226
rect 201306 148170 201374 148226
rect 201430 148170 201498 148226
rect 201554 148170 201622 148226
rect 201678 148170 201774 148226
rect 201154 148102 201774 148170
rect 201154 148046 201250 148102
rect 201306 148046 201374 148102
rect 201430 148046 201498 148102
rect 201554 148046 201622 148102
rect 201678 148046 201774 148102
rect 201154 147978 201774 148046
rect 201154 147922 201250 147978
rect 201306 147922 201374 147978
rect 201430 147922 201498 147978
rect 201554 147922 201622 147978
rect 201678 147922 201774 147978
rect 201154 130350 201774 147922
rect 201154 130294 201250 130350
rect 201306 130294 201374 130350
rect 201430 130294 201498 130350
rect 201554 130294 201622 130350
rect 201678 130294 201774 130350
rect 201154 130226 201774 130294
rect 201154 130170 201250 130226
rect 201306 130170 201374 130226
rect 201430 130170 201498 130226
rect 201554 130170 201622 130226
rect 201678 130170 201774 130226
rect 201154 130102 201774 130170
rect 201154 130046 201250 130102
rect 201306 130046 201374 130102
rect 201430 130046 201498 130102
rect 201554 130046 201622 130102
rect 201678 130046 201774 130102
rect 201154 129978 201774 130046
rect 201154 129922 201250 129978
rect 201306 129922 201374 129978
rect 201430 129922 201498 129978
rect 201554 129922 201622 129978
rect 201678 129922 201774 129978
rect 201154 112350 201774 129922
rect 201154 112294 201250 112350
rect 201306 112294 201374 112350
rect 201430 112294 201498 112350
rect 201554 112294 201622 112350
rect 201678 112294 201774 112350
rect 201154 112226 201774 112294
rect 201154 112170 201250 112226
rect 201306 112170 201374 112226
rect 201430 112170 201498 112226
rect 201554 112170 201622 112226
rect 201678 112170 201774 112226
rect 201154 112102 201774 112170
rect 201154 112046 201250 112102
rect 201306 112046 201374 112102
rect 201430 112046 201498 112102
rect 201554 112046 201622 112102
rect 201678 112046 201774 112102
rect 201154 111978 201774 112046
rect 201154 111922 201250 111978
rect 201306 111922 201374 111978
rect 201430 111922 201498 111978
rect 201554 111922 201622 111978
rect 201678 111922 201774 111978
rect 201154 94350 201774 111922
rect 201154 94294 201250 94350
rect 201306 94294 201374 94350
rect 201430 94294 201498 94350
rect 201554 94294 201622 94350
rect 201678 94294 201774 94350
rect 201154 94226 201774 94294
rect 201154 94170 201250 94226
rect 201306 94170 201374 94226
rect 201430 94170 201498 94226
rect 201554 94170 201622 94226
rect 201678 94170 201774 94226
rect 201154 94102 201774 94170
rect 201154 94046 201250 94102
rect 201306 94046 201374 94102
rect 201430 94046 201498 94102
rect 201554 94046 201622 94102
rect 201678 94046 201774 94102
rect 201154 93978 201774 94046
rect 201154 93922 201250 93978
rect 201306 93922 201374 93978
rect 201430 93922 201498 93978
rect 201554 93922 201622 93978
rect 201678 93922 201774 93978
rect 201154 76350 201774 93922
rect 201154 76294 201250 76350
rect 201306 76294 201374 76350
rect 201430 76294 201498 76350
rect 201554 76294 201622 76350
rect 201678 76294 201774 76350
rect 201154 76226 201774 76294
rect 201154 76170 201250 76226
rect 201306 76170 201374 76226
rect 201430 76170 201498 76226
rect 201554 76170 201622 76226
rect 201678 76170 201774 76226
rect 201154 76102 201774 76170
rect 201154 76046 201250 76102
rect 201306 76046 201374 76102
rect 201430 76046 201498 76102
rect 201554 76046 201622 76102
rect 201678 76046 201774 76102
rect 201154 75978 201774 76046
rect 201154 75922 201250 75978
rect 201306 75922 201374 75978
rect 201430 75922 201498 75978
rect 201554 75922 201622 75978
rect 201678 75922 201774 75978
rect 201154 58350 201774 75922
rect 201154 58294 201250 58350
rect 201306 58294 201374 58350
rect 201430 58294 201498 58350
rect 201554 58294 201622 58350
rect 201678 58294 201774 58350
rect 201154 58226 201774 58294
rect 201154 58170 201250 58226
rect 201306 58170 201374 58226
rect 201430 58170 201498 58226
rect 201554 58170 201622 58226
rect 201678 58170 201774 58226
rect 201154 58102 201774 58170
rect 201154 58046 201250 58102
rect 201306 58046 201374 58102
rect 201430 58046 201498 58102
rect 201554 58046 201622 58102
rect 201678 58046 201774 58102
rect 201154 57978 201774 58046
rect 201154 57922 201250 57978
rect 201306 57922 201374 57978
rect 201430 57922 201498 57978
rect 201554 57922 201622 57978
rect 201678 57922 201774 57978
rect 201154 40350 201774 57922
rect 201154 40294 201250 40350
rect 201306 40294 201374 40350
rect 201430 40294 201498 40350
rect 201554 40294 201622 40350
rect 201678 40294 201774 40350
rect 201154 40226 201774 40294
rect 201154 40170 201250 40226
rect 201306 40170 201374 40226
rect 201430 40170 201498 40226
rect 201554 40170 201622 40226
rect 201678 40170 201774 40226
rect 201154 40102 201774 40170
rect 201154 40046 201250 40102
rect 201306 40046 201374 40102
rect 201430 40046 201498 40102
rect 201554 40046 201622 40102
rect 201678 40046 201774 40102
rect 201154 39978 201774 40046
rect 201154 39922 201250 39978
rect 201306 39922 201374 39978
rect 201430 39922 201498 39978
rect 201554 39922 201622 39978
rect 201678 39922 201774 39978
rect 201154 22350 201774 39922
rect 201154 22294 201250 22350
rect 201306 22294 201374 22350
rect 201430 22294 201498 22350
rect 201554 22294 201622 22350
rect 201678 22294 201774 22350
rect 201154 22226 201774 22294
rect 201154 22170 201250 22226
rect 201306 22170 201374 22226
rect 201430 22170 201498 22226
rect 201554 22170 201622 22226
rect 201678 22170 201774 22226
rect 201154 22102 201774 22170
rect 201154 22046 201250 22102
rect 201306 22046 201374 22102
rect 201430 22046 201498 22102
rect 201554 22046 201622 22102
rect 201678 22046 201774 22102
rect 201154 21978 201774 22046
rect 201154 21922 201250 21978
rect 201306 21922 201374 21978
rect 201430 21922 201498 21978
rect 201554 21922 201622 21978
rect 201678 21922 201774 21978
rect 199052 3266 199108 3276
rect 201154 4350 201774 21922
rect 201154 4294 201250 4350
rect 201306 4294 201374 4350
rect 201430 4294 201498 4350
rect 201554 4294 201622 4350
rect 201678 4294 201774 4350
rect 201154 4226 201774 4294
rect 201154 4170 201250 4226
rect 201306 4170 201374 4226
rect 201430 4170 201498 4226
rect 201554 4170 201622 4226
rect 201678 4170 201774 4226
rect 201154 4102 201774 4170
rect 201154 4046 201250 4102
rect 201306 4046 201374 4102
rect 201430 4046 201498 4102
rect 201554 4046 201622 4102
rect 201678 4046 201774 4102
rect 201154 3978 201774 4046
rect 201154 3922 201250 3978
rect 201306 3922 201374 3978
rect 201430 3922 201498 3978
rect 201554 3922 201622 3978
rect 201678 3922 201774 3978
rect 198044 914 198100 924
rect 186874 -1176 186970 -1120
rect 187026 -1176 187094 -1120
rect 187150 -1176 187218 -1120
rect 187274 -1176 187342 -1120
rect 187398 -1176 187494 -1120
rect 186874 -1244 187494 -1176
rect 186874 -1300 186970 -1244
rect 187026 -1300 187094 -1244
rect 187150 -1300 187218 -1244
rect 187274 -1300 187342 -1244
rect 187398 -1300 187494 -1244
rect 186874 -1368 187494 -1300
rect 186874 -1424 186970 -1368
rect 187026 -1424 187094 -1368
rect 187150 -1424 187218 -1368
rect 187274 -1424 187342 -1368
rect 187398 -1424 187494 -1368
rect 186874 -1492 187494 -1424
rect 186874 -1548 186970 -1492
rect 187026 -1548 187094 -1492
rect 187150 -1548 187218 -1492
rect 187274 -1548 187342 -1492
rect 187398 -1548 187494 -1492
rect 186874 -1644 187494 -1548
rect 201154 -160 201774 3922
rect 201154 -216 201250 -160
rect 201306 -216 201374 -160
rect 201430 -216 201498 -160
rect 201554 -216 201622 -160
rect 201678 -216 201774 -160
rect 201154 -284 201774 -216
rect 201154 -340 201250 -284
rect 201306 -340 201374 -284
rect 201430 -340 201498 -284
rect 201554 -340 201622 -284
rect 201678 -340 201774 -284
rect 201154 -408 201774 -340
rect 201154 -464 201250 -408
rect 201306 -464 201374 -408
rect 201430 -464 201498 -408
rect 201554 -464 201622 -408
rect 201678 -464 201774 -408
rect 201154 -532 201774 -464
rect 201154 -588 201250 -532
rect 201306 -588 201374 -532
rect 201430 -588 201498 -532
rect 201554 -588 201622 -532
rect 201678 -588 201774 -532
rect 201154 -1644 201774 -588
rect 204874 598172 205494 598268
rect 204874 598116 204970 598172
rect 205026 598116 205094 598172
rect 205150 598116 205218 598172
rect 205274 598116 205342 598172
rect 205398 598116 205494 598172
rect 204874 598048 205494 598116
rect 204874 597992 204970 598048
rect 205026 597992 205094 598048
rect 205150 597992 205218 598048
rect 205274 597992 205342 598048
rect 205398 597992 205494 598048
rect 204874 597924 205494 597992
rect 204874 597868 204970 597924
rect 205026 597868 205094 597924
rect 205150 597868 205218 597924
rect 205274 597868 205342 597924
rect 205398 597868 205494 597924
rect 204874 597800 205494 597868
rect 204874 597744 204970 597800
rect 205026 597744 205094 597800
rect 205150 597744 205218 597800
rect 205274 597744 205342 597800
rect 205398 597744 205494 597800
rect 204874 586350 205494 597744
rect 204874 586294 204970 586350
rect 205026 586294 205094 586350
rect 205150 586294 205218 586350
rect 205274 586294 205342 586350
rect 205398 586294 205494 586350
rect 204874 586226 205494 586294
rect 204874 586170 204970 586226
rect 205026 586170 205094 586226
rect 205150 586170 205218 586226
rect 205274 586170 205342 586226
rect 205398 586170 205494 586226
rect 204874 586102 205494 586170
rect 204874 586046 204970 586102
rect 205026 586046 205094 586102
rect 205150 586046 205218 586102
rect 205274 586046 205342 586102
rect 205398 586046 205494 586102
rect 204874 585978 205494 586046
rect 204874 585922 204970 585978
rect 205026 585922 205094 585978
rect 205150 585922 205218 585978
rect 205274 585922 205342 585978
rect 205398 585922 205494 585978
rect 204874 568350 205494 585922
rect 204874 568294 204970 568350
rect 205026 568294 205094 568350
rect 205150 568294 205218 568350
rect 205274 568294 205342 568350
rect 205398 568294 205494 568350
rect 204874 568226 205494 568294
rect 204874 568170 204970 568226
rect 205026 568170 205094 568226
rect 205150 568170 205218 568226
rect 205274 568170 205342 568226
rect 205398 568170 205494 568226
rect 204874 568102 205494 568170
rect 204874 568046 204970 568102
rect 205026 568046 205094 568102
rect 205150 568046 205218 568102
rect 205274 568046 205342 568102
rect 205398 568046 205494 568102
rect 204874 567978 205494 568046
rect 204874 567922 204970 567978
rect 205026 567922 205094 567978
rect 205150 567922 205218 567978
rect 205274 567922 205342 567978
rect 205398 567922 205494 567978
rect 204874 550350 205494 567922
rect 204874 550294 204970 550350
rect 205026 550294 205094 550350
rect 205150 550294 205218 550350
rect 205274 550294 205342 550350
rect 205398 550294 205494 550350
rect 204874 550226 205494 550294
rect 204874 550170 204970 550226
rect 205026 550170 205094 550226
rect 205150 550170 205218 550226
rect 205274 550170 205342 550226
rect 205398 550170 205494 550226
rect 204874 550102 205494 550170
rect 204874 550046 204970 550102
rect 205026 550046 205094 550102
rect 205150 550046 205218 550102
rect 205274 550046 205342 550102
rect 205398 550046 205494 550102
rect 204874 549978 205494 550046
rect 204874 549922 204970 549978
rect 205026 549922 205094 549978
rect 205150 549922 205218 549978
rect 205274 549922 205342 549978
rect 205398 549922 205494 549978
rect 204874 532350 205494 549922
rect 204874 532294 204970 532350
rect 205026 532294 205094 532350
rect 205150 532294 205218 532350
rect 205274 532294 205342 532350
rect 205398 532294 205494 532350
rect 204874 532226 205494 532294
rect 204874 532170 204970 532226
rect 205026 532170 205094 532226
rect 205150 532170 205218 532226
rect 205274 532170 205342 532226
rect 205398 532170 205494 532226
rect 204874 532102 205494 532170
rect 204874 532046 204970 532102
rect 205026 532046 205094 532102
rect 205150 532046 205218 532102
rect 205274 532046 205342 532102
rect 205398 532046 205494 532102
rect 204874 531978 205494 532046
rect 204874 531922 204970 531978
rect 205026 531922 205094 531978
rect 205150 531922 205218 531978
rect 205274 531922 205342 531978
rect 205398 531922 205494 531978
rect 204874 514350 205494 531922
rect 204874 514294 204970 514350
rect 205026 514294 205094 514350
rect 205150 514294 205218 514350
rect 205274 514294 205342 514350
rect 205398 514294 205494 514350
rect 204874 514226 205494 514294
rect 204874 514170 204970 514226
rect 205026 514170 205094 514226
rect 205150 514170 205218 514226
rect 205274 514170 205342 514226
rect 205398 514170 205494 514226
rect 204874 514102 205494 514170
rect 204874 514046 204970 514102
rect 205026 514046 205094 514102
rect 205150 514046 205218 514102
rect 205274 514046 205342 514102
rect 205398 514046 205494 514102
rect 204874 513978 205494 514046
rect 204874 513922 204970 513978
rect 205026 513922 205094 513978
rect 205150 513922 205218 513978
rect 205274 513922 205342 513978
rect 205398 513922 205494 513978
rect 204874 496350 205494 513922
rect 204874 496294 204970 496350
rect 205026 496294 205094 496350
rect 205150 496294 205218 496350
rect 205274 496294 205342 496350
rect 205398 496294 205494 496350
rect 204874 496226 205494 496294
rect 204874 496170 204970 496226
rect 205026 496170 205094 496226
rect 205150 496170 205218 496226
rect 205274 496170 205342 496226
rect 205398 496170 205494 496226
rect 204874 496102 205494 496170
rect 204874 496046 204970 496102
rect 205026 496046 205094 496102
rect 205150 496046 205218 496102
rect 205274 496046 205342 496102
rect 205398 496046 205494 496102
rect 204874 495978 205494 496046
rect 204874 495922 204970 495978
rect 205026 495922 205094 495978
rect 205150 495922 205218 495978
rect 205274 495922 205342 495978
rect 205398 495922 205494 495978
rect 204874 478350 205494 495922
rect 204874 478294 204970 478350
rect 205026 478294 205094 478350
rect 205150 478294 205218 478350
rect 205274 478294 205342 478350
rect 205398 478294 205494 478350
rect 204874 478226 205494 478294
rect 204874 478170 204970 478226
rect 205026 478170 205094 478226
rect 205150 478170 205218 478226
rect 205274 478170 205342 478226
rect 205398 478170 205494 478226
rect 204874 478102 205494 478170
rect 204874 478046 204970 478102
rect 205026 478046 205094 478102
rect 205150 478046 205218 478102
rect 205274 478046 205342 478102
rect 205398 478046 205494 478102
rect 204874 477978 205494 478046
rect 204874 477922 204970 477978
rect 205026 477922 205094 477978
rect 205150 477922 205218 477978
rect 205274 477922 205342 477978
rect 205398 477922 205494 477978
rect 204874 460350 205494 477922
rect 204874 460294 204970 460350
rect 205026 460294 205094 460350
rect 205150 460294 205218 460350
rect 205274 460294 205342 460350
rect 205398 460294 205494 460350
rect 204874 460226 205494 460294
rect 204874 460170 204970 460226
rect 205026 460170 205094 460226
rect 205150 460170 205218 460226
rect 205274 460170 205342 460226
rect 205398 460170 205494 460226
rect 204874 460102 205494 460170
rect 204874 460046 204970 460102
rect 205026 460046 205094 460102
rect 205150 460046 205218 460102
rect 205274 460046 205342 460102
rect 205398 460046 205494 460102
rect 204874 459978 205494 460046
rect 204874 459922 204970 459978
rect 205026 459922 205094 459978
rect 205150 459922 205218 459978
rect 205274 459922 205342 459978
rect 205398 459922 205494 459978
rect 204874 442350 205494 459922
rect 219154 597212 219774 598268
rect 219154 597156 219250 597212
rect 219306 597156 219374 597212
rect 219430 597156 219498 597212
rect 219554 597156 219622 597212
rect 219678 597156 219774 597212
rect 219154 597088 219774 597156
rect 219154 597032 219250 597088
rect 219306 597032 219374 597088
rect 219430 597032 219498 597088
rect 219554 597032 219622 597088
rect 219678 597032 219774 597088
rect 219154 596964 219774 597032
rect 219154 596908 219250 596964
rect 219306 596908 219374 596964
rect 219430 596908 219498 596964
rect 219554 596908 219622 596964
rect 219678 596908 219774 596964
rect 219154 596840 219774 596908
rect 219154 596784 219250 596840
rect 219306 596784 219374 596840
rect 219430 596784 219498 596840
rect 219554 596784 219622 596840
rect 219678 596784 219774 596840
rect 219154 580350 219774 596784
rect 219154 580294 219250 580350
rect 219306 580294 219374 580350
rect 219430 580294 219498 580350
rect 219554 580294 219622 580350
rect 219678 580294 219774 580350
rect 219154 580226 219774 580294
rect 219154 580170 219250 580226
rect 219306 580170 219374 580226
rect 219430 580170 219498 580226
rect 219554 580170 219622 580226
rect 219678 580170 219774 580226
rect 219154 580102 219774 580170
rect 219154 580046 219250 580102
rect 219306 580046 219374 580102
rect 219430 580046 219498 580102
rect 219554 580046 219622 580102
rect 219678 580046 219774 580102
rect 219154 579978 219774 580046
rect 219154 579922 219250 579978
rect 219306 579922 219374 579978
rect 219430 579922 219498 579978
rect 219554 579922 219622 579978
rect 219678 579922 219774 579978
rect 219154 562350 219774 579922
rect 219154 562294 219250 562350
rect 219306 562294 219374 562350
rect 219430 562294 219498 562350
rect 219554 562294 219622 562350
rect 219678 562294 219774 562350
rect 219154 562226 219774 562294
rect 219154 562170 219250 562226
rect 219306 562170 219374 562226
rect 219430 562170 219498 562226
rect 219554 562170 219622 562226
rect 219678 562170 219774 562226
rect 219154 562102 219774 562170
rect 219154 562046 219250 562102
rect 219306 562046 219374 562102
rect 219430 562046 219498 562102
rect 219554 562046 219622 562102
rect 219678 562046 219774 562102
rect 219154 561978 219774 562046
rect 219154 561922 219250 561978
rect 219306 561922 219374 561978
rect 219430 561922 219498 561978
rect 219554 561922 219622 561978
rect 219678 561922 219774 561978
rect 219154 544350 219774 561922
rect 219154 544294 219250 544350
rect 219306 544294 219374 544350
rect 219430 544294 219498 544350
rect 219554 544294 219622 544350
rect 219678 544294 219774 544350
rect 219154 544226 219774 544294
rect 219154 544170 219250 544226
rect 219306 544170 219374 544226
rect 219430 544170 219498 544226
rect 219554 544170 219622 544226
rect 219678 544170 219774 544226
rect 219154 544102 219774 544170
rect 219154 544046 219250 544102
rect 219306 544046 219374 544102
rect 219430 544046 219498 544102
rect 219554 544046 219622 544102
rect 219678 544046 219774 544102
rect 219154 543978 219774 544046
rect 219154 543922 219250 543978
rect 219306 543922 219374 543978
rect 219430 543922 219498 543978
rect 219554 543922 219622 543978
rect 219678 543922 219774 543978
rect 219154 526350 219774 543922
rect 219154 526294 219250 526350
rect 219306 526294 219374 526350
rect 219430 526294 219498 526350
rect 219554 526294 219622 526350
rect 219678 526294 219774 526350
rect 219154 526226 219774 526294
rect 219154 526170 219250 526226
rect 219306 526170 219374 526226
rect 219430 526170 219498 526226
rect 219554 526170 219622 526226
rect 219678 526170 219774 526226
rect 219154 526102 219774 526170
rect 219154 526046 219250 526102
rect 219306 526046 219374 526102
rect 219430 526046 219498 526102
rect 219554 526046 219622 526102
rect 219678 526046 219774 526102
rect 219154 525978 219774 526046
rect 219154 525922 219250 525978
rect 219306 525922 219374 525978
rect 219430 525922 219498 525978
rect 219554 525922 219622 525978
rect 219678 525922 219774 525978
rect 219154 508350 219774 525922
rect 219154 508294 219250 508350
rect 219306 508294 219374 508350
rect 219430 508294 219498 508350
rect 219554 508294 219622 508350
rect 219678 508294 219774 508350
rect 219154 508226 219774 508294
rect 219154 508170 219250 508226
rect 219306 508170 219374 508226
rect 219430 508170 219498 508226
rect 219554 508170 219622 508226
rect 219678 508170 219774 508226
rect 219154 508102 219774 508170
rect 219154 508046 219250 508102
rect 219306 508046 219374 508102
rect 219430 508046 219498 508102
rect 219554 508046 219622 508102
rect 219678 508046 219774 508102
rect 219154 507978 219774 508046
rect 219154 507922 219250 507978
rect 219306 507922 219374 507978
rect 219430 507922 219498 507978
rect 219554 507922 219622 507978
rect 219678 507922 219774 507978
rect 219154 490350 219774 507922
rect 219154 490294 219250 490350
rect 219306 490294 219374 490350
rect 219430 490294 219498 490350
rect 219554 490294 219622 490350
rect 219678 490294 219774 490350
rect 219154 490226 219774 490294
rect 219154 490170 219250 490226
rect 219306 490170 219374 490226
rect 219430 490170 219498 490226
rect 219554 490170 219622 490226
rect 219678 490170 219774 490226
rect 219154 490102 219774 490170
rect 219154 490046 219250 490102
rect 219306 490046 219374 490102
rect 219430 490046 219498 490102
rect 219554 490046 219622 490102
rect 219678 490046 219774 490102
rect 219154 489978 219774 490046
rect 219154 489922 219250 489978
rect 219306 489922 219374 489978
rect 219430 489922 219498 489978
rect 219554 489922 219622 489978
rect 219678 489922 219774 489978
rect 219154 472350 219774 489922
rect 219154 472294 219250 472350
rect 219306 472294 219374 472350
rect 219430 472294 219498 472350
rect 219554 472294 219622 472350
rect 219678 472294 219774 472350
rect 219154 472226 219774 472294
rect 219154 472170 219250 472226
rect 219306 472170 219374 472226
rect 219430 472170 219498 472226
rect 219554 472170 219622 472226
rect 219678 472170 219774 472226
rect 219154 472102 219774 472170
rect 219154 472046 219250 472102
rect 219306 472046 219374 472102
rect 219430 472046 219498 472102
rect 219554 472046 219622 472102
rect 219678 472046 219774 472102
rect 219154 471978 219774 472046
rect 219154 471922 219250 471978
rect 219306 471922 219374 471978
rect 219430 471922 219498 471978
rect 219554 471922 219622 471978
rect 219678 471922 219774 471978
rect 219154 458342 219774 471922
rect 222874 598172 223494 598268
rect 222874 598116 222970 598172
rect 223026 598116 223094 598172
rect 223150 598116 223218 598172
rect 223274 598116 223342 598172
rect 223398 598116 223494 598172
rect 222874 598048 223494 598116
rect 222874 597992 222970 598048
rect 223026 597992 223094 598048
rect 223150 597992 223218 598048
rect 223274 597992 223342 598048
rect 223398 597992 223494 598048
rect 222874 597924 223494 597992
rect 222874 597868 222970 597924
rect 223026 597868 223094 597924
rect 223150 597868 223218 597924
rect 223274 597868 223342 597924
rect 223398 597868 223494 597924
rect 222874 597800 223494 597868
rect 222874 597744 222970 597800
rect 223026 597744 223094 597800
rect 223150 597744 223218 597800
rect 223274 597744 223342 597800
rect 223398 597744 223494 597800
rect 222874 586350 223494 597744
rect 222874 586294 222970 586350
rect 223026 586294 223094 586350
rect 223150 586294 223218 586350
rect 223274 586294 223342 586350
rect 223398 586294 223494 586350
rect 222874 586226 223494 586294
rect 222874 586170 222970 586226
rect 223026 586170 223094 586226
rect 223150 586170 223218 586226
rect 223274 586170 223342 586226
rect 223398 586170 223494 586226
rect 222874 586102 223494 586170
rect 222874 586046 222970 586102
rect 223026 586046 223094 586102
rect 223150 586046 223218 586102
rect 223274 586046 223342 586102
rect 223398 586046 223494 586102
rect 222874 585978 223494 586046
rect 222874 585922 222970 585978
rect 223026 585922 223094 585978
rect 223150 585922 223218 585978
rect 223274 585922 223342 585978
rect 223398 585922 223494 585978
rect 222874 568350 223494 585922
rect 222874 568294 222970 568350
rect 223026 568294 223094 568350
rect 223150 568294 223218 568350
rect 223274 568294 223342 568350
rect 223398 568294 223494 568350
rect 222874 568226 223494 568294
rect 222874 568170 222970 568226
rect 223026 568170 223094 568226
rect 223150 568170 223218 568226
rect 223274 568170 223342 568226
rect 223398 568170 223494 568226
rect 222874 568102 223494 568170
rect 222874 568046 222970 568102
rect 223026 568046 223094 568102
rect 223150 568046 223218 568102
rect 223274 568046 223342 568102
rect 223398 568046 223494 568102
rect 222874 567978 223494 568046
rect 222874 567922 222970 567978
rect 223026 567922 223094 567978
rect 223150 567922 223218 567978
rect 223274 567922 223342 567978
rect 223398 567922 223494 567978
rect 222874 550350 223494 567922
rect 222874 550294 222970 550350
rect 223026 550294 223094 550350
rect 223150 550294 223218 550350
rect 223274 550294 223342 550350
rect 223398 550294 223494 550350
rect 222874 550226 223494 550294
rect 222874 550170 222970 550226
rect 223026 550170 223094 550226
rect 223150 550170 223218 550226
rect 223274 550170 223342 550226
rect 223398 550170 223494 550226
rect 222874 550102 223494 550170
rect 222874 550046 222970 550102
rect 223026 550046 223094 550102
rect 223150 550046 223218 550102
rect 223274 550046 223342 550102
rect 223398 550046 223494 550102
rect 222874 549978 223494 550046
rect 222874 549922 222970 549978
rect 223026 549922 223094 549978
rect 223150 549922 223218 549978
rect 223274 549922 223342 549978
rect 223398 549922 223494 549978
rect 222874 532350 223494 549922
rect 222874 532294 222970 532350
rect 223026 532294 223094 532350
rect 223150 532294 223218 532350
rect 223274 532294 223342 532350
rect 223398 532294 223494 532350
rect 222874 532226 223494 532294
rect 222874 532170 222970 532226
rect 223026 532170 223094 532226
rect 223150 532170 223218 532226
rect 223274 532170 223342 532226
rect 223398 532170 223494 532226
rect 222874 532102 223494 532170
rect 222874 532046 222970 532102
rect 223026 532046 223094 532102
rect 223150 532046 223218 532102
rect 223274 532046 223342 532102
rect 223398 532046 223494 532102
rect 222874 531978 223494 532046
rect 222874 531922 222970 531978
rect 223026 531922 223094 531978
rect 223150 531922 223218 531978
rect 223274 531922 223342 531978
rect 223398 531922 223494 531978
rect 222874 514350 223494 531922
rect 222874 514294 222970 514350
rect 223026 514294 223094 514350
rect 223150 514294 223218 514350
rect 223274 514294 223342 514350
rect 223398 514294 223494 514350
rect 222874 514226 223494 514294
rect 222874 514170 222970 514226
rect 223026 514170 223094 514226
rect 223150 514170 223218 514226
rect 223274 514170 223342 514226
rect 223398 514170 223494 514226
rect 222874 514102 223494 514170
rect 222874 514046 222970 514102
rect 223026 514046 223094 514102
rect 223150 514046 223218 514102
rect 223274 514046 223342 514102
rect 223398 514046 223494 514102
rect 222874 513978 223494 514046
rect 222874 513922 222970 513978
rect 223026 513922 223094 513978
rect 223150 513922 223218 513978
rect 223274 513922 223342 513978
rect 223398 513922 223494 513978
rect 222874 496350 223494 513922
rect 222874 496294 222970 496350
rect 223026 496294 223094 496350
rect 223150 496294 223218 496350
rect 223274 496294 223342 496350
rect 223398 496294 223494 496350
rect 222874 496226 223494 496294
rect 222874 496170 222970 496226
rect 223026 496170 223094 496226
rect 223150 496170 223218 496226
rect 223274 496170 223342 496226
rect 223398 496170 223494 496226
rect 222874 496102 223494 496170
rect 222874 496046 222970 496102
rect 223026 496046 223094 496102
rect 223150 496046 223218 496102
rect 223274 496046 223342 496102
rect 223398 496046 223494 496102
rect 222874 495978 223494 496046
rect 222874 495922 222970 495978
rect 223026 495922 223094 495978
rect 223150 495922 223218 495978
rect 223274 495922 223342 495978
rect 223398 495922 223494 495978
rect 222874 478350 223494 495922
rect 222874 478294 222970 478350
rect 223026 478294 223094 478350
rect 223150 478294 223218 478350
rect 223274 478294 223342 478350
rect 223398 478294 223494 478350
rect 222874 478226 223494 478294
rect 222874 478170 222970 478226
rect 223026 478170 223094 478226
rect 223150 478170 223218 478226
rect 223274 478170 223342 478226
rect 223398 478170 223494 478226
rect 222874 478102 223494 478170
rect 222874 478046 222970 478102
rect 223026 478046 223094 478102
rect 223150 478046 223218 478102
rect 223274 478046 223342 478102
rect 223398 478046 223494 478102
rect 222874 477978 223494 478046
rect 222874 477922 222970 477978
rect 223026 477922 223094 477978
rect 223150 477922 223218 477978
rect 223274 477922 223342 477978
rect 223398 477922 223494 477978
rect 222874 460350 223494 477922
rect 222874 460294 222970 460350
rect 223026 460294 223094 460350
rect 223150 460294 223218 460350
rect 223274 460294 223342 460350
rect 223398 460294 223494 460350
rect 222874 460226 223494 460294
rect 222874 460170 222970 460226
rect 223026 460170 223094 460226
rect 223150 460170 223218 460226
rect 223274 460170 223342 460226
rect 223398 460170 223494 460226
rect 222874 460102 223494 460170
rect 222874 460046 222970 460102
rect 223026 460046 223094 460102
rect 223150 460046 223218 460102
rect 223274 460046 223342 460102
rect 223398 460046 223494 460102
rect 222874 459978 223494 460046
rect 222874 459922 222970 459978
rect 223026 459922 223094 459978
rect 223150 459922 223218 459978
rect 223274 459922 223342 459978
rect 223398 459922 223494 459978
rect 222874 458342 223494 459922
rect 237154 597212 237774 598268
rect 237154 597156 237250 597212
rect 237306 597156 237374 597212
rect 237430 597156 237498 597212
rect 237554 597156 237622 597212
rect 237678 597156 237774 597212
rect 237154 597088 237774 597156
rect 237154 597032 237250 597088
rect 237306 597032 237374 597088
rect 237430 597032 237498 597088
rect 237554 597032 237622 597088
rect 237678 597032 237774 597088
rect 237154 596964 237774 597032
rect 237154 596908 237250 596964
rect 237306 596908 237374 596964
rect 237430 596908 237498 596964
rect 237554 596908 237622 596964
rect 237678 596908 237774 596964
rect 237154 596840 237774 596908
rect 237154 596784 237250 596840
rect 237306 596784 237374 596840
rect 237430 596784 237498 596840
rect 237554 596784 237622 596840
rect 237678 596784 237774 596840
rect 237154 580350 237774 596784
rect 237154 580294 237250 580350
rect 237306 580294 237374 580350
rect 237430 580294 237498 580350
rect 237554 580294 237622 580350
rect 237678 580294 237774 580350
rect 237154 580226 237774 580294
rect 237154 580170 237250 580226
rect 237306 580170 237374 580226
rect 237430 580170 237498 580226
rect 237554 580170 237622 580226
rect 237678 580170 237774 580226
rect 237154 580102 237774 580170
rect 237154 580046 237250 580102
rect 237306 580046 237374 580102
rect 237430 580046 237498 580102
rect 237554 580046 237622 580102
rect 237678 580046 237774 580102
rect 237154 579978 237774 580046
rect 237154 579922 237250 579978
rect 237306 579922 237374 579978
rect 237430 579922 237498 579978
rect 237554 579922 237622 579978
rect 237678 579922 237774 579978
rect 237154 562350 237774 579922
rect 237154 562294 237250 562350
rect 237306 562294 237374 562350
rect 237430 562294 237498 562350
rect 237554 562294 237622 562350
rect 237678 562294 237774 562350
rect 237154 562226 237774 562294
rect 237154 562170 237250 562226
rect 237306 562170 237374 562226
rect 237430 562170 237498 562226
rect 237554 562170 237622 562226
rect 237678 562170 237774 562226
rect 237154 562102 237774 562170
rect 237154 562046 237250 562102
rect 237306 562046 237374 562102
rect 237430 562046 237498 562102
rect 237554 562046 237622 562102
rect 237678 562046 237774 562102
rect 237154 561978 237774 562046
rect 237154 561922 237250 561978
rect 237306 561922 237374 561978
rect 237430 561922 237498 561978
rect 237554 561922 237622 561978
rect 237678 561922 237774 561978
rect 237154 544350 237774 561922
rect 237154 544294 237250 544350
rect 237306 544294 237374 544350
rect 237430 544294 237498 544350
rect 237554 544294 237622 544350
rect 237678 544294 237774 544350
rect 237154 544226 237774 544294
rect 237154 544170 237250 544226
rect 237306 544170 237374 544226
rect 237430 544170 237498 544226
rect 237554 544170 237622 544226
rect 237678 544170 237774 544226
rect 237154 544102 237774 544170
rect 237154 544046 237250 544102
rect 237306 544046 237374 544102
rect 237430 544046 237498 544102
rect 237554 544046 237622 544102
rect 237678 544046 237774 544102
rect 237154 543978 237774 544046
rect 237154 543922 237250 543978
rect 237306 543922 237374 543978
rect 237430 543922 237498 543978
rect 237554 543922 237622 543978
rect 237678 543922 237774 543978
rect 237154 526350 237774 543922
rect 237154 526294 237250 526350
rect 237306 526294 237374 526350
rect 237430 526294 237498 526350
rect 237554 526294 237622 526350
rect 237678 526294 237774 526350
rect 237154 526226 237774 526294
rect 237154 526170 237250 526226
rect 237306 526170 237374 526226
rect 237430 526170 237498 526226
rect 237554 526170 237622 526226
rect 237678 526170 237774 526226
rect 237154 526102 237774 526170
rect 237154 526046 237250 526102
rect 237306 526046 237374 526102
rect 237430 526046 237498 526102
rect 237554 526046 237622 526102
rect 237678 526046 237774 526102
rect 237154 525978 237774 526046
rect 237154 525922 237250 525978
rect 237306 525922 237374 525978
rect 237430 525922 237498 525978
rect 237554 525922 237622 525978
rect 237678 525922 237774 525978
rect 237154 508350 237774 525922
rect 237154 508294 237250 508350
rect 237306 508294 237374 508350
rect 237430 508294 237498 508350
rect 237554 508294 237622 508350
rect 237678 508294 237774 508350
rect 237154 508226 237774 508294
rect 237154 508170 237250 508226
rect 237306 508170 237374 508226
rect 237430 508170 237498 508226
rect 237554 508170 237622 508226
rect 237678 508170 237774 508226
rect 237154 508102 237774 508170
rect 237154 508046 237250 508102
rect 237306 508046 237374 508102
rect 237430 508046 237498 508102
rect 237554 508046 237622 508102
rect 237678 508046 237774 508102
rect 237154 507978 237774 508046
rect 237154 507922 237250 507978
rect 237306 507922 237374 507978
rect 237430 507922 237498 507978
rect 237554 507922 237622 507978
rect 237678 507922 237774 507978
rect 237154 490350 237774 507922
rect 237154 490294 237250 490350
rect 237306 490294 237374 490350
rect 237430 490294 237498 490350
rect 237554 490294 237622 490350
rect 237678 490294 237774 490350
rect 237154 490226 237774 490294
rect 237154 490170 237250 490226
rect 237306 490170 237374 490226
rect 237430 490170 237498 490226
rect 237554 490170 237622 490226
rect 237678 490170 237774 490226
rect 237154 490102 237774 490170
rect 237154 490046 237250 490102
rect 237306 490046 237374 490102
rect 237430 490046 237498 490102
rect 237554 490046 237622 490102
rect 237678 490046 237774 490102
rect 237154 489978 237774 490046
rect 237154 489922 237250 489978
rect 237306 489922 237374 489978
rect 237430 489922 237498 489978
rect 237554 489922 237622 489978
rect 237678 489922 237774 489978
rect 237154 472350 237774 489922
rect 237154 472294 237250 472350
rect 237306 472294 237374 472350
rect 237430 472294 237498 472350
rect 237554 472294 237622 472350
rect 237678 472294 237774 472350
rect 237154 472226 237774 472294
rect 237154 472170 237250 472226
rect 237306 472170 237374 472226
rect 237430 472170 237498 472226
rect 237554 472170 237622 472226
rect 237678 472170 237774 472226
rect 237154 472102 237774 472170
rect 237154 472046 237250 472102
rect 237306 472046 237374 472102
rect 237430 472046 237498 472102
rect 237554 472046 237622 472102
rect 237678 472046 237774 472102
rect 237154 471978 237774 472046
rect 237154 471922 237250 471978
rect 237306 471922 237374 471978
rect 237430 471922 237498 471978
rect 237554 471922 237622 471978
rect 237678 471922 237774 471978
rect 237154 458342 237774 471922
rect 240874 598172 241494 598268
rect 240874 598116 240970 598172
rect 241026 598116 241094 598172
rect 241150 598116 241218 598172
rect 241274 598116 241342 598172
rect 241398 598116 241494 598172
rect 240874 598048 241494 598116
rect 240874 597992 240970 598048
rect 241026 597992 241094 598048
rect 241150 597992 241218 598048
rect 241274 597992 241342 598048
rect 241398 597992 241494 598048
rect 240874 597924 241494 597992
rect 240874 597868 240970 597924
rect 241026 597868 241094 597924
rect 241150 597868 241218 597924
rect 241274 597868 241342 597924
rect 241398 597868 241494 597924
rect 240874 597800 241494 597868
rect 240874 597744 240970 597800
rect 241026 597744 241094 597800
rect 241150 597744 241218 597800
rect 241274 597744 241342 597800
rect 241398 597744 241494 597800
rect 240874 586350 241494 597744
rect 240874 586294 240970 586350
rect 241026 586294 241094 586350
rect 241150 586294 241218 586350
rect 241274 586294 241342 586350
rect 241398 586294 241494 586350
rect 240874 586226 241494 586294
rect 240874 586170 240970 586226
rect 241026 586170 241094 586226
rect 241150 586170 241218 586226
rect 241274 586170 241342 586226
rect 241398 586170 241494 586226
rect 240874 586102 241494 586170
rect 240874 586046 240970 586102
rect 241026 586046 241094 586102
rect 241150 586046 241218 586102
rect 241274 586046 241342 586102
rect 241398 586046 241494 586102
rect 240874 585978 241494 586046
rect 240874 585922 240970 585978
rect 241026 585922 241094 585978
rect 241150 585922 241218 585978
rect 241274 585922 241342 585978
rect 241398 585922 241494 585978
rect 240874 568350 241494 585922
rect 240874 568294 240970 568350
rect 241026 568294 241094 568350
rect 241150 568294 241218 568350
rect 241274 568294 241342 568350
rect 241398 568294 241494 568350
rect 240874 568226 241494 568294
rect 240874 568170 240970 568226
rect 241026 568170 241094 568226
rect 241150 568170 241218 568226
rect 241274 568170 241342 568226
rect 241398 568170 241494 568226
rect 240874 568102 241494 568170
rect 240874 568046 240970 568102
rect 241026 568046 241094 568102
rect 241150 568046 241218 568102
rect 241274 568046 241342 568102
rect 241398 568046 241494 568102
rect 240874 567978 241494 568046
rect 240874 567922 240970 567978
rect 241026 567922 241094 567978
rect 241150 567922 241218 567978
rect 241274 567922 241342 567978
rect 241398 567922 241494 567978
rect 240874 550350 241494 567922
rect 240874 550294 240970 550350
rect 241026 550294 241094 550350
rect 241150 550294 241218 550350
rect 241274 550294 241342 550350
rect 241398 550294 241494 550350
rect 240874 550226 241494 550294
rect 240874 550170 240970 550226
rect 241026 550170 241094 550226
rect 241150 550170 241218 550226
rect 241274 550170 241342 550226
rect 241398 550170 241494 550226
rect 240874 550102 241494 550170
rect 240874 550046 240970 550102
rect 241026 550046 241094 550102
rect 241150 550046 241218 550102
rect 241274 550046 241342 550102
rect 241398 550046 241494 550102
rect 240874 549978 241494 550046
rect 240874 549922 240970 549978
rect 241026 549922 241094 549978
rect 241150 549922 241218 549978
rect 241274 549922 241342 549978
rect 241398 549922 241494 549978
rect 240874 532350 241494 549922
rect 240874 532294 240970 532350
rect 241026 532294 241094 532350
rect 241150 532294 241218 532350
rect 241274 532294 241342 532350
rect 241398 532294 241494 532350
rect 240874 532226 241494 532294
rect 240874 532170 240970 532226
rect 241026 532170 241094 532226
rect 241150 532170 241218 532226
rect 241274 532170 241342 532226
rect 241398 532170 241494 532226
rect 240874 532102 241494 532170
rect 240874 532046 240970 532102
rect 241026 532046 241094 532102
rect 241150 532046 241218 532102
rect 241274 532046 241342 532102
rect 241398 532046 241494 532102
rect 240874 531978 241494 532046
rect 240874 531922 240970 531978
rect 241026 531922 241094 531978
rect 241150 531922 241218 531978
rect 241274 531922 241342 531978
rect 241398 531922 241494 531978
rect 240874 514350 241494 531922
rect 240874 514294 240970 514350
rect 241026 514294 241094 514350
rect 241150 514294 241218 514350
rect 241274 514294 241342 514350
rect 241398 514294 241494 514350
rect 240874 514226 241494 514294
rect 240874 514170 240970 514226
rect 241026 514170 241094 514226
rect 241150 514170 241218 514226
rect 241274 514170 241342 514226
rect 241398 514170 241494 514226
rect 240874 514102 241494 514170
rect 240874 514046 240970 514102
rect 241026 514046 241094 514102
rect 241150 514046 241218 514102
rect 241274 514046 241342 514102
rect 241398 514046 241494 514102
rect 240874 513978 241494 514046
rect 240874 513922 240970 513978
rect 241026 513922 241094 513978
rect 241150 513922 241218 513978
rect 241274 513922 241342 513978
rect 241398 513922 241494 513978
rect 240874 496350 241494 513922
rect 240874 496294 240970 496350
rect 241026 496294 241094 496350
rect 241150 496294 241218 496350
rect 241274 496294 241342 496350
rect 241398 496294 241494 496350
rect 240874 496226 241494 496294
rect 240874 496170 240970 496226
rect 241026 496170 241094 496226
rect 241150 496170 241218 496226
rect 241274 496170 241342 496226
rect 241398 496170 241494 496226
rect 240874 496102 241494 496170
rect 240874 496046 240970 496102
rect 241026 496046 241094 496102
rect 241150 496046 241218 496102
rect 241274 496046 241342 496102
rect 241398 496046 241494 496102
rect 240874 495978 241494 496046
rect 240874 495922 240970 495978
rect 241026 495922 241094 495978
rect 241150 495922 241218 495978
rect 241274 495922 241342 495978
rect 241398 495922 241494 495978
rect 240874 478350 241494 495922
rect 240874 478294 240970 478350
rect 241026 478294 241094 478350
rect 241150 478294 241218 478350
rect 241274 478294 241342 478350
rect 241398 478294 241494 478350
rect 240874 478226 241494 478294
rect 240874 478170 240970 478226
rect 241026 478170 241094 478226
rect 241150 478170 241218 478226
rect 241274 478170 241342 478226
rect 241398 478170 241494 478226
rect 240874 478102 241494 478170
rect 240874 478046 240970 478102
rect 241026 478046 241094 478102
rect 241150 478046 241218 478102
rect 241274 478046 241342 478102
rect 241398 478046 241494 478102
rect 240874 477978 241494 478046
rect 240874 477922 240970 477978
rect 241026 477922 241094 477978
rect 241150 477922 241218 477978
rect 241274 477922 241342 477978
rect 241398 477922 241494 477978
rect 240874 460350 241494 477922
rect 240874 460294 240970 460350
rect 241026 460294 241094 460350
rect 241150 460294 241218 460350
rect 241274 460294 241342 460350
rect 241398 460294 241494 460350
rect 240874 460226 241494 460294
rect 240874 460170 240970 460226
rect 241026 460170 241094 460226
rect 241150 460170 241218 460226
rect 241274 460170 241342 460226
rect 241398 460170 241494 460226
rect 240874 460102 241494 460170
rect 240874 460046 240970 460102
rect 241026 460046 241094 460102
rect 241150 460046 241218 460102
rect 241274 460046 241342 460102
rect 241398 460046 241494 460102
rect 240874 459978 241494 460046
rect 240874 459922 240970 459978
rect 241026 459922 241094 459978
rect 241150 459922 241218 459978
rect 241274 459922 241342 459978
rect 241398 459922 241494 459978
rect 240874 458342 241494 459922
rect 255154 597212 255774 598268
rect 255154 597156 255250 597212
rect 255306 597156 255374 597212
rect 255430 597156 255498 597212
rect 255554 597156 255622 597212
rect 255678 597156 255774 597212
rect 255154 597088 255774 597156
rect 255154 597032 255250 597088
rect 255306 597032 255374 597088
rect 255430 597032 255498 597088
rect 255554 597032 255622 597088
rect 255678 597032 255774 597088
rect 255154 596964 255774 597032
rect 255154 596908 255250 596964
rect 255306 596908 255374 596964
rect 255430 596908 255498 596964
rect 255554 596908 255622 596964
rect 255678 596908 255774 596964
rect 255154 596840 255774 596908
rect 255154 596784 255250 596840
rect 255306 596784 255374 596840
rect 255430 596784 255498 596840
rect 255554 596784 255622 596840
rect 255678 596784 255774 596840
rect 255154 580350 255774 596784
rect 255154 580294 255250 580350
rect 255306 580294 255374 580350
rect 255430 580294 255498 580350
rect 255554 580294 255622 580350
rect 255678 580294 255774 580350
rect 255154 580226 255774 580294
rect 255154 580170 255250 580226
rect 255306 580170 255374 580226
rect 255430 580170 255498 580226
rect 255554 580170 255622 580226
rect 255678 580170 255774 580226
rect 255154 580102 255774 580170
rect 255154 580046 255250 580102
rect 255306 580046 255374 580102
rect 255430 580046 255498 580102
rect 255554 580046 255622 580102
rect 255678 580046 255774 580102
rect 255154 579978 255774 580046
rect 255154 579922 255250 579978
rect 255306 579922 255374 579978
rect 255430 579922 255498 579978
rect 255554 579922 255622 579978
rect 255678 579922 255774 579978
rect 255154 562350 255774 579922
rect 255154 562294 255250 562350
rect 255306 562294 255374 562350
rect 255430 562294 255498 562350
rect 255554 562294 255622 562350
rect 255678 562294 255774 562350
rect 255154 562226 255774 562294
rect 255154 562170 255250 562226
rect 255306 562170 255374 562226
rect 255430 562170 255498 562226
rect 255554 562170 255622 562226
rect 255678 562170 255774 562226
rect 255154 562102 255774 562170
rect 255154 562046 255250 562102
rect 255306 562046 255374 562102
rect 255430 562046 255498 562102
rect 255554 562046 255622 562102
rect 255678 562046 255774 562102
rect 255154 561978 255774 562046
rect 255154 561922 255250 561978
rect 255306 561922 255374 561978
rect 255430 561922 255498 561978
rect 255554 561922 255622 561978
rect 255678 561922 255774 561978
rect 255154 544350 255774 561922
rect 255154 544294 255250 544350
rect 255306 544294 255374 544350
rect 255430 544294 255498 544350
rect 255554 544294 255622 544350
rect 255678 544294 255774 544350
rect 255154 544226 255774 544294
rect 255154 544170 255250 544226
rect 255306 544170 255374 544226
rect 255430 544170 255498 544226
rect 255554 544170 255622 544226
rect 255678 544170 255774 544226
rect 255154 544102 255774 544170
rect 255154 544046 255250 544102
rect 255306 544046 255374 544102
rect 255430 544046 255498 544102
rect 255554 544046 255622 544102
rect 255678 544046 255774 544102
rect 255154 543978 255774 544046
rect 255154 543922 255250 543978
rect 255306 543922 255374 543978
rect 255430 543922 255498 543978
rect 255554 543922 255622 543978
rect 255678 543922 255774 543978
rect 255154 526350 255774 543922
rect 255154 526294 255250 526350
rect 255306 526294 255374 526350
rect 255430 526294 255498 526350
rect 255554 526294 255622 526350
rect 255678 526294 255774 526350
rect 255154 526226 255774 526294
rect 255154 526170 255250 526226
rect 255306 526170 255374 526226
rect 255430 526170 255498 526226
rect 255554 526170 255622 526226
rect 255678 526170 255774 526226
rect 255154 526102 255774 526170
rect 255154 526046 255250 526102
rect 255306 526046 255374 526102
rect 255430 526046 255498 526102
rect 255554 526046 255622 526102
rect 255678 526046 255774 526102
rect 255154 525978 255774 526046
rect 255154 525922 255250 525978
rect 255306 525922 255374 525978
rect 255430 525922 255498 525978
rect 255554 525922 255622 525978
rect 255678 525922 255774 525978
rect 255154 508350 255774 525922
rect 255154 508294 255250 508350
rect 255306 508294 255374 508350
rect 255430 508294 255498 508350
rect 255554 508294 255622 508350
rect 255678 508294 255774 508350
rect 255154 508226 255774 508294
rect 255154 508170 255250 508226
rect 255306 508170 255374 508226
rect 255430 508170 255498 508226
rect 255554 508170 255622 508226
rect 255678 508170 255774 508226
rect 255154 508102 255774 508170
rect 255154 508046 255250 508102
rect 255306 508046 255374 508102
rect 255430 508046 255498 508102
rect 255554 508046 255622 508102
rect 255678 508046 255774 508102
rect 255154 507978 255774 508046
rect 255154 507922 255250 507978
rect 255306 507922 255374 507978
rect 255430 507922 255498 507978
rect 255554 507922 255622 507978
rect 255678 507922 255774 507978
rect 255154 490350 255774 507922
rect 255154 490294 255250 490350
rect 255306 490294 255374 490350
rect 255430 490294 255498 490350
rect 255554 490294 255622 490350
rect 255678 490294 255774 490350
rect 255154 490226 255774 490294
rect 255154 490170 255250 490226
rect 255306 490170 255374 490226
rect 255430 490170 255498 490226
rect 255554 490170 255622 490226
rect 255678 490170 255774 490226
rect 255154 490102 255774 490170
rect 255154 490046 255250 490102
rect 255306 490046 255374 490102
rect 255430 490046 255498 490102
rect 255554 490046 255622 490102
rect 255678 490046 255774 490102
rect 255154 489978 255774 490046
rect 255154 489922 255250 489978
rect 255306 489922 255374 489978
rect 255430 489922 255498 489978
rect 255554 489922 255622 489978
rect 255678 489922 255774 489978
rect 255154 472350 255774 489922
rect 255154 472294 255250 472350
rect 255306 472294 255374 472350
rect 255430 472294 255498 472350
rect 255554 472294 255622 472350
rect 255678 472294 255774 472350
rect 255154 472226 255774 472294
rect 255154 472170 255250 472226
rect 255306 472170 255374 472226
rect 255430 472170 255498 472226
rect 255554 472170 255622 472226
rect 255678 472170 255774 472226
rect 255154 472102 255774 472170
rect 255154 472046 255250 472102
rect 255306 472046 255374 472102
rect 255430 472046 255498 472102
rect 255554 472046 255622 472102
rect 255678 472046 255774 472102
rect 255154 471978 255774 472046
rect 255154 471922 255250 471978
rect 255306 471922 255374 471978
rect 255430 471922 255498 471978
rect 255554 471922 255622 471978
rect 255678 471922 255774 471978
rect 255154 458342 255774 471922
rect 258874 598172 259494 598268
rect 258874 598116 258970 598172
rect 259026 598116 259094 598172
rect 259150 598116 259218 598172
rect 259274 598116 259342 598172
rect 259398 598116 259494 598172
rect 258874 598048 259494 598116
rect 258874 597992 258970 598048
rect 259026 597992 259094 598048
rect 259150 597992 259218 598048
rect 259274 597992 259342 598048
rect 259398 597992 259494 598048
rect 258874 597924 259494 597992
rect 258874 597868 258970 597924
rect 259026 597868 259094 597924
rect 259150 597868 259218 597924
rect 259274 597868 259342 597924
rect 259398 597868 259494 597924
rect 258874 597800 259494 597868
rect 258874 597744 258970 597800
rect 259026 597744 259094 597800
rect 259150 597744 259218 597800
rect 259274 597744 259342 597800
rect 259398 597744 259494 597800
rect 258874 586350 259494 597744
rect 258874 586294 258970 586350
rect 259026 586294 259094 586350
rect 259150 586294 259218 586350
rect 259274 586294 259342 586350
rect 259398 586294 259494 586350
rect 258874 586226 259494 586294
rect 258874 586170 258970 586226
rect 259026 586170 259094 586226
rect 259150 586170 259218 586226
rect 259274 586170 259342 586226
rect 259398 586170 259494 586226
rect 258874 586102 259494 586170
rect 258874 586046 258970 586102
rect 259026 586046 259094 586102
rect 259150 586046 259218 586102
rect 259274 586046 259342 586102
rect 259398 586046 259494 586102
rect 258874 585978 259494 586046
rect 258874 585922 258970 585978
rect 259026 585922 259094 585978
rect 259150 585922 259218 585978
rect 259274 585922 259342 585978
rect 259398 585922 259494 585978
rect 258874 568350 259494 585922
rect 258874 568294 258970 568350
rect 259026 568294 259094 568350
rect 259150 568294 259218 568350
rect 259274 568294 259342 568350
rect 259398 568294 259494 568350
rect 258874 568226 259494 568294
rect 258874 568170 258970 568226
rect 259026 568170 259094 568226
rect 259150 568170 259218 568226
rect 259274 568170 259342 568226
rect 259398 568170 259494 568226
rect 258874 568102 259494 568170
rect 258874 568046 258970 568102
rect 259026 568046 259094 568102
rect 259150 568046 259218 568102
rect 259274 568046 259342 568102
rect 259398 568046 259494 568102
rect 258874 567978 259494 568046
rect 258874 567922 258970 567978
rect 259026 567922 259094 567978
rect 259150 567922 259218 567978
rect 259274 567922 259342 567978
rect 259398 567922 259494 567978
rect 258874 550350 259494 567922
rect 258874 550294 258970 550350
rect 259026 550294 259094 550350
rect 259150 550294 259218 550350
rect 259274 550294 259342 550350
rect 259398 550294 259494 550350
rect 258874 550226 259494 550294
rect 258874 550170 258970 550226
rect 259026 550170 259094 550226
rect 259150 550170 259218 550226
rect 259274 550170 259342 550226
rect 259398 550170 259494 550226
rect 258874 550102 259494 550170
rect 258874 550046 258970 550102
rect 259026 550046 259094 550102
rect 259150 550046 259218 550102
rect 259274 550046 259342 550102
rect 259398 550046 259494 550102
rect 258874 549978 259494 550046
rect 258874 549922 258970 549978
rect 259026 549922 259094 549978
rect 259150 549922 259218 549978
rect 259274 549922 259342 549978
rect 259398 549922 259494 549978
rect 258874 532350 259494 549922
rect 258874 532294 258970 532350
rect 259026 532294 259094 532350
rect 259150 532294 259218 532350
rect 259274 532294 259342 532350
rect 259398 532294 259494 532350
rect 258874 532226 259494 532294
rect 258874 532170 258970 532226
rect 259026 532170 259094 532226
rect 259150 532170 259218 532226
rect 259274 532170 259342 532226
rect 259398 532170 259494 532226
rect 258874 532102 259494 532170
rect 258874 532046 258970 532102
rect 259026 532046 259094 532102
rect 259150 532046 259218 532102
rect 259274 532046 259342 532102
rect 259398 532046 259494 532102
rect 258874 531978 259494 532046
rect 258874 531922 258970 531978
rect 259026 531922 259094 531978
rect 259150 531922 259218 531978
rect 259274 531922 259342 531978
rect 259398 531922 259494 531978
rect 258874 514350 259494 531922
rect 258874 514294 258970 514350
rect 259026 514294 259094 514350
rect 259150 514294 259218 514350
rect 259274 514294 259342 514350
rect 259398 514294 259494 514350
rect 258874 514226 259494 514294
rect 258874 514170 258970 514226
rect 259026 514170 259094 514226
rect 259150 514170 259218 514226
rect 259274 514170 259342 514226
rect 259398 514170 259494 514226
rect 258874 514102 259494 514170
rect 258874 514046 258970 514102
rect 259026 514046 259094 514102
rect 259150 514046 259218 514102
rect 259274 514046 259342 514102
rect 259398 514046 259494 514102
rect 258874 513978 259494 514046
rect 258874 513922 258970 513978
rect 259026 513922 259094 513978
rect 259150 513922 259218 513978
rect 259274 513922 259342 513978
rect 259398 513922 259494 513978
rect 258874 496350 259494 513922
rect 258874 496294 258970 496350
rect 259026 496294 259094 496350
rect 259150 496294 259218 496350
rect 259274 496294 259342 496350
rect 259398 496294 259494 496350
rect 258874 496226 259494 496294
rect 258874 496170 258970 496226
rect 259026 496170 259094 496226
rect 259150 496170 259218 496226
rect 259274 496170 259342 496226
rect 259398 496170 259494 496226
rect 258874 496102 259494 496170
rect 258874 496046 258970 496102
rect 259026 496046 259094 496102
rect 259150 496046 259218 496102
rect 259274 496046 259342 496102
rect 259398 496046 259494 496102
rect 258874 495978 259494 496046
rect 258874 495922 258970 495978
rect 259026 495922 259094 495978
rect 259150 495922 259218 495978
rect 259274 495922 259342 495978
rect 259398 495922 259494 495978
rect 258874 478350 259494 495922
rect 258874 478294 258970 478350
rect 259026 478294 259094 478350
rect 259150 478294 259218 478350
rect 259274 478294 259342 478350
rect 259398 478294 259494 478350
rect 258874 478226 259494 478294
rect 258874 478170 258970 478226
rect 259026 478170 259094 478226
rect 259150 478170 259218 478226
rect 259274 478170 259342 478226
rect 259398 478170 259494 478226
rect 258874 478102 259494 478170
rect 258874 478046 258970 478102
rect 259026 478046 259094 478102
rect 259150 478046 259218 478102
rect 259274 478046 259342 478102
rect 259398 478046 259494 478102
rect 258874 477978 259494 478046
rect 258874 477922 258970 477978
rect 259026 477922 259094 477978
rect 259150 477922 259218 477978
rect 259274 477922 259342 477978
rect 259398 477922 259494 477978
rect 258874 460350 259494 477922
rect 258874 460294 258970 460350
rect 259026 460294 259094 460350
rect 259150 460294 259218 460350
rect 259274 460294 259342 460350
rect 259398 460294 259494 460350
rect 258874 460226 259494 460294
rect 258874 460170 258970 460226
rect 259026 460170 259094 460226
rect 259150 460170 259218 460226
rect 259274 460170 259342 460226
rect 259398 460170 259494 460226
rect 258874 460102 259494 460170
rect 258874 460046 258970 460102
rect 259026 460046 259094 460102
rect 259150 460046 259218 460102
rect 259274 460046 259342 460102
rect 259398 460046 259494 460102
rect 258874 459978 259494 460046
rect 258874 459922 258970 459978
rect 259026 459922 259094 459978
rect 259150 459922 259218 459978
rect 259274 459922 259342 459978
rect 259398 459922 259494 459978
rect 258874 458342 259494 459922
rect 273154 597212 273774 598268
rect 273154 597156 273250 597212
rect 273306 597156 273374 597212
rect 273430 597156 273498 597212
rect 273554 597156 273622 597212
rect 273678 597156 273774 597212
rect 273154 597088 273774 597156
rect 273154 597032 273250 597088
rect 273306 597032 273374 597088
rect 273430 597032 273498 597088
rect 273554 597032 273622 597088
rect 273678 597032 273774 597088
rect 273154 596964 273774 597032
rect 273154 596908 273250 596964
rect 273306 596908 273374 596964
rect 273430 596908 273498 596964
rect 273554 596908 273622 596964
rect 273678 596908 273774 596964
rect 273154 596840 273774 596908
rect 273154 596784 273250 596840
rect 273306 596784 273374 596840
rect 273430 596784 273498 596840
rect 273554 596784 273622 596840
rect 273678 596784 273774 596840
rect 273154 580350 273774 596784
rect 273154 580294 273250 580350
rect 273306 580294 273374 580350
rect 273430 580294 273498 580350
rect 273554 580294 273622 580350
rect 273678 580294 273774 580350
rect 273154 580226 273774 580294
rect 273154 580170 273250 580226
rect 273306 580170 273374 580226
rect 273430 580170 273498 580226
rect 273554 580170 273622 580226
rect 273678 580170 273774 580226
rect 273154 580102 273774 580170
rect 273154 580046 273250 580102
rect 273306 580046 273374 580102
rect 273430 580046 273498 580102
rect 273554 580046 273622 580102
rect 273678 580046 273774 580102
rect 273154 579978 273774 580046
rect 273154 579922 273250 579978
rect 273306 579922 273374 579978
rect 273430 579922 273498 579978
rect 273554 579922 273622 579978
rect 273678 579922 273774 579978
rect 273154 562350 273774 579922
rect 273154 562294 273250 562350
rect 273306 562294 273374 562350
rect 273430 562294 273498 562350
rect 273554 562294 273622 562350
rect 273678 562294 273774 562350
rect 273154 562226 273774 562294
rect 273154 562170 273250 562226
rect 273306 562170 273374 562226
rect 273430 562170 273498 562226
rect 273554 562170 273622 562226
rect 273678 562170 273774 562226
rect 273154 562102 273774 562170
rect 273154 562046 273250 562102
rect 273306 562046 273374 562102
rect 273430 562046 273498 562102
rect 273554 562046 273622 562102
rect 273678 562046 273774 562102
rect 273154 561978 273774 562046
rect 273154 561922 273250 561978
rect 273306 561922 273374 561978
rect 273430 561922 273498 561978
rect 273554 561922 273622 561978
rect 273678 561922 273774 561978
rect 273154 544350 273774 561922
rect 273154 544294 273250 544350
rect 273306 544294 273374 544350
rect 273430 544294 273498 544350
rect 273554 544294 273622 544350
rect 273678 544294 273774 544350
rect 273154 544226 273774 544294
rect 273154 544170 273250 544226
rect 273306 544170 273374 544226
rect 273430 544170 273498 544226
rect 273554 544170 273622 544226
rect 273678 544170 273774 544226
rect 273154 544102 273774 544170
rect 273154 544046 273250 544102
rect 273306 544046 273374 544102
rect 273430 544046 273498 544102
rect 273554 544046 273622 544102
rect 273678 544046 273774 544102
rect 273154 543978 273774 544046
rect 273154 543922 273250 543978
rect 273306 543922 273374 543978
rect 273430 543922 273498 543978
rect 273554 543922 273622 543978
rect 273678 543922 273774 543978
rect 273154 526350 273774 543922
rect 273154 526294 273250 526350
rect 273306 526294 273374 526350
rect 273430 526294 273498 526350
rect 273554 526294 273622 526350
rect 273678 526294 273774 526350
rect 273154 526226 273774 526294
rect 273154 526170 273250 526226
rect 273306 526170 273374 526226
rect 273430 526170 273498 526226
rect 273554 526170 273622 526226
rect 273678 526170 273774 526226
rect 273154 526102 273774 526170
rect 273154 526046 273250 526102
rect 273306 526046 273374 526102
rect 273430 526046 273498 526102
rect 273554 526046 273622 526102
rect 273678 526046 273774 526102
rect 273154 525978 273774 526046
rect 273154 525922 273250 525978
rect 273306 525922 273374 525978
rect 273430 525922 273498 525978
rect 273554 525922 273622 525978
rect 273678 525922 273774 525978
rect 273154 508350 273774 525922
rect 273154 508294 273250 508350
rect 273306 508294 273374 508350
rect 273430 508294 273498 508350
rect 273554 508294 273622 508350
rect 273678 508294 273774 508350
rect 273154 508226 273774 508294
rect 273154 508170 273250 508226
rect 273306 508170 273374 508226
rect 273430 508170 273498 508226
rect 273554 508170 273622 508226
rect 273678 508170 273774 508226
rect 273154 508102 273774 508170
rect 273154 508046 273250 508102
rect 273306 508046 273374 508102
rect 273430 508046 273498 508102
rect 273554 508046 273622 508102
rect 273678 508046 273774 508102
rect 273154 507978 273774 508046
rect 273154 507922 273250 507978
rect 273306 507922 273374 507978
rect 273430 507922 273498 507978
rect 273554 507922 273622 507978
rect 273678 507922 273774 507978
rect 273154 490350 273774 507922
rect 273154 490294 273250 490350
rect 273306 490294 273374 490350
rect 273430 490294 273498 490350
rect 273554 490294 273622 490350
rect 273678 490294 273774 490350
rect 273154 490226 273774 490294
rect 273154 490170 273250 490226
rect 273306 490170 273374 490226
rect 273430 490170 273498 490226
rect 273554 490170 273622 490226
rect 273678 490170 273774 490226
rect 273154 490102 273774 490170
rect 273154 490046 273250 490102
rect 273306 490046 273374 490102
rect 273430 490046 273498 490102
rect 273554 490046 273622 490102
rect 273678 490046 273774 490102
rect 273154 489978 273774 490046
rect 273154 489922 273250 489978
rect 273306 489922 273374 489978
rect 273430 489922 273498 489978
rect 273554 489922 273622 489978
rect 273678 489922 273774 489978
rect 273154 472350 273774 489922
rect 273154 472294 273250 472350
rect 273306 472294 273374 472350
rect 273430 472294 273498 472350
rect 273554 472294 273622 472350
rect 273678 472294 273774 472350
rect 273154 472226 273774 472294
rect 273154 472170 273250 472226
rect 273306 472170 273374 472226
rect 273430 472170 273498 472226
rect 273554 472170 273622 472226
rect 273678 472170 273774 472226
rect 273154 472102 273774 472170
rect 273154 472046 273250 472102
rect 273306 472046 273374 472102
rect 273430 472046 273498 472102
rect 273554 472046 273622 472102
rect 273678 472046 273774 472102
rect 273154 471978 273774 472046
rect 273154 471922 273250 471978
rect 273306 471922 273374 471978
rect 273430 471922 273498 471978
rect 273554 471922 273622 471978
rect 273678 471922 273774 471978
rect 273154 458342 273774 471922
rect 276874 598172 277494 598268
rect 276874 598116 276970 598172
rect 277026 598116 277094 598172
rect 277150 598116 277218 598172
rect 277274 598116 277342 598172
rect 277398 598116 277494 598172
rect 276874 598048 277494 598116
rect 276874 597992 276970 598048
rect 277026 597992 277094 598048
rect 277150 597992 277218 598048
rect 277274 597992 277342 598048
rect 277398 597992 277494 598048
rect 276874 597924 277494 597992
rect 276874 597868 276970 597924
rect 277026 597868 277094 597924
rect 277150 597868 277218 597924
rect 277274 597868 277342 597924
rect 277398 597868 277494 597924
rect 276874 597800 277494 597868
rect 276874 597744 276970 597800
rect 277026 597744 277094 597800
rect 277150 597744 277218 597800
rect 277274 597744 277342 597800
rect 277398 597744 277494 597800
rect 276874 586350 277494 597744
rect 276874 586294 276970 586350
rect 277026 586294 277094 586350
rect 277150 586294 277218 586350
rect 277274 586294 277342 586350
rect 277398 586294 277494 586350
rect 276874 586226 277494 586294
rect 276874 586170 276970 586226
rect 277026 586170 277094 586226
rect 277150 586170 277218 586226
rect 277274 586170 277342 586226
rect 277398 586170 277494 586226
rect 276874 586102 277494 586170
rect 276874 586046 276970 586102
rect 277026 586046 277094 586102
rect 277150 586046 277218 586102
rect 277274 586046 277342 586102
rect 277398 586046 277494 586102
rect 276874 585978 277494 586046
rect 276874 585922 276970 585978
rect 277026 585922 277094 585978
rect 277150 585922 277218 585978
rect 277274 585922 277342 585978
rect 277398 585922 277494 585978
rect 276874 568350 277494 585922
rect 276874 568294 276970 568350
rect 277026 568294 277094 568350
rect 277150 568294 277218 568350
rect 277274 568294 277342 568350
rect 277398 568294 277494 568350
rect 276874 568226 277494 568294
rect 276874 568170 276970 568226
rect 277026 568170 277094 568226
rect 277150 568170 277218 568226
rect 277274 568170 277342 568226
rect 277398 568170 277494 568226
rect 276874 568102 277494 568170
rect 276874 568046 276970 568102
rect 277026 568046 277094 568102
rect 277150 568046 277218 568102
rect 277274 568046 277342 568102
rect 277398 568046 277494 568102
rect 276874 567978 277494 568046
rect 276874 567922 276970 567978
rect 277026 567922 277094 567978
rect 277150 567922 277218 567978
rect 277274 567922 277342 567978
rect 277398 567922 277494 567978
rect 276874 550350 277494 567922
rect 276874 550294 276970 550350
rect 277026 550294 277094 550350
rect 277150 550294 277218 550350
rect 277274 550294 277342 550350
rect 277398 550294 277494 550350
rect 276874 550226 277494 550294
rect 276874 550170 276970 550226
rect 277026 550170 277094 550226
rect 277150 550170 277218 550226
rect 277274 550170 277342 550226
rect 277398 550170 277494 550226
rect 276874 550102 277494 550170
rect 276874 550046 276970 550102
rect 277026 550046 277094 550102
rect 277150 550046 277218 550102
rect 277274 550046 277342 550102
rect 277398 550046 277494 550102
rect 276874 549978 277494 550046
rect 276874 549922 276970 549978
rect 277026 549922 277094 549978
rect 277150 549922 277218 549978
rect 277274 549922 277342 549978
rect 277398 549922 277494 549978
rect 276874 532350 277494 549922
rect 276874 532294 276970 532350
rect 277026 532294 277094 532350
rect 277150 532294 277218 532350
rect 277274 532294 277342 532350
rect 277398 532294 277494 532350
rect 276874 532226 277494 532294
rect 276874 532170 276970 532226
rect 277026 532170 277094 532226
rect 277150 532170 277218 532226
rect 277274 532170 277342 532226
rect 277398 532170 277494 532226
rect 276874 532102 277494 532170
rect 276874 532046 276970 532102
rect 277026 532046 277094 532102
rect 277150 532046 277218 532102
rect 277274 532046 277342 532102
rect 277398 532046 277494 532102
rect 276874 531978 277494 532046
rect 276874 531922 276970 531978
rect 277026 531922 277094 531978
rect 277150 531922 277218 531978
rect 277274 531922 277342 531978
rect 277398 531922 277494 531978
rect 276874 514350 277494 531922
rect 276874 514294 276970 514350
rect 277026 514294 277094 514350
rect 277150 514294 277218 514350
rect 277274 514294 277342 514350
rect 277398 514294 277494 514350
rect 276874 514226 277494 514294
rect 276874 514170 276970 514226
rect 277026 514170 277094 514226
rect 277150 514170 277218 514226
rect 277274 514170 277342 514226
rect 277398 514170 277494 514226
rect 276874 514102 277494 514170
rect 276874 514046 276970 514102
rect 277026 514046 277094 514102
rect 277150 514046 277218 514102
rect 277274 514046 277342 514102
rect 277398 514046 277494 514102
rect 276874 513978 277494 514046
rect 276874 513922 276970 513978
rect 277026 513922 277094 513978
rect 277150 513922 277218 513978
rect 277274 513922 277342 513978
rect 277398 513922 277494 513978
rect 276874 496350 277494 513922
rect 276874 496294 276970 496350
rect 277026 496294 277094 496350
rect 277150 496294 277218 496350
rect 277274 496294 277342 496350
rect 277398 496294 277494 496350
rect 276874 496226 277494 496294
rect 276874 496170 276970 496226
rect 277026 496170 277094 496226
rect 277150 496170 277218 496226
rect 277274 496170 277342 496226
rect 277398 496170 277494 496226
rect 276874 496102 277494 496170
rect 276874 496046 276970 496102
rect 277026 496046 277094 496102
rect 277150 496046 277218 496102
rect 277274 496046 277342 496102
rect 277398 496046 277494 496102
rect 276874 495978 277494 496046
rect 276874 495922 276970 495978
rect 277026 495922 277094 495978
rect 277150 495922 277218 495978
rect 277274 495922 277342 495978
rect 277398 495922 277494 495978
rect 276874 478350 277494 495922
rect 276874 478294 276970 478350
rect 277026 478294 277094 478350
rect 277150 478294 277218 478350
rect 277274 478294 277342 478350
rect 277398 478294 277494 478350
rect 276874 478226 277494 478294
rect 276874 478170 276970 478226
rect 277026 478170 277094 478226
rect 277150 478170 277218 478226
rect 277274 478170 277342 478226
rect 277398 478170 277494 478226
rect 276874 478102 277494 478170
rect 276874 478046 276970 478102
rect 277026 478046 277094 478102
rect 277150 478046 277218 478102
rect 277274 478046 277342 478102
rect 277398 478046 277494 478102
rect 276874 477978 277494 478046
rect 276874 477922 276970 477978
rect 277026 477922 277094 477978
rect 277150 477922 277218 477978
rect 277274 477922 277342 477978
rect 277398 477922 277494 477978
rect 276874 460350 277494 477922
rect 276874 460294 276970 460350
rect 277026 460294 277094 460350
rect 277150 460294 277218 460350
rect 277274 460294 277342 460350
rect 277398 460294 277494 460350
rect 276874 460226 277494 460294
rect 276874 460170 276970 460226
rect 277026 460170 277094 460226
rect 277150 460170 277218 460226
rect 277274 460170 277342 460226
rect 277398 460170 277494 460226
rect 276874 460102 277494 460170
rect 276874 460046 276970 460102
rect 277026 460046 277094 460102
rect 277150 460046 277218 460102
rect 277274 460046 277342 460102
rect 277398 460046 277494 460102
rect 276874 459978 277494 460046
rect 276874 459922 276970 459978
rect 277026 459922 277094 459978
rect 277150 459922 277218 459978
rect 277274 459922 277342 459978
rect 277398 459922 277494 459978
rect 276874 458342 277494 459922
rect 291154 597212 291774 598268
rect 291154 597156 291250 597212
rect 291306 597156 291374 597212
rect 291430 597156 291498 597212
rect 291554 597156 291622 597212
rect 291678 597156 291774 597212
rect 291154 597088 291774 597156
rect 291154 597032 291250 597088
rect 291306 597032 291374 597088
rect 291430 597032 291498 597088
rect 291554 597032 291622 597088
rect 291678 597032 291774 597088
rect 291154 596964 291774 597032
rect 291154 596908 291250 596964
rect 291306 596908 291374 596964
rect 291430 596908 291498 596964
rect 291554 596908 291622 596964
rect 291678 596908 291774 596964
rect 291154 596840 291774 596908
rect 291154 596784 291250 596840
rect 291306 596784 291374 596840
rect 291430 596784 291498 596840
rect 291554 596784 291622 596840
rect 291678 596784 291774 596840
rect 291154 580350 291774 596784
rect 291154 580294 291250 580350
rect 291306 580294 291374 580350
rect 291430 580294 291498 580350
rect 291554 580294 291622 580350
rect 291678 580294 291774 580350
rect 291154 580226 291774 580294
rect 291154 580170 291250 580226
rect 291306 580170 291374 580226
rect 291430 580170 291498 580226
rect 291554 580170 291622 580226
rect 291678 580170 291774 580226
rect 291154 580102 291774 580170
rect 291154 580046 291250 580102
rect 291306 580046 291374 580102
rect 291430 580046 291498 580102
rect 291554 580046 291622 580102
rect 291678 580046 291774 580102
rect 291154 579978 291774 580046
rect 291154 579922 291250 579978
rect 291306 579922 291374 579978
rect 291430 579922 291498 579978
rect 291554 579922 291622 579978
rect 291678 579922 291774 579978
rect 291154 562350 291774 579922
rect 291154 562294 291250 562350
rect 291306 562294 291374 562350
rect 291430 562294 291498 562350
rect 291554 562294 291622 562350
rect 291678 562294 291774 562350
rect 291154 562226 291774 562294
rect 291154 562170 291250 562226
rect 291306 562170 291374 562226
rect 291430 562170 291498 562226
rect 291554 562170 291622 562226
rect 291678 562170 291774 562226
rect 291154 562102 291774 562170
rect 291154 562046 291250 562102
rect 291306 562046 291374 562102
rect 291430 562046 291498 562102
rect 291554 562046 291622 562102
rect 291678 562046 291774 562102
rect 291154 561978 291774 562046
rect 291154 561922 291250 561978
rect 291306 561922 291374 561978
rect 291430 561922 291498 561978
rect 291554 561922 291622 561978
rect 291678 561922 291774 561978
rect 291154 544350 291774 561922
rect 291154 544294 291250 544350
rect 291306 544294 291374 544350
rect 291430 544294 291498 544350
rect 291554 544294 291622 544350
rect 291678 544294 291774 544350
rect 291154 544226 291774 544294
rect 291154 544170 291250 544226
rect 291306 544170 291374 544226
rect 291430 544170 291498 544226
rect 291554 544170 291622 544226
rect 291678 544170 291774 544226
rect 291154 544102 291774 544170
rect 291154 544046 291250 544102
rect 291306 544046 291374 544102
rect 291430 544046 291498 544102
rect 291554 544046 291622 544102
rect 291678 544046 291774 544102
rect 291154 543978 291774 544046
rect 291154 543922 291250 543978
rect 291306 543922 291374 543978
rect 291430 543922 291498 543978
rect 291554 543922 291622 543978
rect 291678 543922 291774 543978
rect 291154 526350 291774 543922
rect 291154 526294 291250 526350
rect 291306 526294 291374 526350
rect 291430 526294 291498 526350
rect 291554 526294 291622 526350
rect 291678 526294 291774 526350
rect 291154 526226 291774 526294
rect 291154 526170 291250 526226
rect 291306 526170 291374 526226
rect 291430 526170 291498 526226
rect 291554 526170 291622 526226
rect 291678 526170 291774 526226
rect 291154 526102 291774 526170
rect 291154 526046 291250 526102
rect 291306 526046 291374 526102
rect 291430 526046 291498 526102
rect 291554 526046 291622 526102
rect 291678 526046 291774 526102
rect 291154 525978 291774 526046
rect 291154 525922 291250 525978
rect 291306 525922 291374 525978
rect 291430 525922 291498 525978
rect 291554 525922 291622 525978
rect 291678 525922 291774 525978
rect 291154 508350 291774 525922
rect 291154 508294 291250 508350
rect 291306 508294 291374 508350
rect 291430 508294 291498 508350
rect 291554 508294 291622 508350
rect 291678 508294 291774 508350
rect 291154 508226 291774 508294
rect 291154 508170 291250 508226
rect 291306 508170 291374 508226
rect 291430 508170 291498 508226
rect 291554 508170 291622 508226
rect 291678 508170 291774 508226
rect 291154 508102 291774 508170
rect 291154 508046 291250 508102
rect 291306 508046 291374 508102
rect 291430 508046 291498 508102
rect 291554 508046 291622 508102
rect 291678 508046 291774 508102
rect 291154 507978 291774 508046
rect 291154 507922 291250 507978
rect 291306 507922 291374 507978
rect 291430 507922 291498 507978
rect 291554 507922 291622 507978
rect 291678 507922 291774 507978
rect 291154 490350 291774 507922
rect 291154 490294 291250 490350
rect 291306 490294 291374 490350
rect 291430 490294 291498 490350
rect 291554 490294 291622 490350
rect 291678 490294 291774 490350
rect 291154 490226 291774 490294
rect 291154 490170 291250 490226
rect 291306 490170 291374 490226
rect 291430 490170 291498 490226
rect 291554 490170 291622 490226
rect 291678 490170 291774 490226
rect 291154 490102 291774 490170
rect 291154 490046 291250 490102
rect 291306 490046 291374 490102
rect 291430 490046 291498 490102
rect 291554 490046 291622 490102
rect 291678 490046 291774 490102
rect 291154 489978 291774 490046
rect 291154 489922 291250 489978
rect 291306 489922 291374 489978
rect 291430 489922 291498 489978
rect 291554 489922 291622 489978
rect 291678 489922 291774 489978
rect 291154 472350 291774 489922
rect 291154 472294 291250 472350
rect 291306 472294 291374 472350
rect 291430 472294 291498 472350
rect 291554 472294 291622 472350
rect 291678 472294 291774 472350
rect 291154 472226 291774 472294
rect 291154 472170 291250 472226
rect 291306 472170 291374 472226
rect 291430 472170 291498 472226
rect 291554 472170 291622 472226
rect 291678 472170 291774 472226
rect 291154 472102 291774 472170
rect 291154 472046 291250 472102
rect 291306 472046 291374 472102
rect 291430 472046 291498 472102
rect 291554 472046 291622 472102
rect 291678 472046 291774 472102
rect 291154 471978 291774 472046
rect 291154 471922 291250 471978
rect 291306 471922 291374 471978
rect 291430 471922 291498 471978
rect 291554 471922 291622 471978
rect 291678 471922 291774 471978
rect 291154 458342 291774 471922
rect 294874 598172 295494 598268
rect 294874 598116 294970 598172
rect 295026 598116 295094 598172
rect 295150 598116 295218 598172
rect 295274 598116 295342 598172
rect 295398 598116 295494 598172
rect 294874 598048 295494 598116
rect 294874 597992 294970 598048
rect 295026 597992 295094 598048
rect 295150 597992 295218 598048
rect 295274 597992 295342 598048
rect 295398 597992 295494 598048
rect 294874 597924 295494 597992
rect 294874 597868 294970 597924
rect 295026 597868 295094 597924
rect 295150 597868 295218 597924
rect 295274 597868 295342 597924
rect 295398 597868 295494 597924
rect 294874 597800 295494 597868
rect 294874 597744 294970 597800
rect 295026 597744 295094 597800
rect 295150 597744 295218 597800
rect 295274 597744 295342 597800
rect 295398 597744 295494 597800
rect 294874 586350 295494 597744
rect 294874 586294 294970 586350
rect 295026 586294 295094 586350
rect 295150 586294 295218 586350
rect 295274 586294 295342 586350
rect 295398 586294 295494 586350
rect 294874 586226 295494 586294
rect 294874 586170 294970 586226
rect 295026 586170 295094 586226
rect 295150 586170 295218 586226
rect 295274 586170 295342 586226
rect 295398 586170 295494 586226
rect 294874 586102 295494 586170
rect 294874 586046 294970 586102
rect 295026 586046 295094 586102
rect 295150 586046 295218 586102
rect 295274 586046 295342 586102
rect 295398 586046 295494 586102
rect 294874 585978 295494 586046
rect 294874 585922 294970 585978
rect 295026 585922 295094 585978
rect 295150 585922 295218 585978
rect 295274 585922 295342 585978
rect 295398 585922 295494 585978
rect 294874 568350 295494 585922
rect 294874 568294 294970 568350
rect 295026 568294 295094 568350
rect 295150 568294 295218 568350
rect 295274 568294 295342 568350
rect 295398 568294 295494 568350
rect 294874 568226 295494 568294
rect 294874 568170 294970 568226
rect 295026 568170 295094 568226
rect 295150 568170 295218 568226
rect 295274 568170 295342 568226
rect 295398 568170 295494 568226
rect 294874 568102 295494 568170
rect 294874 568046 294970 568102
rect 295026 568046 295094 568102
rect 295150 568046 295218 568102
rect 295274 568046 295342 568102
rect 295398 568046 295494 568102
rect 294874 567978 295494 568046
rect 294874 567922 294970 567978
rect 295026 567922 295094 567978
rect 295150 567922 295218 567978
rect 295274 567922 295342 567978
rect 295398 567922 295494 567978
rect 294874 550350 295494 567922
rect 294874 550294 294970 550350
rect 295026 550294 295094 550350
rect 295150 550294 295218 550350
rect 295274 550294 295342 550350
rect 295398 550294 295494 550350
rect 294874 550226 295494 550294
rect 294874 550170 294970 550226
rect 295026 550170 295094 550226
rect 295150 550170 295218 550226
rect 295274 550170 295342 550226
rect 295398 550170 295494 550226
rect 294874 550102 295494 550170
rect 294874 550046 294970 550102
rect 295026 550046 295094 550102
rect 295150 550046 295218 550102
rect 295274 550046 295342 550102
rect 295398 550046 295494 550102
rect 294874 549978 295494 550046
rect 294874 549922 294970 549978
rect 295026 549922 295094 549978
rect 295150 549922 295218 549978
rect 295274 549922 295342 549978
rect 295398 549922 295494 549978
rect 294874 532350 295494 549922
rect 294874 532294 294970 532350
rect 295026 532294 295094 532350
rect 295150 532294 295218 532350
rect 295274 532294 295342 532350
rect 295398 532294 295494 532350
rect 294874 532226 295494 532294
rect 294874 532170 294970 532226
rect 295026 532170 295094 532226
rect 295150 532170 295218 532226
rect 295274 532170 295342 532226
rect 295398 532170 295494 532226
rect 294874 532102 295494 532170
rect 294874 532046 294970 532102
rect 295026 532046 295094 532102
rect 295150 532046 295218 532102
rect 295274 532046 295342 532102
rect 295398 532046 295494 532102
rect 294874 531978 295494 532046
rect 294874 531922 294970 531978
rect 295026 531922 295094 531978
rect 295150 531922 295218 531978
rect 295274 531922 295342 531978
rect 295398 531922 295494 531978
rect 294874 514350 295494 531922
rect 294874 514294 294970 514350
rect 295026 514294 295094 514350
rect 295150 514294 295218 514350
rect 295274 514294 295342 514350
rect 295398 514294 295494 514350
rect 294874 514226 295494 514294
rect 294874 514170 294970 514226
rect 295026 514170 295094 514226
rect 295150 514170 295218 514226
rect 295274 514170 295342 514226
rect 295398 514170 295494 514226
rect 294874 514102 295494 514170
rect 294874 514046 294970 514102
rect 295026 514046 295094 514102
rect 295150 514046 295218 514102
rect 295274 514046 295342 514102
rect 295398 514046 295494 514102
rect 294874 513978 295494 514046
rect 294874 513922 294970 513978
rect 295026 513922 295094 513978
rect 295150 513922 295218 513978
rect 295274 513922 295342 513978
rect 295398 513922 295494 513978
rect 294874 496350 295494 513922
rect 294874 496294 294970 496350
rect 295026 496294 295094 496350
rect 295150 496294 295218 496350
rect 295274 496294 295342 496350
rect 295398 496294 295494 496350
rect 294874 496226 295494 496294
rect 294874 496170 294970 496226
rect 295026 496170 295094 496226
rect 295150 496170 295218 496226
rect 295274 496170 295342 496226
rect 295398 496170 295494 496226
rect 294874 496102 295494 496170
rect 294874 496046 294970 496102
rect 295026 496046 295094 496102
rect 295150 496046 295218 496102
rect 295274 496046 295342 496102
rect 295398 496046 295494 496102
rect 294874 495978 295494 496046
rect 294874 495922 294970 495978
rect 295026 495922 295094 495978
rect 295150 495922 295218 495978
rect 295274 495922 295342 495978
rect 295398 495922 295494 495978
rect 294874 478350 295494 495922
rect 294874 478294 294970 478350
rect 295026 478294 295094 478350
rect 295150 478294 295218 478350
rect 295274 478294 295342 478350
rect 295398 478294 295494 478350
rect 294874 478226 295494 478294
rect 294874 478170 294970 478226
rect 295026 478170 295094 478226
rect 295150 478170 295218 478226
rect 295274 478170 295342 478226
rect 295398 478170 295494 478226
rect 294874 478102 295494 478170
rect 294874 478046 294970 478102
rect 295026 478046 295094 478102
rect 295150 478046 295218 478102
rect 295274 478046 295342 478102
rect 295398 478046 295494 478102
rect 294874 477978 295494 478046
rect 294874 477922 294970 477978
rect 295026 477922 295094 477978
rect 295150 477922 295218 477978
rect 295274 477922 295342 477978
rect 295398 477922 295494 477978
rect 294874 460350 295494 477922
rect 294874 460294 294970 460350
rect 295026 460294 295094 460350
rect 295150 460294 295218 460350
rect 295274 460294 295342 460350
rect 295398 460294 295494 460350
rect 294874 460226 295494 460294
rect 294874 460170 294970 460226
rect 295026 460170 295094 460226
rect 295150 460170 295218 460226
rect 295274 460170 295342 460226
rect 295398 460170 295494 460226
rect 294874 460102 295494 460170
rect 294874 460046 294970 460102
rect 295026 460046 295094 460102
rect 295150 460046 295218 460102
rect 295274 460046 295342 460102
rect 295398 460046 295494 460102
rect 294874 459978 295494 460046
rect 294874 459922 294970 459978
rect 295026 459922 295094 459978
rect 295150 459922 295218 459978
rect 295274 459922 295342 459978
rect 295398 459922 295494 459978
rect 294874 458342 295494 459922
rect 309154 597212 309774 598268
rect 309154 597156 309250 597212
rect 309306 597156 309374 597212
rect 309430 597156 309498 597212
rect 309554 597156 309622 597212
rect 309678 597156 309774 597212
rect 309154 597088 309774 597156
rect 309154 597032 309250 597088
rect 309306 597032 309374 597088
rect 309430 597032 309498 597088
rect 309554 597032 309622 597088
rect 309678 597032 309774 597088
rect 309154 596964 309774 597032
rect 309154 596908 309250 596964
rect 309306 596908 309374 596964
rect 309430 596908 309498 596964
rect 309554 596908 309622 596964
rect 309678 596908 309774 596964
rect 309154 596840 309774 596908
rect 309154 596784 309250 596840
rect 309306 596784 309374 596840
rect 309430 596784 309498 596840
rect 309554 596784 309622 596840
rect 309678 596784 309774 596840
rect 309154 580350 309774 596784
rect 309154 580294 309250 580350
rect 309306 580294 309374 580350
rect 309430 580294 309498 580350
rect 309554 580294 309622 580350
rect 309678 580294 309774 580350
rect 309154 580226 309774 580294
rect 309154 580170 309250 580226
rect 309306 580170 309374 580226
rect 309430 580170 309498 580226
rect 309554 580170 309622 580226
rect 309678 580170 309774 580226
rect 309154 580102 309774 580170
rect 309154 580046 309250 580102
rect 309306 580046 309374 580102
rect 309430 580046 309498 580102
rect 309554 580046 309622 580102
rect 309678 580046 309774 580102
rect 309154 579978 309774 580046
rect 309154 579922 309250 579978
rect 309306 579922 309374 579978
rect 309430 579922 309498 579978
rect 309554 579922 309622 579978
rect 309678 579922 309774 579978
rect 309154 562350 309774 579922
rect 309154 562294 309250 562350
rect 309306 562294 309374 562350
rect 309430 562294 309498 562350
rect 309554 562294 309622 562350
rect 309678 562294 309774 562350
rect 309154 562226 309774 562294
rect 309154 562170 309250 562226
rect 309306 562170 309374 562226
rect 309430 562170 309498 562226
rect 309554 562170 309622 562226
rect 309678 562170 309774 562226
rect 309154 562102 309774 562170
rect 309154 562046 309250 562102
rect 309306 562046 309374 562102
rect 309430 562046 309498 562102
rect 309554 562046 309622 562102
rect 309678 562046 309774 562102
rect 309154 561978 309774 562046
rect 309154 561922 309250 561978
rect 309306 561922 309374 561978
rect 309430 561922 309498 561978
rect 309554 561922 309622 561978
rect 309678 561922 309774 561978
rect 309154 544350 309774 561922
rect 309154 544294 309250 544350
rect 309306 544294 309374 544350
rect 309430 544294 309498 544350
rect 309554 544294 309622 544350
rect 309678 544294 309774 544350
rect 309154 544226 309774 544294
rect 309154 544170 309250 544226
rect 309306 544170 309374 544226
rect 309430 544170 309498 544226
rect 309554 544170 309622 544226
rect 309678 544170 309774 544226
rect 309154 544102 309774 544170
rect 309154 544046 309250 544102
rect 309306 544046 309374 544102
rect 309430 544046 309498 544102
rect 309554 544046 309622 544102
rect 309678 544046 309774 544102
rect 309154 543978 309774 544046
rect 309154 543922 309250 543978
rect 309306 543922 309374 543978
rect 309430 543922 309498 543978
rect 309554 543922 309622 543978
rect 309678 543922 309774 543978
rect 309154 526350 309774 543922
rect 309154 526294 309250 526350
rect 309306 526294 309374 526350
rect 309430 526294 309498 526350
rect 309554 526294 309622 526350
rect 309678 526294 309774 526350
rect 309154 526226 309774 526294
rect 309154 526170 309250 526226
rect 309306 526170 309374 526226
rect 309430 526170 309498 526226
rect 309554 526170 309622 526226
rect 309678 526170 309774 526226
rect 309154 526102 309774 526170
rect 309154 526046 309250 526102
rect 309306 526046 309374 526102
rect 309430 526046 309498 526102
rect 309554 526046 309622 526102
rect 309678 526046 309774 526102
rect 309154 525978 309774 526046
rect 309154 525922 309250 525978
rect 309306 525922 309374 525978
rect 309430 525922 309498 525978
rect 309554 525922 309622 525978
rect 309678 525922 309774 525978
rect 309154 508350 309774 525922
rect 309154 508294 309250 508350
rect 309306 508294 309374 508350
rect 309430 508294 309498 508350
rect 309554 508294 309622 508350
rect 309678 508294 309774 508350
rect 309154 508226 309774 508294
rect 309154 508170 309250 508226
rect 309306 508170 309374 508226
rect 309430 508170 309498 508226
rect 309554 508170 309622 508226
rect 309678 508170 309774 508226
rect 309154 508102 309774 508170
rect 309154 508046 309250 508102
rect 309306 508046 309374 508102
rect 309430 508046 309498 508102
rect 309554 508046 309622 508102
rect 309678 508046 309774 508102
rect 309154 507978 309774 508046
rect 309154 507922 309250 507978
rect 309306 507922 309374 507978
rect 309430 507922 309498 507978
rect 309554 507922 309622 507978
rect 309678 507922 309774 507978
rect 309154 490350 309774 507922
rect 309154 490294 309250 490350
rect 309306 490294 309374 490350
rect 309430 490294 309498 490350
rect 309554 490294 309622 490350
rect 309678 490294 309774 490350
rect 309154 490226 309774 490294
rect 309154 490170 309250 490226
rect 309306 490170 309374 490226
rect 309430 490170 309498 490226
rect 309554 490170 309622 490226
rect 309678 490170 309774 490226
rect 309154 490102 309774 490170
rect 309154 490046 309250 490102
rect 309306 490046 309374 490102
rect 309430 490046 309498 490102
rect 309554 490046 309622 490102
rect 309678 490046 309774 490102
rect 309154 489978 309774 490046
rect 309154 489922 309250 489978
rect 309306 489922 309374 489978
rect 309430 489922 309498 489978
rect 309554 489922 309622 489978
rect 309678 489922 309774 489978
rect 309154 472350 309774 489922
rect 309154 472294 309250 472350
rect 309306 472294 309374 472350
rect 309430 472294 309498 472350
rect 309554 472294 309622 472350
rect 309678 472294 309774 472350
rect 309154 472226 309774 472294
rect 309154 472170 309250 472226
rect 309306 472170 309374 472226
rect 309430 472170 309498 472226
rect 309554 472170 309622 472226
rect 309678 472170 309774 472226
rect 309154 472102 309774 472170
rect 309154 472046 309250 472102
rect 309306 472046 309374 472102
rect 309430 472046 309498 472102
rect 309554 472046 309622 472102
rect 309678 472046 309774 472102
rect 309154 471978 309774 472046
rect 309154 471922 309250 471978
rect 309306 471922 309374 471978
rect 309430 471922 309498 471978
rect 309554 471922 309622 471978
rect 309678 471922 309774 471978
rect 309154 458342 309774 471922
rect 312874 598172 313494 598268
rect 312874 598116 312970 598172
rect 313026 598116 313094 598172
rect 313150 598116 313218 598172
rect 313274 598116 313342 598172
rect 313398 598116 313494 598172
rect 312874 598048 313494 598116
rect 312874 597992 312970 598048
rect 313026 597992 313094 598048
rect 313150 597992 313218 598048
rect 313274 597992 313342 598048
rect 313398 597992 313494 598048
rect 312874 597924 313494 597992
rect 312874 597868 312970 597924
rect 313026 597868 313094 597924
rect 313150 597868 313218 597924
rect 313274 597868 313342 597924
rect 313398 597868 313494 597924
rect 312874 597800 313494 597868
rect 312874 597744 312970 597800
rect 313026 597744 313094 597800
rect 313150 597744 313218 597800
rect 313274 597744 313342 597800
rect 313398 597744 313494 597800
rect 312874 586350 313494 597744
rect 312874 586294 312970 586350
rect 313026 586294 313094 586350
rect 313150 586294 313218 586350
rect 313274 586294 313342 586350
rect 313398 586294 313494 586350
rect 312874 586226 313494 586294
rect 312874 586170 312970 586226
rect 313026 586170 313094 586226
rect 313150 586170 313218 586226
rect 313274 586170 313342 586226
rect 313398 586170 313494 586226
rect 312874 586102 313494 586170
rect 312874 586046 312970 586102
rect 313026 586046 313094 586102
rect 313150 586046 313218 586102
rect 313274 586046 313342 586102
rect 313398 586046 313494 586102
rect 312874 585978 313494 586046
rect 312874 585922 312970 585978
rect 313026 585922 313094 585978
rect 313150 585922 313218 585978
rect 313274 585922 313342 585978
rect 313398 585922 313494 585978
rect 312874 568350 313494 585922
rect 312874 568294 312970 568350
rect 313026 568294 313094 568350
rect 313150 568294 313218 568350
rect 313274 568294 313342 568350
rect 313398 568294 313494 568350
rect 312874 568226 313494 568294
rect 312874 568170 312970 568226
rect 313026 568170 313094 568226
rect 313150 568170 313218 568226
rect 313274 568170 313342 568226
rect 313398 568170 313494 568226
rect 312874 568102 313494 568170
rect 312874 568046 312970 568102
rect 313026 568046 313094 568102
rect 313150 568046 313218 568102
rect 313274 568046 313342 568102
rect 313398 568046 313494 568102
rect 312874 567978 313494 568046
rect 312874 567922 312970 567978
rect 313026 567922 313094 567978
rect 313150 567922 313218 567978
rect 313274 567922 313342 567978
rect 313398 567922 313494 567978
rect 312874 550350 313494 567922
rect 312874 550294 312970 550350
rect 313026 550294 313094 550350
rect 313150 550294 313218 550350
rect 313274 550294 313342 550350
rect 313398 550294 313494 550350
rect 312874 550226 313494 550294
rect 312874 550170 312970 550226
rect 313026 550170 313094 550226
rect 313150 550170 313218 550226
rect 313274 550170 313342 550226
rect 313398 550170 313494 550226
rect 312874 550102 313494 550170
rect 312874 550046 312970 550102
rect 313026 550046 313094 550102
rect 313150 550046 313218 550102
rect 313274 550046 313342 550102
rect 313398 550046 313494 550102
rect 312874 549978 313494 550046
rect 312874 549922 312970 549978
rect 313026 549922 313094 549978
rect 313150 549922 313218 549978
rect 313274 549922 313342 549978
rect 313398 549922 313494 549978
rect 312874 532350 313494 549922
rect 312874 532294 312970 532350
rect 313026 532294 313094 532350
rect 313150 532294 313218 532350
rect 313274 532294 313342 532350
rect 313398 532294 313494 532350
rect 312874 532226 313494 532294
rect 312874 532170 312970 532226
rect 313026 532170 313094 532226
rect 313150 532170 313218 532226
rect 313274 532170 313342 532226
rect 313398 532170 313494 532226
rect 312874 532102 313494 532170
rect 312874 532046 312970 532102
rect 313026 532046 313094 532102
rect 313150 532046 313218 532102
rect 313274 532046 313342 532102
rect 313398 532046 313494 532102
rect 312874 531978 313494 532046
rect 312874 531922 312970 531978
rect 313026 531922 313094 531978
rect 313150 531922 313218 531978
rect 313274 531922 313342 531978
rect 313398 531922 313494 531978
rect 312874 514350 313494 531922
rect 312874 514294 312970 514350
rect 313026 514294 313094 514350
rect 313150 514294 313218 514350
rect 313274 514294 313342 514350
rect 313398 514294 313494 514350
rect 312874 514226 313494 514294
rect 312874 514170 312970 514226
rect 313026 514170 313094 514226
rect 313150 514170 313218 514226
rect 313274 514170 313342 514226
rect 313398 514170 313494 514226
rect 312874 514102 313494 514170
rect 312874 514046 312970 514102
rect 313026 514046 313094 514102
rect 313150 514046 313218 514102
rect 313274 514046 313342 514102
rect 313398 514046 313494 514102
rect 312874 513978 313494 514046
rect 312874 513922 312970 513978
rect 313026 513922 313094 513978
rect 313150 513922 313218 513978
rect 313274 513922 313342 513978
rect 313398 513922 313494 513978
rect 312874 496350 313494 513922
rect 312874 496294 312970 496350
rect 313026 496294 313094 496350
rect 313150 496294 313218 496350
rect 313274 496294 313342 496350
rect 313398 496294 313494 496350
rect 312874 496226 313494 496294
rect 312874 496170 312970 496226
rect 313026 496170 313094 496226
rect 313150 496170 313218 496226
rect 313274 496170 313342 496226
rect 313398 496170 313494 496226
rect 312874 496102 313494 496170
rect 312874 496046 312970 496102
rect 313026 496046 313094 496102
rect 313150 496046 313218 496102
rect 313274 496046 313342 496102
rect 313398 496046 313494 496102
rect 312874 495978 313494 496046
rect 312874 495922 312970 495978
rect 313026 495922 313094 495978
rect 313150 495922 313218 495978
rect 313274 495922 313342 495978
rect 313398 495922 313494 495978
rect 312874 478350 313494 495922
rect 312874 478294 312970 478350
rect 313026 478294 313094 478350
rect 313150 478294 313218 478350
rect 313274 478294 313342 478350
rect 313398 478294 313494 478350
rect 312874 478226 313494 478294
rect 312874 478170 312970 478226
rect 313026 478170 313094 478226
rect 313150 478170 313218 478226
rect 313274 478170 313342 478226
rect 313398 478170 313494 478226
rect 312874 478102 313494 478170
rect 312874 478046 312970 478102
rect 313026 478046 313094 478102
rect 313150 478046 313218 478102
rect 313274 478046 313342 478102
rect 313398 478046 313494 478102
rect 312874 477978 313494 478046
rect 312874 477922 312970 477978
rect 313026 477922 313094 477978
rect 313150 477922 313218 477978
rect 313274 477922 313342 477978
rect 313398 477922 313494 477978
rect 312874 460350 313494 477922
rect 312874 460294 312970 460350
rect 313026 460294 313094 460350
rect 313150 460294 313218 460350
rect 313274 460294 313342 460350
rect 313398 460294 313494 460350
rect 312874 460226 313494 460294
rect 312874 460170 312970 460226
rect 313026 460170 313094 460226
rect 313150 460170 313218 460226
rect 313274 460170 313342 460226
rect 313398 460170 313494 460226
rect 312874 460102 313494 460170
rect 312874 460046 312970 460102
rect 313026 460046 313094 460102
rect 313150 460046 313218 460102
rect 313274 460046 313342 460102
rect 313398 460046 313494 460102
rect 312874 459978 313494 460046
rect 312874 459922 312970 459978
rect 313026 459922 313094 459978
rect 313150 459922 313218 459978
rect 313274 459922 313342 459978
rect 313398 459922 313494 459978
rect 312874 458342 313494 459922
rect 327154 597212 327774 598268
rect 327154 597156 327250 597212
rect 327306 597156 327374 597212
rect 327430 597156 327498 597212
rect 327554 597156 327622 597212
rect 327678 597156 327774 597212
rect 327154 597088 327774 597156
rect 327154 597032 327250 597088
rect 327306 597032 327374 597088
rect 327430 597032 327498 597088
rect 327554 597032 327622 597088
rect 327678 597032 327774 597088
rect 327154 596964 327774 597032
rect 327154 596908 327250 596964
rect 327306 596908 327374 596964
rect 327430 596908 327498 596964
rect 327554 596908 327622 596964
rect 327678 596908 327774 596964
rect 327154 596840 327774 596908
rect 327154 596784 327250 596840
rect 327306 596784 327374 596840
rect 327430 596784 327498 596840
rect 327554 596784 327622 596840
rect 327678 596784 327774 596840
rect 327154 580350 327774 596784
rect 327154 580294 327250 580350
rect 327306 580294 327374 580350
rect 327430 580294 327498 580350
rect 327554 580294 327622 580350
rect 327678 580294 327774 580350
rect 327154 580226 327774 580294
rect 327154 580170 327250 580226
rect 327306 580170 327374 580226
rect 327430 580170 327498 580226
rect 327554 580170 327622 580226
rect 327678 580170 327774 580226
rect 327154 580102 327774 580170
rect 327154 580046 327250 580102
rect 327306 580046 327374 580102
rect 327430 580046 327498 580102
rect 327554 580046 327622 580102
rect 327678 580046 327774 580102
rect 327154 579978 327774 580046
rect 327154 579922 327250 579978
rect 327306 579922 327374 579978
rect 327430 579922 327498 579978
rect 327554 579922 327622 579978
rect 327678 579922 327774 579978
rect 327154 562350 327774 579922
rect 327154 562294 327250 562350
rect 327306 562294 327374 562350
rect 327430 562294 327498 562350
rect 327554 562294 327622 562350
rect 327678 562294 327774 562350
rect 327154 562226 327774 562294
rect 327154 562170 327250 562226
rect 327306 562170 327374 562226
rect 327430 562170 327498 562226
rect 327554 562170 327622 562226
rect 327678 562170 327774 562226
rect 327154 562102 327774 562170
rect 327154 562046 327250 562102
rect 327306 562046 327374 562102
rect 327430 562046 327498 562102
rect 327554 562046 327622 562102
rect 327678 562046 327774 562102
rect 327154 561978 327774 562046
rect 327154 561922 327250 561978
rect 327306 561922 327374 561978
rect 327430 561922 327498 561978
rect 327554 561922 327622 561978
rect 327678 561922 327774 561978
rect 327154 544350 327774 561922
rect 327154 544294 327250 544350
rect 327306 544294 327374 544350
rect 327430 544294 327498 544350
rect 327554 544294 327622 544350
rect 327678 544294 327774 544350
rect 327154 544226 327774 544294
rect 327154 544170 327250 544226
rect 327306 544170 327374 544226
rect 327430 544170 327498 544226
rect 327554 544170 327622 544226
rect 327678 544170 327774 544226
rect 327154 544102 327774 544170
rect 327154 544046 327250 544102
rect 327306 544046 327374 544102
rect 327430 544046 327498 544102
rect 327554 544046 327622 544102
rect 327678 544046 327774 544102
rect 327154 543978 327774 544046
rect 327154 543922 327250 543978
rect 327306 543922 327374 543978
rect 327430 543922 327498 543978
rect 327554 543922 327622 543978
rect 327678 543922 327774 543978
rect 327154 526350 327774 543922
rect 327154 526294 327250 526350
rect 327306 526294 327374 526350
rect 327430 526294 327498 526350
rect 327554 526294 327622 526350
rect 327678 526294 327774 526350
rect 327154 526226 327774 526294
rect 327154 526170 327250 526226
rect 327306 526170 327374 526226
rect 327430 526170 327498 526226
rect 327554 526170 327622 526226
rect 327678 526170 327774 526226
rect 327154 526102 327774 526170
rect 327154 526046 327250 526102
rect 327306 526046 327374 526102
rect 327430 526046 327498 526102
rect 327554 526046 327622 526102
rect 327678 526046 327774 526102
rect 327154 525978 327774 526046
rect 327154 525922 327250 525978
rect 327306 525922 327374 525978
rect 327430 525922 327498 525978
rect 327554 525922 327622 525978
rect 327678 525922 327774 525978
rect 327154 508350 327774 525922
rect 327154 508294 327250 508350
rect 327306 508294 327374 508350
rect 327430 508294 327498 508350
rect 327554 508294 327622 508350
rect 327678 508294 327774 508350
rect 327154 508226 327774 508294
rect 327154 508170 327250 508226
rect 327306 508170 327374 508226
rect 327430 508170 327498 508226
rect 327554 508170 327622 508226
rect 327678 508170 327774 508226
rect 327154 508102 327774 508170
rect 327154 508046 327250 508102
rect 327306 508046 327374 508102
rect 327430 508046 327498 508102
rect 327554 508046 327622 508102
rect 327678 508046 327774 508102
rect 327154 507978 327774 508046
rect 327154 507922 327250 507978
rect 327306 507922 327374 507978
rect 327430 507922 327498 507978
rect 327554 507922 327622 507978
rect 327678 507922 327774 507978
rect 327154 490350 327774 507922
rect 327154 490294 327250 490350
rect 327306 490294 327374 490350
rect 327430 490294 327498 490350
rect 327554 490294 327622 490350
rect 327678 490294 327774 490350
rect 327154 490226 327774 490294
rect 327154 490170 327250 490226
rect 327306 490170 327374 490226
rect 327430 490170 327498 490226
rect 327554 490170 327622 490226
rect 327678 490170 327774 490226
rect 327154 490102 327774 490170
rect 327154 490046 327250 490102
rect 327306 490046 327374 490102
rect 327430 490046 327498 490102
rect 327554 490046 327622 490102
rect 327678 490046 327774 490102
rect 327154 489978 327774 490046
rect 327154 489922 327250 489978
rect 327306 489922 327374 489978
rect 327430 489922 327498 489978
rect 327554 489922 327622 489978
rect 327678 489922 327774 489978
rect 327154 472350 327774 489922
rect 327154 472294 327250 472350
rect 327306 472294 327374 472350
rect 327430 472294 327498 472350
rect 327554 472294 327622 472350
rect 327678 472294 327774 472350
rect 327154 472226 327774 472294
rect 327154 472170 327250 472226
rect 327306 472170 327374 472226
rect 327430 472170 327498 472226
rect 327554 472170 327622 472226
rect 327678 472170 327774 472226
rect 327154 472102 327774 472170
rect 327154 472046 327250 472102
rect 327306 472046 327374 472102
rect 327430 472046 327498 472102
rect 327554 472046 327622 472102
rect 327678 472046 327774 472102
rect 327154 471978 327774 472046
rect 327154 471922 327250 471978
rect 327306 471922 327374 471978
rect 327430 471922 327498 471978
rect 327554 471922 327622 471978
rect 327678 471922 327774 471978
rect 327154 458342 327774 471922
rect 330874 598172 331494 598268
rect 330874 598116 330970 598172
rect 331026 598116 331094 598172
rect 331150 598116 331218 598172
rect 331274 598116 331342 598172
rect 331398 598116 331494 598172
rect 330874 598048 331494 598116
rect 330874 597992 330970 598048
rect 331026 597992 331094 598048
rect 331150 597992 331218 598048
rect 331274 597992 331342 598048
rect 331398 597992 331494 598048
rect 330874 597924 331494 597992
rect 330874 597868 330970 597924
rect 331026 597868 331094 597924
rect 331150 597868 331218 597924
rect 331274 597868 331342 597924
rect 331398 597868 331494 597924
rect 330874 597800 331494 597868
rect 330874 597744 330970 597800
rect 331026 597744 331094 597800
rect 331150 597744 331218 597800
rect 331274 597744 331342 597800
rect 331398 597744 331494 597800
rect 330874 586350 331494 597744
rect 330874 586294 330970 586350
rect 331026 586294 331094 586350
rect 331150 586294 331218 586350
rect 331274 586294 331342 586350
rect 331398 586294 331494 586350
rect 330874 586226 331494 586294
rect 330874 586170 330970 586226
rect 331026 586170 331094 586226
rect 331150 586170 331218 586226
rect 331274 586170 331342 586226
rect 331398 586170 331494 586226
rect 330874 586102 331494 586170
rect 330874 586046 330970 586102
rect 331026 586046 331094 586102
rect 331150 586046 331218 586102
rect 331274 586046 331342 586102
rect 331398 586046 331494 586102
rect 330874 585978 331494 586046
rect 330874 585922 330970 585978
rect 331026 585922 331094 585978
rect 331150 585922 331218 585978
rect 331274 585922 331342 585978
rect 331398 585922 331494 585978
rect 330874 568350 331494 585922
rect 330874 568294 330970 568350
rect 331026 568294 331094 568350
rect 331150 568294 331218 568350
rect 331274 568294 331342 568350
rect 331398 568294 331494 568350
rect 330874 568226 331494 568294
rect 330874 568170 330970 568226
rect 331026 568170 331094 568226
rect 331150 568170 331218 568226
rect 331274 568170 331342 568226
rect 331398 568170 331494 568226
rect 330874 568102 331494 568170
rect 330874 568046 330970 568102
rect 331026 568046 331094 568102
rect 331150 568046 331218 568102
rect 331274 568046 331342 568102
rect 331398 568046 331494 568102
rect 330874 567978 331494 568046
rect 330874 567922 330970 567978
rect 331026 567922 331094 567978
rect 331150 567922 331218 567978
rect 331274 567922 331342 567978
rect 331398 567922 331494 567978
rect 330874 550350 331494 567922
rect 330874 550294 330970 550350
rect 331026 550294 331094 550350
rect 331150 550294 331218 550350
rect 331274 550294 331342 550350
rect 331398 550294 331494 550350
rect 330874 550226 331494 550294
rect 330874 550170 330970 550226
rect 331026 550170 331094 550226
rect 331150 550170 331218 550226
rect 331274 550170 331342 550226
rect 331398 550170 331494 550226
rect 330874 550102 331494 550170
rect 330874 550046 330970 550102
rect 331026 550046 331094 550102
rect 331150 550046 331218 550102
rect 331274 550046 331342 550102
rect 331398 550046 331494 550102
rect 330874 549978 331494 550046
rect 330874 549922 330970 549978
rect 331026 549922 331094 549978
rect 331150 549922 331218 549978
rect 331274 549922 331342 549978
rect 331398 549922 331494 549978
rect 330874 532350 331494 549922
rect 330874 532294 330970 532350
rect 331026 532294 331094 532350
rect 331150 532294 331218 532350
rect 331274 532294 331342 532350
rect 331398 532294 331494 532350
rect 330874 532226 331494 532294
rect 330874 532170 330970 532226
rect 331026 532170 331094 532226
rect 331150 532170 331218 532226
rect 331274 532170 331342 532226
rect 331398 532170 331494 532226
rect 330874 532102 331494 532170
rect 330874 532046 330970 532102
rect 331026 532046 331094 532102
rect 331150 532046 331218 532102
rect 331274 532046 331342 532102
rect 331398 532046 331494 532102
rect 330874 531978 331494 532046
rect 330874 531922 330970 531978
rect 331026 531922 331094 531978
rect 331150 531922 331218 531978
rect 331274 531922 331342 531978
rect 331398 531922 331494 531978
rect 330874 514350 331494 531922
rect 330874 514294 330970 514350
rect 331026 514294 331094 514350
rect 331150 514294 331218 514350
rect 331274 514294 331342 514350
rect 331398 514294 331494 514350
rect 330874 514226 331494 514294
rect 330874 514170 330970 514226
rect 331026 514170 331094 514226
rect 331150 514170 331218 514226
rect 331274 514170 331342 514226
rect 331398 514170 331494 514226
rect 330874 514102 331494 514170
rect 330874 514046 330970 514102
rect 331026 514046 331094 514102
rect 331150 514046 331218 514102
rect 331274 514046 331342 514102
rect 331398 514046 331494 514102
rect 330874 513978 331494 514046
rect 330874 513922 330970 513978
rect 331026 513922 331094 513978
rect 331150 513922 331218 513978
rect 331274 513922 331342 513978
rect 331398 513922 331494 513978
rect 330874 496350 331494 513922
rect 330874 496294 330970 496350
rect 331026 496294 331094 496350
rect 331150 496294 331218 496350
rect 331274 496294 331342 496350
rect 331398 496294 331494 496350
rect 330874 496226 331494 496294
rect 330874 496170 330970 496226
rect 331026 496170 331094 496226
rect 331150 496170 331218 496226
rect 331274 496170 331342 496226
rect 331398 496170 331494 496226
rect 330874 496102 331494 496170
rect 330874 496046 330970 496102
rect 331026 496046 331094 496102
rect 331150 496046 331218 496102
rect 331274 496046 331342 496102
rect 331398 496046 331494 496102
rect 330874 495978 331494 496046
rect 330874 495922 330970 495978
rect 331026 495922 331094 495978
rect 331150 495922 331218 495978
rect 331274 495922 331342 495978
rect 331398 495922 331494 495978
rect 330874 478350 331494 495922
rect 330874 478294 330970 478350
rect 331026 478294 331094 478350
rect 331150 478294 331218 478350
rect 331274 478294 331342 478350
rect 331398 478294 331494 478350
rect 330874 478226 331494 478294
rect 330874 478170 330970 478226
rect 331026 478170 331094 478226
rect 331150 478170 331218 478226
rect 331274 478170 331342 478226
rect 331398 478170 331494 478226
rect 330874 478102 331494 478170
rect 330874 478046 330970 478102
rect 331026 478046 331094 478102
rect 331150 478046 331218 478102
rect 331274 478046 331342 478102
rect 331398 478046 331494 478102
rect 330874 477978 331494 478046
rect 330874 477922 330970 477978
rect 331026 477922 331094 477978
rect 331150 477922 331218 477978
rect 331274 477922 331342 477978
rect 331398 477922 331494 477978
rect 330874 460350 331494 477922
rect 330874 460294 330970 460350
rect 331026 460294 331094 460350
rect 331150 460294 331218 460350
rect 331274 460294 331342 460350
rect 331398 460294 331494 460350
rect 330874 460226 331494 460294
rect 330874 460170 330970 460226
rect 331026 460170 331094 460226
rect 331150 460170 331218 460226
rect 331274 460170 331342 460226
rect 331398 460170 331494 460226
rect 330874 460102 331494 460170
rect 330874 460046 330970 460102
rect 331026 460046 331094 460102
rect 331150 460046 331218 460102
rect 331274 460046 331342 460102
rect 331398 460046 331494 460102
rect 330874 459978 331494 460046
rect 330874 459922 330970 459978
rect 331026 459922 331094 459978
rect 331150 459922 331218 459978
rect 331274 459922 331342 459978
rect 331398 459922 331494 459978
rect 330874 458342 331494 459922
rect 345154 597212 345774 598268
rect 345154 597156 345250 597212
rect 345306 597156 345374 597212
rect 345430 597156 345498 597212
rect 345554 597156 345622 597212
rect 345678 597156 345774 597212
rect 345154 597088 345774 597156
rect 345154 597032 345250 597088
rect 345306 597032 345374 597088
rect 345430 597032 345498 597088
rect 345554 597032 345622 597088
rect 345678 597032 345774 597088
rect 345154 596964 345774 597032
rect 345154 596908 345250 596964
rect 345306 596908 345374 596964
rect 345430 596908 345498 596964
rect 345554 596908 345622 596964
rect 345678 596908 345774 596964
rect 345154 596840 345774 596908
rect 345154 596784 345250 596840
rect 345306 596784 345374 596840
rect 345430 596784 345498 596840
rect 345554 596784 345622 596840
rect 345678 596784 345774 596840
rect 345154 580350 345774 596784
rect 345154 580294 345250 580350
rect 345306 580294 345374 580350
rect 345430 580294 345498 580350
rect 345554 580294 345622 580350
rect 345678 580294 345774 580350
rect 345154 580226 345774 580294
rect 345154 580170 345250 580226
rect 345306 580170 345374 580226
rect 345430 580170 345498 580226
rect 345554 580170 345622 580226
rect 345678 580170 345774 580226
rect 345154 580102 345774 580170
rect 345154 580046 345250 580102
rect 345306 580046 345374 580102
rect 345430 580046 345498 580102
rect 345554 580046 345622 580102
rect 345678 580046 345774 580102
rect 345154 579978 345774 580046
rect 345154 579922 345250 579978
rect 345306 579922 345374 579978
rect 345430 579922 345498 579978
rect 345554 579922 345622 579978
rect 345678 579922 345774 579978
rect 345154 562350 345774 579922
rect 345154 562294 345250 562350
rect 345306 562294 345374 562350
rect 345430 562294 345498 562350
rect 345554 562294 345622 562350
rect 345678 562294 345774 562350
rect 345154 562226 345774 562294
rect 345154 562170 345250 562226
rect 345306 562170 345374 562226
rect 345430 562170 345498 562226
rect 345554 562170 345622 562226
rect 345678 562170 345774 562226
rect 345154 562102 345774 562170
rect 345154 562046 345250 562102
rect 345306 562046 345374 562102
rect 345430 562046 345498 562102
rect 345554 562046 345622 562102
rect 345678 562046 345774 562102
rect 345154 561978 345774 562046
rect 345154 561922 345250 561978
rect 345306 561922 345374 561978
rect 345430 561922 345498 561978
rect 345554 561922 345622 561978
rect 345678 561922 345774 561978
rect 345154 544350 345774 561922
rect 345154 544294 345250 544350
rect 345306 544294 345374 544350
rect 345430 544294 345498 544350
rect 345554 544294 345622 544350
rect 345678 544294 345774 544350
rect 345154 544226 345774 544294
rect 345154 544170 345250 544226
rect 345306 544170 345374 544226
rect 345430 544170 345498 544226
rect 345554 544170 345622 544226
rect 345678 544170 345774 544226
rect 345154 544102 345774 544170
rect 345154 544046 345250 544102
rect 345306 544046 345374 544102
rect 345430 544046 345498 544102
rect 345554 544046 345622 544102
rect 345678 544046 345774 544102
rect 345154 543978 345774 544046
rect 345154 543922 345250 543978
rect 345306 543922 345374 543978
rect 345430 543922 345498 543978
rect 345554 543922 345622 543978
rect 345678 543922 345774 543978
rect 345154 526350 345774 543922
rect 345154 526294 345250 526350
rect 345306 526294 345374 526350
rect 345430 526294 345498 526350
rect 345554 526294 345622 526350
rect 345678 526294 345774 526350
rect 345154 526226 345774 526294
rect 345154 526170 345250 526226
rect 345306 526170 345374 526226
rect 345430 526170 345498 526226
rect 345554 526170 345622 526226
rect 345678 526170 345774 526226
rect 345154 526102 345774 526170
rect 345154 526046 345250 526102
rect 345306 526046 345374 526102
rect 345430 526046 345498 526102
rect 345554 526046 345622 526102
rect 345678 526046 345774 526102
rect 345154 525978 345774 526046
rect 345154 525922 345250 525978
rect 345306 525922 345374 525978
rect 345430 525922 345498 525978
rect 345554 525922 345622 525978
rect 345678 525922 345774 525978
rect 345154 508350 345774 525922
rect 345154 508294 345250 508350
rect 345306 508294 345374 508350
rect 345430 508294 345498 508350
rect 345554 508294 345622 508350
rect 345678 508294 345774 508350
rect 345154 508226 345774 508294
rect 345154 508170 345250 508226
rect 345306 508170 345374 508226
rect 345430 508170 345498 508226
rect 345554 508170 345622 508226
rect 345678 508170 345774 508226
rect 345154 508102 345774 508170
rect 345154 508046 345250 508102
rect 345306 508046 345374 508102
rect 345430 508046 345498 508102
rect 345554 508046 345622 508102
rect 345678 508046 345774 508102
rect 345154 507978 345774 508046
rect 345154 507922 345250 507978
rect 345306 507922 345374 507978
rect 345430 507922 345498 507978
rect 345554 507922 345622 507978
rect 345678 507922 345774 507978
rect 345154 490350 345774 507922
rect 345154 490294 345250 490350
rect 345306 490294 345374 490350
rect 345430 490294 345498 490350
rect 345554 490294 345622 490350
rect 345678 490294 345774 490350
rect 345154 490226 345774 490294
rect 345154 490170 345250 490226
rect 345306 490170 345374 490226
rect 345430 490170 345498 490226
rect 345554 490170 345622 490226
rect 345678 490170 345774 490226
rect 345154 490102 345774 490170
rect 345154 490046 345250 490102
rect 345306 490046 345374 490102
rect 345430 490046 345498 490102
rect 345554 490046 345622 490102
rect 345678 490046 345774 490102
rect 345154 489978 345774 490046
rect 345154 489922 345250 489978
rect 345306 489922 345374 489978
rect 345430 489922 345498 489978
rect 345554 489922 345622 489978
rect 345678 489922 345774 489978
rect 345154 472350 345774 489922
rect 345154 472294 345250 472350
rect 345306 472294 345374 472350
rect 345430 472294 345498 472350
rect 345554 472294 345622 472350
rect 345678 472294 345774 472350
rect 345154 472226 345774 472294
rect 345154 472170 345250 472226
rect 345306 472170 345374 472226
rect 345430 472170 345498 472226
rect 345554 472170 345622 472226
rect 345678 472170 345774 472226
rect 345154 472102 345774 472170
rect 345154 472046 345250 472102
rect 345306 472046 345374 472102
rect 345430 472046 345498 472102
rect 345554 472046 345622 472102
rect 345678 472046 345774 472102
rect 345154 471978 345774 472046
rect 345154 471922 345250 471978
rect 345306 471922 345374 471978
rect 345430 471922 345498 471978
rect 345554 471922 345622 471978
rect 345678 471922 345774 471978
rect 345154 458342 345774 471922
rect 348874 598172 349494 598268
rect 348874 598116 348970 598172
rect 349026 598116 349094 598172
rect 349150 598116 349218 598172
rect 349274 598116 349342 598172
rect 349398 598116 349494 598172
rect 348874 598048 349494 598116
rect 348874 597992 348970 598048
rect 349026 597992 349094 598048
rect 349150 597992 349218 598048
rect 349274 597992 349342 598048
rect 349398 597992 349494 598048
rect 348874 597924 349494 597992
rect 348874 597868 348970 597924
rect 349026 597868 349094 597924
rect 349150 597868 349218 597924
rect 349274 597868 349342 597924
rect 349398 597868 349494 597924
rect 348874 597800 349494 597868
rect 348874 597744 348970 597800
rect 349026 597744 349094 597800
rect 349150 597744 349218 597800
rect 349274 597744 349342 597800
rect 349398 597744 349494 597800
rect 348874 586350 349494 597744
rect 348874 586294 348970 586350
rect 349026 586294 349094 586350
rect 349150 586294 349218 586350
rect 349274 586294 349342 586350
rect 349398 586294 349494 586350
rect 348874 586226 349494 586294
rect 348874 586170 348970 586226
rect 349026 586170 349094 586226
rect 349150 586170 349218 586226
rect 349274 586170 349342 586226
rect 349398 586170 349494 586226
rect 348874 586102 349494 586170
rect 348874 586046 348970 586102
rect 349026 586046 349094 586102
rect 349150 586046 349218 586102
rect 349274 586046 349342 586102
rect 349398 586046 349494 586102
rect 348874 585978 349494 586046
rect 348874 585922 348970 585978
rect 349026 585922 349094 585978
rect 349150 585922 349218 585978
rect 349274 585922 349342 585978
rect 349398 585922 349494 585978
rect 348874 568350 349494 585922
rect 348874 568294 348970 568350
rect 349026 568294 349094 568350
rect 349150 568294 349218 568350
rect 349274 568294 349342 568350
rect 349398 568294 349494 568350
rect 348874 568226 349494 568294
rect 348874 568170 348970 568226
rect 349026 568170 349094 568226
rect 349150 568170 349218 568226
rect 349274 568170 349342 568226
rect 349398 568170 349494 568226
rect 348874 568102 349494 568170
rect 348874 568046 348970 568102
rect 349026 568046 349094 568102
rect 349150 568046 349218 568102
rect 349274 568046 349342 568102
rect 349398 568046 349494 568102
rect 348874 567978 349494 568046
rect 348874 567922 348970 567978
rect 349026 567922 349094 567978
rect 349150 567922 349218 567978
rect 349274 567922 349342 567978
rect 349398 567922 349494 567978
rect 348874 550350 349494 567922
rect 348874 550294 348970 550350
rect 349026 550294 349094 550350
rect 349150 550294 349218 550350
rect 349274 550294 349342 550350
rect 349398 550294 349494 550350
rect 348874 550226 349494 550294
rect 348874 550170 348970 550226
rect 349026 550170 349094 550226
rect 349150 550170 349218 550226
rect 349274 550170 349342 550226
rect 349398 550170 349494 550226
rect 348874 550102 349494 550170
rect 348874 550046 348970 550102
rect 349026 550046 349094 550102
rect 349150 550046 349218 550102
rect 349274 550046 349342 550102
rect 349398 550046 349494 550102
rect 348874 549978 349494 550046
rect 348874 549922 348970 549978
rect 349026 549922 349094 549978
rect 349150 549922 349218 549978
rect 349274 549922 349342 549978
rect 349398 549922 349494 549978
rect 348874 532350 349494 549922
rect 348874 532294 348970 532350
rect 349026 532294 349094 532350
rect 349150 532294 349218 532350
rect 349274 532294 349342 532350
rect 349398 532294 349494 532350
rect 348874 532226 349494 532294
rect 348874 532170 348970 532226
rect 349026 532170 349094 532226
rect 349150 532170 349218 532226
rect 349274 532170 349342 532226
rect 349398 532170 349494 532226
rect 348874 532102 349494 532170
rect 348874 532046 348970 532102
rect 349026 532046 349094 532102
rect 349150 532046 349218 532102
rect 349274 532046 349342 532102
rect 349398 532046 349494 532102
rect 348874 531978 349494 532046
rect 348874 531922 348970 531978
rect 349026 531922 349094 531978
rect 349150 531922 349218 531978
rect 349274 531922 349342 531978
rect 349398 531922 349494 531978
rect 348874 514350 349494 531922
rect 348874 514294 348970 514350
rect 349026 514294 349094 514350
rect 349150 514294 349218 514350
rect 349274 514294 349342 514350
rect 349398 514294 349494 514350
rect 348874 514226 349494 514294
rect 348874 514170 348970 514226
rect 349026 514170 349094 514226
rect 349150 514170 349218 514226
rect 349274 514170 349342 514226
rect 349398 514170 349494 514226
rect 348874 514102 349494 514170
rect 348874 514046 348970 514102
rect 349026 514046 349094 514102
rect 349150 514046 349218 514102
rect 349274 514046 349342 514102
rect 349398 514046 349494 514102
rect 348874 513978 349494 514046
rect 348874 513922 348970 513978
rect 349026 513922 349094 513978
rect 349150 513922 349218 513978
rect 349274 513922 349342 513978
rect 349398 513922 349494 513978
rect 348874 496350 349494 513922
rect 348874 496294 348970 496350
rect 349026 496294 349094 496350
rect 349150 496294 349218 496350
rect 349274 496294 349342 496350
rect 349398 496294 349494 496350
rect 348874 496226 349494 496294
rect 348874 496170 348970 496226
rect 349026 496170 349094 496226
rect 349150 496170 349218 496226
rect 349274 496170 349342 496226
rect 349398 496170 349494 496226
rect 348874 496102 349494 496170
rect 348874 496046 348970 496102
rect 349026 496046 349094 496102
rect 349150 496046 349218 496102
rect 349274 496046 349342 496102
rect 349398 496046 349494 496102
rect 348874 495978 349494 496046
rect 348874 495922 348970 495978
rect 349026 495922 349094 495978
rect 349150 495922 349218 495978
rect 349274 495922 349342 495978
rect 349398 495922 349494 495978
rect 348874 478350 349494 495922
rect 348874 478294 348970 478350
rect 349026 478294 349094 478350
rect 349150 478294 349218 478350
rect 349274 478294 349342 478350
rect 349398 478294 349494 478350
rect 348874 478226 349494 478294
rect 348874 478170 348970 478226
rect 349026 478170 349094 478226
rect 349150 478170 349218 478226
rect 349274 478170 349342 478226
rect 349398 478170 349494 478226
rect 348874 478102 349494 478170
rect 348874 478046 348970 478102
rect 349026 478046 349094 478102
rect 349150 478046 349218 478102
rect 349274 478046 349342 478102
rect 349398 478046 349494 478102
rect 348874 477978 349494 478046
rect 348874 477922 348970 477978
rect 349026 477922 349094 477978
rect 349150 477922 349218 477978
rect 349274 477922 349342 477978
rect 349398 477922 349494 477978
rect 348874 460350 349494 477922
rect 348874 460294 348970 460350
rect 349026 460294 349094 460350
rect 349150 460294 349218 460350
rect 349274 460294 349342 460350
rect 349398 460294 349494 460350
rect 348874 460226 349494 460294
rect 348874 460170 348970 460226
rect 349026 460170 349094 460226
rect 349150 460170 349218 460226
rect 349274 460170 349342 460226
rect 349398 460170 349494 460226
rect 348874 460102 349494 460170
rect 348874 460046 348970 460102
rect 349026 460046 349094 460102
rect 349150 460046 349218 460102
rect 349274 460046 349342 460102
rect 349398 460046 349494 460102
rect 348874 459978 349494 460046
rect 348874 459922 348970 459978
rect 349026 459922 349094 459978
rect 349150 459922 349218 459978
rect 349274 459922 349342 459978
rect 349398 459922 349494 459978
rect 348874 458342 349494 459922
rect 363154 597212 363774 598268
rect 363154 597156 363250 597212
rect 363306 597156 363374 597212
rect 363430 597156 363498 597212
rect 363554 597156 363622 597212
rect 363678 597156 363774 597212
rect 363154 597088 363774 597156
rect 363154 597032 363250 597088
rect 363306 597032 363374 597088
rect 363430 597032 363498 597088
rect 363554 597032 363622 597088
rect 363678 597032 363774 597088
rect 363154 596964 363774 597032
rect 363154 596908 363250 596964
rect 363306 596908 363374 596964
rect 363430 596908 363498 596964
rect 363554 596908 363622 596964
rect 363678 596908 363774 596964
rect 363154 596840 363774 596908
rect 363154 596784 363250 596840
rect 363306 596784 363374 596840
rect 363430 596784 363498 596840
rect 363554 596784 363622 596840
rect 363678 596784 363774 596840
rect 363154 580350 363774 596784
rect 363154 580294 363250 580350
rect 363306 580294 363374 580350
rect 363430 580294 363498 580350
rect 363554 580294 363622 580350
rect 363678 580294 363774 580350
rect 363154 580226 363774 580294
rect 363154 580170 363250 580226
rect 363306 580170 363374 580226
rect 363430 580170 363498 580226
rect 363554 580170 363622 580226
rect 363678 580170 363774 580226
rect 363154 580102 363774 580170
rect 363154 580046 363250 580102
rect 363306 580046 363374 580102
rect 363430 580046 363498 580102
rect 363554 580046 363622 580102
rect 363678 580046 363774 580102
rect 363154 579978 363774 580046
rect 363154 579922 363250 579978
rect 363306 579922 363374 579978
rect 363430 579922 363498 579978
rect 363554 579922 363622 579978
rect 363678 579922 363774 579978
rect 363154 562350 363774 579922
rect 363154 562294 363250 562350
rect 363306 562294 363374 562350
rect 363430 562294 363498 562350
rect 363554 562294 363622 562350
rect 363678 562294 363774 562350
rect 363154 562226 363774 562294
rect 363154 562170 363250 562226
rect 363306 562170 363374 562226
rect 363430 562170 363498 562226
rect 363554 562170 363622 562226
rect 363678 562170 363774 562226
rect 363154 562102 363774 562170
rect 363154 562046 363250 562102
rect 363306 562046 363374 562102
rect 363430 562046 363498 562102
rect 363554 562046 363622 562102
rect 363678 562046 363774 562102
rect 363154 561978 363774 562046
rect 363154 561922 363250 561978
rect 363306 561922 363374 561978
rect 363430 561922 363498 561978
rect 363554 561922 363622 561978
rect 363678 561922 363774 561978
rect 363154 544350 363774 561922
rect 363154 544294 363250 544350
rect 363306 544294 363374 544350
rect 363430 544294 363498 544350
rect 363554 544294 363622 544350
rect 363678 544294 363774 544350
rect 363154 544226 363774 544294
rect 363154 544170 363250 544226
rect 363306 544170 363374 544226
rect 363430 544170 363498 544226
rect 363554 544170 363622 544226
rect 363678 544170 363774 544226
rect 363154 544102 363774 544170
rect 363154 544046 363250 544102
rect 363306 544046 363374 544102
rect 363430 544046 363498 544102
rect 363554 544046 363622 544102
rect 363678 544046 363774 544102
rect 363154 543978 363774 544046
rect 363154 543922 363250 543978
rect 363306 543922 363374 543978
rect 363430 543922 363498 543978
rect 363554 543922 363622 543978
rect 363678 543922 363774 543978
rect 363154 526350 363774 543922
rect 363154 526294 363250 526350
rect 363306 526294 363374 526350
rect 363430 526294 363498 526350
rect 363554 526294 363622 526350
rect 363678 526294 363774 526350
rect 363154 526226 363774 526294
rect 363154 526170 363250 526226
rect 363306 526170 363374 526226
rect 363430 526170 363498 526226
rect 363554 526170 363622 526226
rect 363678 526170 363774 526226
rect 363154 526102 363774 526170
rect 363154 526046 363250 526102
rect 363306 526046 363374 526102
rect 363430 526046 363498 526102
rect 363554 526046 363622 526102
rect 363678 526046 363774 526102
rect 363154 525978 363774 526046
rect 363154 525922 363250 525978
rect 363306 525922 363374 525978
rect 363430 525922 363498 525978
rect 363554 525922 363622 525978
rect 363678 525922 363774 525978
rect 363154 508350 363774 525922
rect 363154 508294 363250 508350
rect 363306 508294 363374 508350
rect 363430 508294 363498 508350
rect 363554 508294 363622 508350
rect 363678 508294 363774 508350
rect 363154 508226 363774 508294
rect 363154 508170 363250 508226
rect 363306 508170 363374 508226
rect 363430 508170 363498 508226
rect 363554 508170 363622 508226
rect 363678 508170 363774 508226
rect 363154 508102 363774 508170
rect 363154 508046 363250 508102
rect 363306 508046 363374 508102
rect 363430 508046 363498 508102
rect 363554 508046 363622 508102
rect 363678 508046 363774 508102
rect 363154 507978 363774 508046
rect 363154 507922 363250 507978
rect 363306 507922 363374 507978
rect 363430 507922 363498 507978
rect 363554 507922 363622 507978
rect 363678 507922 363774 507978
rect 363154 490350 363774 507922
rect 363154 490294 363250 490350
rect 363306 490294 363374 490350
rect 363430 490294 363498 490350
rect 363554 490294 363622 490350
rect 363678 490294 363774 490350
rect 363154 490226 363774 490294
rect 363154 490170 363250 490226
rect 363306 490170 363374 490226
rect 363430 490170 363498 490226
rect 363554 490170 363622 490226
rect 363678 490170 363774 490226
rect 363154 490102 363774 490170
rect 363154 490046 363250 490102
rect 363306 490046 363374 490102
rect 363430 490046 363498 490102
rect 363554 490046 363622 490102
rect 363678 490046 363774 490102
rect 363154 489978 363774 490046
rect 363154 489922 363250 489978
rect 363306 489922 363374 489978
rect 363430 489922 363498 489978
rect 363554 489922 363622 489978
rect 363678 489922 363774 489978
rect 363154 472350 363774 489922
rect 363154 472294 363250 472350
rect 363306 472294 363374 472350
rect 363430 472294 363498 472350
rect 363554 472294 363622 472350
rect 363678 472294 363774 472350
rect 363154 472226 363774 472294
rect 363154 472170 363250 472226
rect 363306 472170 363374 472226
rect 363430 472170 363498 472226
rect 363554 472170 363622 472226
rect 363678 472170 363774 472226
rect 363154 472102 363774 472170
rect 363154 472046 363250 472102
rect 363306 472046 363374 472102
rect 363430 472046 363498 472102
rect 363554 472046 363622 472102
rect 363678 472046 363774 472102
rect 363154 471978 363774 472046
rect 363154 471922 363250 471978
rect 363306 471922 363374 471978
rect 363430 471922 363498 471978
rect 363554 471922 363622 471978
rect 363678 471922 363774 471978
rect 363154 458342 363774 471922
rect 366874 598172 367494 598268
rect 366874 598116 366970 598172
rect 367026 598116 367094 598172
rect 367150 598116 367218 598172
rect 367274 598116 367342 598172
rect 367398 598116 367494 598172
rect 366874 598048 367494 598116
rect 366874 597992 366970 598048
rect 367026 597992 367094 598048
rect 367150 597992 367218 598048
rect 367274 597992 367342 598048
rect 367398 597992 367494 598048
rect 366874 597924 367494 597992
rect 366874 597868 366970 597924
rect 367026 597868 367094 597924
rect 367150 597868 367218 597924
rect 367274 597868 367342 597924
rect 367398 597868 367494 597924
rect 366874 597800 367494 597868
rect 366874 597744 366970 597800
rect 367026 597744 367094 597800
rect 367150 597744 367218 597800
rect 367274 597744 367342 597800
rect 367398 597744 367494 597800
rect 366874 586350 367494 597744
rect 366874 586294 366970 586350
rect 367026 586294 367094 586350
rect 367150 586294 367218 586350
rect 367274 586294 367342 586350
rect 367398 586294 367494 586350
rect 366874 586226 367494 586294
rect 366874 586170 366970 586226
rect 367026 586170 367094 586226
rect 367150 586170 367218 586226
rect 367274 586170 367342 586226
rect 367398 586170 367494 586226
rect 366874 586102 367494 586170
rect 366874 586046 366970 586102
rect 367026 586046 367094 586102
rect 367150 586046 367218 586102
rect 367274 586046 367342 586102
rect 367398 586046 367494 586102
rect 366874 585978 367494 586046
rect 366874 585922 366970 585978
rect 367026 585922 367094 585978
rect 367150 585922 367218 585978
rect 367274 585922 367342 585978
rect 367398 585922 367494 585978
rect 366874 568350 367494 585922
rect 366874 568294 366970 568350
rect 367026 568294 367094 568350
rect 367150 568294 367218 568350
rect 367274 568294 367342 568350
rect 367398 568294 367494 568350
rect 366874 568226 367494 568294
rect 366874 568170 366970 568226
rect 367026 568170 367094 568226
rect 367150 568170 367218 568226
rect 367274 568170 367342 568226
rect 367398 568170 367494 568226
rect 366874 568102 367494 568170
rect 366874 568046 366970 568102
rect 367026 568046 367094 568102
rect 367150 568046 367218 568102
rect 367274 568046 367342 568102
rect 367398 568046 367494 568102
rect 366874 567978 367494 568046
rect 366874 567922 366970 567978
rect 367026 567922 367094 567978
rect 367150 567922 367218 567978
rect 367274 567922 367342 567978
rect 367398 567922 367494 567978
rect 366874 550350 367494 567922
rect 366874 550294 366970 550350
rect 367026 550294 367094 550350
rect 367150 550294 367218 550350
rect 367274 550294 367342 550350
rect 367398 550294 367494 550350
rect 366874 550226 367494 550294
rect 366874 550170 366970 550226
rect 367026 550170 367094 550226
rect 367150 550170 367218 550226
rect 367274 550170 367342 550226
rect 367398 550170 367494 550226
rect 366874 550102 367494 550170
rect 366874 550046 366970 550102
rect 367026 550046 367094 550102
rect 367150 550046 367218 550102
rect 367274 550046 367342 550102
rect 367398 550046 367494 550102
rect 366874 549978 367494 550046
rect 366874 549922 366970 549978
rect 367026 549922 367094 549978
rect 367150 549922 367218 549978
rect 367274 549922 367342 549978
rect 367398 549922 367494 549978
rect 366874 532350 367494 549922
rect 366874 532294 366970 532350
rect 367026 532294 367094 532350
rect 367150 532294 367218 532350
rect 367274 532294 367342 532350
rect 367398 532294 367494 532350
rect 366874 532226 367494 532294
rect 366874 532170 366970 532226
rect 367026 532170 367094 532226
rect 367150 532170 367218 532226
rect 367274 532170 367342 532226
rect 367398 532170 367494 532226
rect 366874 532102 367494 532170
rect 366874 532046 366970 532102
rect 367026 532046 367094 532102
rect 367150 532046 367218 532102
rect 367274 532046 367342 532102
rect 367398 532046 367494 532102
rect 366874 531978 367494 532046
rect 366874 531922 366970 531978
rect 367026 531922 367094 531978
rect 367150 531922 367218 531978
rect 367274 531922 367342 531978
rect 367398 531922 367494 531978
rect 366874 514350 367494 531922
rect 366874 514294 366970 514350
rect 367026 514294 367094 514350
rect 367150 514294 367218 514350
rect 367274 514294 367342 514350
rect 367398 514294 367494 514350
rect 366874 514226 367494 514294
rect 366874 514170 366970 514226
rect 367026 514170 367094 514226
rect 367150 514170 367218 514226
rect 367274 514170 367342 514226
rect 367398 514170 367494 514226
rect 366874 514102 367494 514170
rect 366874 514046 366970 514102
rect 367026 514046 367094 514102
rect 367150 514046 367218 514102
rect 367274 514046 367342 514102
rect 367398 514046 367494 514102
rect 366874 513978 367494 514046
rect 366874 513922 366970 513978
rect 367026 513922 367094 513978
rect 367150 513922 367218 513978
rect 367274 513922 367342 513978
rect 367398 513922 367494 513978
rect 366874 496350 367494 513922
rect 366874 496294 366970 496350
rect 367026 496294 367094 496350
rect 367150 496294 367218 496350
rect 367274 496294 367342 496350
rect 367398 496294 367494 496350
rect 366874 496226 367494 496294
rect 366874 496170 366970 496226
rect 367026 496170 367094 496226
rect 367150 496170 367218 496226
rect 367274 496170 367342 496226
rect 367398 496170 367494 496226
rect 366874 496102 367494 496170
rect 366874 496046 366970 496102
rect 367026 496046 367094 496102
rect 367150 496046 367218 496102
rect 367274 496046 367342 496102
rect 367398 496046 367494 496102
rect 366874 495978 367494 496046
rect 366874 495922 366970 495978
rect 367026 495922 367094 495978
rect 367150 495922 367218 495978
rect 367274 495922 367342 495978
rect 367398 495922 367494 495978
rect 366874 478350 367494 495922
rect 366874 478294 366970 478350
rect 367026 478294 367094 478350
rect 367150 478294 367218 478350
rect 367274 478294 367342 478350
rect 367398 478294 367494 478350
rect 366874 478226 367494 478294
rect 366874 478170 366970 478226
rect 367026 478170 367094 478226
rect 367150 478170 367218 478226
rect 367274 478170 367342 478226
rect 367398 478170 367494 478226
rect 366874 478102 367494 478170
rect 366874 478046 366970 478102
rect 367026 478046 367094 478102
rect 367150 478046 367218 478102
rect 367274 478046 367342 478102
rect 367398 478046 367494 478102
rect 366874 477978 367494 478046
rect 366874 477922 366970 477978
rect 367026 477922 367094 477978
rect 367150 477922 367218 477978
rect 367274 477922 367342 477978
rect 367398 477922 367494 477978
rect 366874 460350 367494 477922
rect 366874 460294 366970 460350
rect 367026 460294 367094 460350
rect 367150 460294 367218 460350
rect 367274 460294 367342 460350
rect 367398 460294 367494 460350
rect 366874 460226 367494 460294
rect 366874 460170 366970 460226
rect 367026 460170 367094 460226
rect 367150 460170 367218 460226
rect 367274 460170 367342 460226
rect 367398 460170 367494 460226
rect 366874 460102 367494 460170
rect 366874 460046 366970 460102
rect 367026 460046 367094 460102
rect 367150 460046 367218 460102
rect 367274 460046 367342 460102
rect 367398 460046 367494 460102
rect 366874 459978 367494 460046
rect 366874 459922 366970 459978
rect 367026 459922 367094 459978
rect 367150 459922 367218 459978
rect 367274 459922 367342 459978
rect 367398 459922 367494 459978
rect 366874 458342 367494 459922
rect 381154 597212 381774 598268
rect 381154 597156 381250 597212
rect 381306 597156 381374 597212
rect 381430 597156 381498 597212
rect 381554 597156 381622 597212
rect 381678 597156 381774 597212
rect 381154 597088 381774 597156
rect 381154 597032 381250 597088
rect 381306 597032 381374 597088
rect 381430 597032 381498 597088
rect 381554 597032 381622 597088
rect 381678 597032 381774 597088
rect 381154 596964 381774 597032
rect 381154 596908 381250 596964
rect 381306 596908 381374 596964
rect 381430 596908 381498 596964
rect 381554 596908 381622 596964
rect 381678 596908 381774 596964
rect 381154 596840 381774 596908
rect 381154 596784 381250 596840
rect 381306 596784 381374 596840
rect 381430 596784 381498 596840
rect 381554 596784 381622 596840
rect 381678 596784 381774 596840
rect 381154 580350 381774 596784
rect 381154 580294 381250 580350
rect 381306 580294 381374 580350
rect 381430 580294 381498 580350
rect 381554 580294 381622 580350
rect 381678 580294 381774 580350
rect 381154 580226 381774 580294
rect 381154 580170 381250 580226
rect 381306 580170 381374 580226
rect 381430 580170 381498 580226
rect 381554 580170 381622 580226
rect 381678 580170 381774 580226
rect 381154 580102 381774 580170
rect 381154 580046 381250 580102
rect 381306 580046 381374 580102
rect 381430 580046 381498 580102
rect 381554 580046 381622 580102
rect 381678 580046 381774 580102
rect 381154 579978 381774 580046
rect 381154 579922 381250 579978
rect 381306 579922 381374 579978
rect 381430 579922 381498 579978
rect 381554 579922 381622 579978
rect 381678 579922 381774 579978
rect 381154 562350 381774 579922
rect 381154 562294 381250 562350
rect 381306 562294 381374 562350
rect 381430 562294 381498 562350
rect 381554 562294 381622 562350
rect 381678 562294 381774 562350
rect 381154 562226 381774 562294
rect 381154 562170 381250 562226
rect 381306 562170 381374 562226
rect 381430 562170 381498 562226
rect 381554 562170 381622 562226
rect 381678 562170 381774 562226
rect 381154 562102 381774 562170
rect 381154 562046 381250 562102
rect 381306 562046 381374 562102
rect 381430 562046 381498 562102
rect 381554 562046 381622 562102
rect 381678 562046 381774 562102
rect 381154 561978 381774 562046
rect 381154 561922 381250 561978
rect 381306 561922 381374 561978
rect 381430 561922 381498 561978
rect 381554 561922 381622 561978
rect 381678 561922 381774 561978
rect 381154 544350 381774 561922
rect 381154 544294 381250 544350
rect 381306 544294 381374 544350
rect 381430 544294 381498 544350
rect 381554 544294 381622 544350
rect 381678 544294 381774 544350
rect 381154 544226 381774 544294
rect 381154 544170 381250 544226
rect 381306 544170 381374 544226
rect 381430 544170 381498 544226
rect 381554 544170 381622 544226
rect 381678 544170 381774 544226
rect 381154 544102 381774 544170
rect 381154 544046 381250 544102
rect 381306 544046 381374 544102
rect 381430 544046 381498 544102
rect 381554 544046 381622 544102
rect 381678 544046 381774 544102
rect 381154 543978 381774 544046
rect 381154 543922 381250 543978
rect 381306 543922 381374 543978
rect 381430 543922 381498 543978
rect 381554 543922 381622 543978
rect 381678 543922 381774 543978
rect 381154 526350 381774 543922
rect 381154 526294 381250 526350
rect 381306 526294 381374 526350
rect 381430 526294 381498 526350
rect 381554 526294 381622 526350
rect 381678 526294 381774 526350
rect 381154 526226 381774 526294
rect 381154 526170 381250 526226
rect 381306 526170 381374 526226
rect 381430 526170 381498 526226
rect 381554 526170 381622 526226
rect 381678 526170 381774 526226
rect 381154 526102 381774 526170
rect 381154 526046 381250 526102
rect 381306 526046 381374 526102
rect 381430 526046 381498 526102
rect 381554 526046 381622 526102
rect 381678 526046 381774 526102
rect 381154 525978 381774 526046
rect 381154 525922 381250 525978
rect 381306 525922 381374 525978
rect 381430 525922 381498 525978
rect 381554 525922 381622 525978
rect 381678 525922 381774 525978
rect 381154 508350 381774 525922
rect 381154 508294 381250 508350
rect 381306 508294 381374 508350
rect 381430 508294 381498 508350
rect 381554 508294 381622 508350
rect 381678 508294 381774 508350
rect 381154 508226 381774 508294
rect 381154 508170 381250 508226
rect 381306 508170 381374 508226
rect 381430 508170 381498 508226
rect 381554 508170 381622 508226
rect 381678 508170 381774 508226
rect 381154 508102 381774 508170
rect 381154 508046 381250 508102
rect 381306 508046 381374 508102
rect 381430 508046 381498 508102
rect 381554 508046 381622 508102
rect 381678 508046 381774 508102
rect 381154 507978 381774 508046
rect 381154 507922 381250 507978
rect 381306 507922 381374 507978
rect 381430 507922 381498 507978
rect 381554 507922 381622 507978
rect 381678 507922 381774 507978
rect 381154 490350 381774 507922
rect 381154 490294 381250 490350
rect 381306 490294 381374 490350
rect 381430 490294 381498 490350
rect 381554 490294 381622 490350
rect 381678 490294 381774 490350
rect 381154 490226 381774 490294
rect 381154 490170 381250 490226
rect 381306 490170 381374 490226
rect 381430 490170 381498 490226
rect 381554 490170 381622 490226
rect 381678 490170 381774 490226
rect 381154 490102 381774 490170
rect 381154 490046 381250 490102
rect 381306 490046 381374 490102
rect 381430 490046 381498 490102
rect 381554 490046 381622 490102
rect 381678 490046 381774 490102
rect 381154 489978 381774 490046
rect 381154 489922 381250 489978
rect 381306 489922 381374 489978
rect 381430 489922 381498 489978
rect 381554 489922 381622 489978
rect 381678 489922 381774 489978
rect 381154 472350 381774 489922
rect 381154 472294 381250 472350
rect 381306 472294 381374 472350
rect 381430 472294 381498 472350
rect 381554 472294 381622 472350
rect 381678 472294 381774 472350
rect 381154 472226 381774 472294
rect 381154 472170 381250 472226
rect 381306 472170 381374 472226
rect 381430 472170 381498 472226
rect 381554 472170 381622 472226
rect 381678 472170 381774 472226
rect 381154 472102 381774 472170
rect 381154 472046 381250 472102
rect 381306 472046 381374 472102
rect 381430 472046 381498 472102
rect 381554 472046 381622 472102
rect 381678 472046 381774 472102
rect 381154 471978 381774 472046
rect 381154 471922 381250 471978
rect 381306 471922 381374 471978
rect 381430 471922 381498 471978
rect 381554 471922 381622 471978
rect 381678 471922 381774 471978
rect 204874 442294 204970 442350
rect 205026 442294 205094 442350
rect 205150 442294 205218 442350
rect 205274 442294 205342 442350
rect 205398 442294 205494 442350
rect 204874 442226 205494 442294
rect 204874 442170 204970 442226
rect 205026 442170 205094 442226
rect 205150 442170 205218 442226
rect 205274 442170 205342 442226
rect 205398 442170 205494 442226
rect 204874 442102 205494 442170
rect 204874 442046 204970 442102
rect 205026 442046 205094 442102
rect 205150 442046 205218 442102
rect 205274 442046 205342 442102
rect 205398 442046 205494 442102
rect 204874 441978 205494 442046
rect 204874 441922 204970 441978
rect 205026 441922 205094 441978
rect 205150 441922 205218 441978
rect 205274 441922 205342 441978
rect 205398 441922 205494 441978
rect 204874 424350 205494 441922
rect 204874 424294 204970 424350
rect 205026 424294 205094 424350
rect 205150 424294 205218 424350
rect 205274 424294 205342 424350
rect 205398 424294 205494 424350
rect 204874 424226 205494 424294
rect 204874 424170 204970 424226
rect 205026 424170 205094 424226
rect 205150 424170 205218 424226
rect 205274 424170 205342 424226
rect 205398 424170 205494 424226
rect 204874 424102 205494 424170
rect 204874 424046 204970 424102
rect 205026 424046 205094 424102
rect 205150 424046 205218 424102
rect 205274 424046 205342 424102
rect 205398 424046 205494 424102
rect 204874 423978 205494 424046
rect 204874 423922 204970 423978
rect 205026 423922 205094 423978
rect 205150 423922 205218 423978
rect 205274 423922 205342 423978
rect 205398 423922 205494 423978
rect 204874 406350 205494 423922
rect 204874 406294 204970 406350
rect 205026 406294 205094 406350
rect 205150 406294 205218 406350
rect 205274 406294 205342 406350
rect 205398 406294 205494 406350
rect 204874 406226 205494 406294
rect 204874 406170 204970 406226
rect 205026 406170 205094 406226
rect 205150 406170 205218 406226
rect 205274 406170 205342 406226
rect 205398 406170 205494 406226
rect 204874 406102 205494 406170
rect 204874 406046 204970 406102
rect 205026 406046 205094 406102
rect 205150 406046 205218 406102
rect 205274 406046 205342 406102
rect 205398 406046 205494 406102
rect 204874 405978 205494 406046
rect 204874 405922 204970 405978
rect 205026 405922 205094 405978
rect 205150 405922 205218 405978
rect 205274 405922 205342 405978
rect 205398 405922 205494 405978
rect 204874 388350 205494 405922
rect 204874 388294 204970 388350
rect 205026 388294 205094 388350
rect 205150 388294 205218 388350
rect 205274 388294 205342 388350
rect 205398 388294 205494 388350
rect 204874 388226 205494 388294
rect 204874 388170 204970 388226
rect 205026 388170 205094 388226
rect 205150 388170 205218 388226
rect 205274 388170 205342 388226
rect 205398 388170 205494 388226
rect 204874 388102 205494 388170
rect 204874 388046 204970 388102
rect 205026 388046 205094 388102
rect 205150 388046 205218 388102
rect 205274 388046 205342 388102
rect 205398 388046 205494 388102
rect 204874 387978 205494 388046
rect 204874 387922 204970 387978
rect 205026 387922 205094 387978
rect 205150 387922 205218 387978
rect 205274 387922 205342 387978
rect 205398 387922 205494 387978
rect 204874 370350 205494 387922
rect 204874 370294 204970 370350
rect 205026 370294 205094 370350
rect 205150 370294 205218 370350
rect 205274 370294 205342 370350
rect 205398 370294 205494 370350
rect 204874 370226 205494 370294
rect 204874 370170 204970 370226
rect 205026 370170 205094 370226
rect 205150 370170 205218 370226
rect 205274 370170 205342 370226
rect 205398 370170 205494 370226
rect 204874 370102 205494 370170
rect 204874 370046 204970 370102
rect 205026 370046 205094 370102
rect 205150 370046 205218 370102
rect 205274 370046 205342 370102
rect 205398 370046 205494 370102
rect 204874 369978 205494 370046
rect 204874 369922 204970 369978
rect 205026 369922 205094 369978
rect 205150 369922 205218 369978
rect 205274 369922 205342 369978
rect 205398 369922 205494 369978
rect 204874 352350 205494 369922
rect 204874 352294 204970 352350
rect 205026 352294 205094 352350
rect 205150 352294 205218 352350
rect 205274 352294 205342 352350
rect 205398 352294 205494 352350
rect 204874 352226 205494 352294
rect 204874 352170 204970 352226
rect 205026 352170 205094 352226
rect 205150 352170 205218 352226
rect 205274 352170 205342 352226
rect 205398 352170 205494 352226
rect 204874 352102 205494 352170
rect 204874 352046 204970 352102
rect 205026 352046 205094 352102
rect 205150 352046 205218 352102
rect 205274 352046 205342 352102
rect 205398 352046 205494 352102
rect 204874 351978 205494 352046
rect 204874 351922 204970 351978
rect 205026 351922 205094 351978
rect 205150 351922 205218 351978
rect 205274 351922 205342 351978
rect 205398 351922 205494 351978
rect 204874 334350 205494 351922
rect 204874 334294 204970 334350
rect 205026 334294 205094 334350
rect 205150 334294 205218 334350
rect 205274 334294 205342 334350
rect 205398 334294 205494 334350
rect 204874 334226 205494 334294
rect 204874 334170 204970 334226
rect 205026 334170 205094 334226
rect 205150 334170 205218 334226
rect 205274 334170 205342 334226
rect 205398 334170 205494 334226
rect 204874 334102 205494 334170
rect 204874 334046 204970 334102
rect 205026 334046 205094 334102
rect 205150 334046 205218 334102
rect 205274 334046 205342 334102
rect 205398 334046 205494 334102
rect 204874 333978 205494 334046
rect 204874 333922 204970 333978
rect 205026 333922 205094 333978
rect 205150 333922 205218 333978
rect 205274 333922 205342 333978
rect 205398 333922 205494 333978
rect 204874 316350 205494 333922
rect 381154 454350 381774 471922
rect 381154 454294 381250 454350
rect 381306 454294 381374 454350
rect 381430 454294 381498 454350
rect 381554 454294 381622 454350
rect 381678 454294 381774 454350
rect 381154 454226 381774 454294
rect 381154 454170 381250 454226
rect 381306 454170 381374 454226
rect 381430 454170 381498 454226
rect 381554 454170 381622 454226
rect 381678 454170 381774 454226
rect 381154 454102 381774 454170
rect 381154 454046 381250 454102
rect 381306 454046 381374 454102
rect 381430 454046 381498 454102
rect 381554 454046 381622 454102
rect 381678 454046 381774 454102
rect 381154 453978 381774 454046
rect 381154 453922 381250 453978
rect 381306 453922 381374 453978
rect 381430 453922 381498 453978
rect 381554 453922 381622 453978
rect 381678 453922 381774 453978
rect 381154 436350 381774 453922
rect 381154 436294 381250 436350
rect 381306 436294 381374 436350
rect 381430 436294 381498 436350
rect 381554 436294 381622 436350
rect 381678 436294 381774 436350
rect 381154 436226 381774 436294
rect 381154 436170 381250 436226
rect 381306 436170 381374 436226
rect 381430 436170 381498 436226
rect 381554 436170 381622 436226
rect 381678 436170 381774 436226
rect 381154 436102 381774 436170
rect 381154 436046 381250 436102
rect 381306 436046 381374 436102
rect 381430 436046 381498 436102
rect 381554 436046 381622 436102
rect 381678 436046 381774 436102
rect 381154 435978 381774 436046
rect 381154 435922 381250 435978
rect 381306 435922 381374 435978
rect 381430 435922 381498 435978
rect 381554 435922 381622 435978
rect 381678 435922 381774 435978
rect 381154 418350 381774 435922
rect 381154 418294 381250 418350
rect 381306 418294 381374 418350
rect 381430 418294 381498 418350
rect 381554 418294 381622 418350
rect 381678 418294 381774 418350
rect 381154 418226 381774 418294
rect 381154 418170 381250 418226
rect 381306 418170 381374 418226
rect 381430 418170 381498 418226
rect 381554 418170 381622 418226
rect 381678 418170 381774 418226
rect 381154 418102 381774 418170
rect 381154 418046 381250 418102
rect 381306 418046 381374 418102
rect 381430 418046 381498 418102
rect 381554 418046 381622 418102
rect 381678 418046 381774 418102
rect 381154 417978 381774 418046
rect 381154 417922 381250 417978
rect 381306 417922 381374 417978
rect 381430 417922 381498 417978
rect 381554 417922 381622 417978
rect 381678 417922 381774 417978
rect 381154 400350 381774 417922
rect 381154 400294 381250 400350
rect 381306 400294 381374 400350
rect 381430 400294 381498 400350
rect 381554 400294 381622 400350
rect 381678 400294 381774 400350
rect 381154 400226 381774 400294
rect 381154 400170 381250 400226
rect 381306 400170 381374 400226
rect 381430 400170 381498 400226
rect 381554 400170 381622 400226
rect 381678 400170 381774 400226
rect 381154 400102 381774 400170
rect 381154 400046 381250 400102
rect 381306 400046 381374 400102
rect 381430 400046 381498 400102
rect 381554 400046 381622 400102
rect 381678 400046 381774 400102
rect 381154 399978 381774 400046
rect 381154 399922 381250 399978
rect 381306 399922 381374 399978
rect 381430 399922 381498 399978
rect 381554 399922 381622 399978
rect 381678 399922 381774 399978
rect 381154 382350 381774 399922
rect 381154 382294 381250 382350
rect 381306 382294 381374 382350
rect 381430 382294 381498 382350
rect 381554 382294 381622 382350
rect 381678 382294 381774 382350
rect 381154 382226 381774 382294
rect 381154 382170 381250 382226
rect 381306 382170 381374 382226
rect 381430 382170 381498 382226
rect 381554 382170 381622 382226
rect 381678 382170 381774 382226
rect 381154 382102 381774 382170
rect 381154 382046 381250 382102
rect 381306 382046 381374 382102
rect 381430 382046 381498 382102
rect 381554 382046 381622 382102
rect 381678 382046 381774 382102
rect 381154 381978 381774 382046
rect 381154 381922 381250 381978
rect 381306 381922 381374 381978
rect 381430 381922 381498 381978
rect 381554 381922 381622 381978
rect 381678 381922 381774 381978
rect 381154 364350 381774 381922
rect 381154 364294 381250 364350
rect 381306 364294 381374 364350
rect 381430 364294 381498 364350
rect 381554 364294 381622 364350
rect 381678 364294 381774 364350
rect 381154 364226 381774 364294
rect 381154 364170 381250 364226
rect 381306 364170 381374 364226
rect 381430 364170 381498 364226
rect 381554 364170 381622 364226
rect 381678 364170 381774 364226
rect 381154 364102 381774 364170
rect 381154 364046 381250 364102
rect 381306 364046 381374 364102
rect 381430 364046 381498 364102
rect 381554 364046 381622 364102
rect 381678 364046 381774 364102
rect 381154 363978 381774 364046
rect 381154 363922 381250 363978
rect 381306 363922 381374 363978
rect 381430 363922 381498 363978
rect 381554 363922 381622 363978
rect 381678 363922 381774 363978
rect 381154 346350 381774 363922
rect 381154 346294 381250 346350
rect 381306 346294 381374 346350
rect 381430 346294 381498 346350
rect 381554 346294 381622 346350
rect 381678 346294 381774 346350
rect 381154 346226 381774 346294
rect 381154 346170 381250 346226
rect 381306 346170 381374 346226
rect 381430 346170 381498 346226
rect 381554 346170 381622 346226
rect 381678 346170 381774 346226
rect 381154 346102 381774 346170
rect 381154 346046 381250 346102
rect 381306 346046 381374 346102
rect 381430 346046 381498 346102
rect 381554 346046 381622 346102
rect 381678 346046 381774 346102
rect 381154 345978 381774 346046
rect 381154 345922 381250 345978
rect 381306 345922 381374 345978
rect 381430 345922 381498 345978
rect 381554 345922 381622 345978
rect 381678 345922 381774 345978
rect 381154 328350 381774 345922
rect 381154 328294 381250 328350
rect 381306 328294 381374 328350
rect 381430 328294 381498 328350
rect 381554 328294 381622 328350
rect 381678 328294 381774 328350
rect 381154 328226 381774 328294
rect 381154 328170 381250 328226
rect 381306 328170 381374 328226
rect 381430 328170 381498 328226
rect 381554 328170 381622 328226
rect 381678 328170 381774 328226
rect 381154 328102 381774 328170
rect 381154 328046 381250 328102
rect 381306 328046 381374 328102
rect 381430 328046 381498 328102
rect 381554 328046 381622 328102
rect 381678 328046 381774 328102
rect 381154 327978 381774 328046
rect 381154 327922 381250 327978
rect 381306 327922 381374 327978
rect 381430 327922 381498 327978
rect 381554 327922 381622 327978
rect 381678 327922 381774 327978
rect 204874 316294 204970 316350
rect 205026 316294 205094 316350
rect 205150 316294 205218 316350
rect 205274 316294 205342 316350
rect 205398 316294 205494 316350
rect 204874 316226 205494 316294
rect 204874 316170 204970 316226
rect 205026 316170 205094 316226
rect 205150 316170 205218 316226
rect 205274 316170 205342 316226
rect 205398 316170 205494 316226
rect 204874 316102 205494 316170
rect 204874 316046 204970 316102
rect 205026 316046 205094 316102
rect 205150 316046 205218 316102
rect 205274 316046 205342 316102
rect 205398 316046 205494 316102
rect 204874 315978 205494 316046
rect 204874 315922 204970 315978
rect 205026 315922 205094 315978
rect 205150 315922 205218 315978
rect 205274 315922 205342 315978
rect 205398 315922 205494 315978
rect 204874 298350 205494 315922
rect 204874 298294 204970 298350
rect 205026 298294 205094 298350
rect 205150 298294 205218 298350
rect 205274 298294 205342 298350
rect 205398 298294 205494 298350
rect 222874 316350 223494 318858
rect 222874 316294 222970 316350
rect 223026 316294 223094 316350
rect 223150 316294 223218 316350
rect 223274 316294 223342 316350
rect 223398 316294 223494 316350
rect 222874 316226 223494 316294
rect 222874 316170 222970 316226
rect 223026 316170 223094 316226
rect 223150 316170 223218 316226
rect 223274 316170 223342 316226
rect 223398 316170 223494 316226
rect 222874 316102 223494 316170
rect 222874 316046 222970 316102
rect 223026 316046 223094 316102
rect 223150 316046 223218 316102
rect 223274 316046 223342 316102
rect 223398 316046 223494 316102
rect 222874 315978 223494 316046
rect 222874 315922 222970 315978
rect 223026 315922 223094 315978
rect 223150 315922 223218 315978
rect 223274 315922 223342 315978
rect 223398 315922 223494 315978
rect 222874 298422 223494 315922
rect 222874 298366 222970 298422
rect 223026 298366 223094 298422
rect 223150 298366 223218 298422
rect 223274 298366 223342 298422
rect 223398 298366 223494 298422
rect 222874 298342 223494 298366
rect 240874 316350 241494 318858
rect 240874 316294 240970 316350
rect 241026 316294 241094 316350
rect 241150 316294 241218 316350
rect 241274 316294 241342 316350
rect 241398 316294 241494 316350
rect 240874 316226 241494 316294
rect 240874 316170 240970 316226
rect 241026 316170 241094 316226
rect 241150 316170 241218 316226
rect 241274 316170 241342 316226
rect 241398 316170 241494 316226
rect 240874 316102 241494 316170
rect 240874 316046 240970 316102
rect 241026 316046 241094 316102
rect 241150 316046 241218 316102
rect 241274 316046 241342 316102
rect 241398 316046 241494 316102
rect 240874 315978 241494 316046
rect 240874 315922 240970 315978
rect 241026 315922 241094 315978
rect 241150 315922 241218 315978
rect 241274 315922 241342 315978
rect 241398 315922 241494 315978
rect 240874 298422 241494 315922
rect 240874 298366 240970 298422
rect 241026 298366 241094 298422
rect 241150 298366 241218 298422
rect 241274 298366 241342 298422
rect 241398 298366 241494 298422
rect 240874 298342 241494 298366
rect 258874 316350 259494 318858
rect 258874 316294 258970 316350
rect 259026 316294 259094 316350
rect 259150 316294 259218 316350
rect 259274 316294 259342 316350
rect 259398 316294 259494 316350
rect 258874 316226 259494 316294
rect 258874 316170 258970 316226
rect 259026 316170 259094 316226
rect 259150 316170 259218 316226
rect 259274 316170 259342 316226
rect 259398 316170 259494 316226
rect 258874 316102 259494 316170
rect 258874 316046 258970 316102
rect 259026 316046 259094 316102
rect 259150 316046 259218 316102
rect 259274 316046 259342 316102
rect 259398 316046 259494 316102
rect 258874 315978 259494 316046
rect 258874 315922 258970 315978
rect 259026 315922 259094 315978
rect 259150 315922 259218 315978
rect 259274 315922 259342 315978
rect 259398 315922 259494 315978
rect 258874 298422 259494 315922
rect 258874 298366 258970 298422
rect 259026 298366 259094 298422
rect 259150 298366 259218 298422
rect 259274 298366 259342 298422
rect 259398 298366 259494 298422
rect 258874 298342 259494 298366
rect 276874 316350 277494 318858
rect 276874 316294 276970 316350
rect 277026 316294 277094 316350
rect 277150 316294 277218 316350
rect 277274 316294 277342 316350
rect 277398 316294 277494 316350
rect 276874 316226 277494 316294
rect 276874 316170 276970 316226
rect 277026 316170 277094 316226
rect 277150 316170 277218 316226
rect 277274 316170 277342 316226
rect 277398 316170 277494 316226
rect 276874 316102 277494 316170
rect 276874 316046 276970 316102
rect 277026 316046 277094 316102
rect 277150 316046 277218 316102
rect 277274 316046 277342 316102
rect 277398 316046 277494 316102
rect 276874 315978 277494 316046
rect 276874 315922 276970 315978
rect 277026 315922 277094 315978
rect 277150 315922 277218 315978
rect 277274 315922 277342 315978
rect 277398 315922 277494 315978
rect 276874 298422 277494 315922
rect 276874 298366 276970 298422
rect 277026 298366 277094 298422
rect 277150 298366 277218 298422
rect 277274 298366 277342 298422
rect 277398 298366 277494 298422
rect 276874 298342 277494 298366
rect 294874 316350 295494 318858
rect 294874 316294 294970 316350
rect 295026 316294 295094 316350
rect 295150 316294 295218 316350
rect 295274 316294 295342 316350
rect 295398 316294 295494 316350
rect 294874 316226 295494 316294
rect 294874 316170 294970 316226
rect 295026 316170 295094 316226
rect 295150 316170 295218 316226
rect 295274 316170 295342 316226
rect 295398 316170 295494 316226
rect 294874 316102 295494 316170
rect 294874 316046 294970 316102
rect 295026 316046 295094 316102
rect 295150 316046 295218 316102
rect 295274 316046 295342 316102
rect 295398 316046 295494 316102
rect 294874 315978 295494 316046
rect 294874 315922 294970 315978
rect 295026 315922 295094 315978
rect 295150 315922 295218 315978
rect 295274 315922 295342 315978
rect 295398 315922 295494 315978
rect 294874 298422 295494 315922
rect 294874 298366 294970 298422
rect 295026 298366 295094 298422
rect 295150 298366 295218 298422
rect 295274 298366 295342 298422
rect 295398 298366 295494 298422
rect 294874 298342 295494 298366
rect 312874 316350 313494 318858
rect 312874 316294 312970 316350
rect 313026 316294 313094 316350
rect 313150 316294 313218 316350
rect 313274 316294 313342 316350
rect 313398 316294 313494 316350
rect 312874 316226 313494 316294
rect 312874 316170 312970 316226
rect 313026 316170 313094 316226
rect 313150 316170 313218 316226
rect 313274 316170 313342 316226
rect 313398 316170 313494 316226
rect 312874 316102 313494 316170
rect 312874 316046 312970 316102
rect 313026 316046 313094 316102
rect 313150 316046 313218 316102
rect 313274 316046 313342 316102
rect 313398 316046 313494 316102
rect 312874 315978 313494 316046
rect 312874 315922 312970 315978
rect 313026 315922 313094 315978
rect 313150 315922 313218 315978
rect 313274 315922 313342 315978
rect 313398 315922 313494 315978
rect 312874 298422 313494 315922
rect 312874 298366 312970 298422
rect 313026 298366 313094 298422
rect 313150 298366 313218 298422
rect 313274 298366 313342 298422
rect 313398 298366 313494 298422
rect 312874 298342 313494 298366
rect 330874 316350 331494 318858
rect 330874 316294 330970 316350
rect 331026 316294 331094 316350
rect 331150 316294 331218 316350
rect 331274 316294 331342 316350
rect 331398 316294 331494 316350
rect 330874 316226 331494 316294
rect 330874 316170 330970 316226
rect 331026 316170 331094 316226
rect 331150 316170 331218 316226
rect 331274 316170 331342 316226
rect 331398 316170 331494 316226
rect 330874 316102 331494 316170
rect 330874 316046 330970 316102
rect 331026 316046 331094 316102
rect 331150 316046 331218 316102
rect 331274 316046 331342 316102
rect 331398 316046 331494 316102
rect 330874 315978 331494 316046
rect 330874 315922 330970 315978
rect 331026 315922 331094 315978
rect 331150 315922 331218 315978
rect 331274 315922 331342 315978
rect 331398 315922 331494 315978
rect 330874 298422 331494 315922
rect 330874 298366 330970 298422
rect 331026 298366 331094 298422
rect 331150 298366 331218 298422
rect 331274 298366 331342 298422
rect 331398 298366 331494 298422
rect 330874 298342 331494 298366
rect 348874 316350 349494 318858
rect 348874 316294 348970 316350
rect 349026 316294 349094 316350
rect 349150 316294 349218 316350
rect 349274 316294 349342 316350
rect 349398 316294 349494 316350
rect 348874 316226 349494 316294
rect 348874 316170 348970 316226
rect 349026 316170 349094 316226
rect 349150 316170 349218 316226
rect 349274 316170 349342 316226
rect 349398 316170 349494 316226
rect 348874 316102 349494 316170
rect 348874 316046 348970 316102
rect 349026 316046 349094 316102
rect 349150 316046 349218 316102
rect 349274 316046 349342 316102
rect 349398 316046 349494 316102
rect 348874 315978 349494 316046
rect 348874 315922 348970 315978
rect 349026 315922 349094 315978
rect 349150 315922 349218 315978
rect 349274 315922 349342 315978
rect 349398 315922 349494 315978
rect 348874 298422 349494 315922
rect 348874 298366 348970 298422
rect 349026 298366 349094 298422
rect 349150 298366 349218 298422
rect 349274 298366 349342 298422
rect 349398 298366 349494 298422
rect 348874 298342 349494 298366
rect 366874 316350 367494 318858
rect 366874 316294 366970 316350
rect 367026 316294 367094 316350
rect 367150 316294 367218 316350
rect 367274 316294 367342 316350
rect 367398 316294 367494 316350
rect 366874 316226 367494 316294
rect 366874 316170 366970 316226
rect 367026 316170 367094 316226
rect 367150 316170 367218 316226
rect 367274 316170 367342 316226
rect 367398 316170 367494 316226
rect 366874 316102 367494 316170
rect 366874 316046 366970 316102
rect 367026 316046 367094 316102
rect 367150 316046 367218 316102
rect 367274 316046 367342 316102
rect 367398 316046 367494 316102
rect 366874 315978 367494 316046
rect 366874 315922 366970 315978
rect 367026 315922 367094 315978
rect 367150 315922 367218 315978
rect 367274 315922 367342 315978
rect 367398 315922 367494 315978
rect 366874 298422 367494 315922
rect 381154 310350 381774 327922
rect 381154 310294 381250 310350
rect 381306 310294 381374 310350
rect 381430 310294 381498 310350
rect 381554 310294 381622 310350
rect 381678 310294 381774 310350
rect 381154 310226 381774 310294
rect 381154 310170 381250 310226
rect 381306 310170 381374 310226
rect 381430 310170 381498 310226
rect 381554 310170 381622 310226
rect 381678 310170 381774 310226
rect 381154 310102 381774 310170
rect 381154 310046 381250 310102
rect 381306 310046 381374 310102
rect 381430 310046 381498 310102
rect 381554 310046 381622 310102
rect 381678 310046 381774 310102
rect 366874 298366 366970 298422
rect 367026 298366 367094 298422
rect 367150 298366 367218 298422
rect 367274 298366 367342 298422
rect 367398 298366 367494 298422
rect 366874 298342 367494 298366
rect 376348 309988 376404 309998
rect 204874 298226 205494 298294
rect 204874 298170 204970 298226
rect 205026 298170 205094 298226
rect 205150 298170 205218 298226
rect 205274 298170 205342 298226
rect 205398 298170 205494 298226
rect 204874 298102 205494 298170
rect 204874 298046 204970 298102
rect 205026 298046 205094 298102
rect 205150 298046 205218 298102
rect 205274 298046 205342 298102
rect 205398 298046 205494 298102
rect 204874 297978 205494 298046
rect 204874 297922 204970 297978
rect 205026 297922 205094 297978
rect 205150 297922 205218 297978
rect 205274 297922 205342 297978
rect 205398 297922 205494 297978
rect 204874 280350 205494 297922
rect 204874 280294 204970 280350
rect 205026 280294 205094 280350
rect 205150 280294 205218 280350
rect 205274 280294 205342 280350
rect 205398 280294 205494 280350
rect 204874 280226 205494 280294
rect 204874 280170 204970 280226
rect 205026 280170 205094 280226
rect 205150 280170 205218 280226
rect 205274 280170 205342 280226
rect 205398 280170 205494 280226
rect 204874 280102 205494 280170
rect 204874 280046 204970 280102
rect 205026 280046 205094 280102
rect 205150 280046 205218 280102
rect 205274 280046 205342 280102
rect 205398 280046 205494 280102
rect 204874 279978 205494 280046
rect 204874 279922 204970 279978
rect 205026 279922 205094 279978
rect 205150 279922 205218 279978
rect 205274 279922 205342 279978
rect 205398 279922 205494 279978
rect 204874 262350 205494 279922
rect 204874 262294 204970 262350
rect 205026 262294 205094 262350
rect 205150 262294 205218 262350
rect 205274 262294 205342 262350
rect 205398 262294 205494 262350
rect 204874 262226 205494 262294
rect 204874 262170 204970 262226
rect 205026 262170 205094 262226
rect 205150 262170 205218 262226
rect 205274 262170 205342 262226
rect 205398 262170 205494 262226
rect 204874 262102 205494 262170
rect 204874 262046 204970 262102
rect 205026 262046 205094 262102
rect 205150 262046 205218 262102
rect 205274 262046 205342 262102
rect 205398 262046 205494 262102
rect 204874 261978 205494 262046
rect 204874 261922 204970 261978
rect 205026 261922 205094 261978
rect 205150 261922 205218 261978
rect 205274 261922 205342 261978
rect 205398 261922 205494 261978
rect 204874 244350 205494 261922
rect 204874 244294 204970 244350
rect 205026 244294 205094 244350
rect 205150 244294 205218 244350
rect 205274 244294 205342 244350
rect 205398 244294 205494 244350
rect 204874 244226 205494 244294
rect 204874 244170 204970 244226
rect 205026 244170 205094 244226
rect 205150 244170 205218 244226
rect 205274 244170 205342 244226
rect 205398 244170 205494 244226
rect 204874 244102 205494 244170
rect 204874 244046 204970 244102
rect 205026 244046 205094 244102
rect 205150 244046 205218 244102
rect 205274 244046 205342 244102
rect 205398 244046 205494 244102
rect 204874 243978 205494 244046
rect 204874 243922 204970 243978
rect 205026 243922 205094 243978
rect 205150 243922 205218 243978
rect 205274 243922 205342 243978
rect 205398 243922 205494 243978
rect 204874 226350 205494 243922
rect 204874 226294 204970 226350
rect 205026 226294 205094 226350
rect 205150 226294 205218 226350
rect 205274 226294 205342 226350
rect 205398 226294 205494 226350
rect 204874 226226 205494 226294
rect 204874 226170 204970 226226
rect 205026 226170 205094 226226
rect 205150 226170 205218 226226
rect 205274 226170 205342 226226
rect 205398 226170 205494 226226
rect 204874 226102 205494 226170
rect 204874 226046 204970 226102
rect 205026 226046 205094 226102
rect 205150 226046 205218 226102
rect 205274 226046 205342 226102
rect 205398 226046 205494 226102
rect 204874 225978 205494 226046
rect 204874 225922 204970 225978
rect 205026 225922 205094 225978
rect 205150 225922 205218 225978
rect 205274 225922 205342 225978
rect 205398 225922 205494 225978
rect 204874 208350 205494 225922
rect 204874 208294 204970 208350
rect 205026 208294 205094 208350
rect 205150 208294 205218 208350
rect 205274 208294 205342 208350
rect 205398 208294 205494 208350
rect 204874 208226 205494 208294
rect 204874 208170 204970 208226
rect 205026 208170 205094 208226
rect 205150 208170 205218 208226
rect 205274 208170 205342 208226
rect 205398 208170 205494 208226
rect 204874 208102 205494 208170
rect 204874 208046 204970 208102
rect 205026 208046 205094 208102
rect 205150 208046 205218 208102
rect 205274 208046 205342 208102
rect 205398 208046 205494 208102
rect 204874 207978 205494 208046
rect 204874 207922 204970 207978
rect 205026 207922 205094 207978
rect 205150 207922 205218 207978
rect 205274 207922 205342 207978
rect 205398 207922 205494 207978
rect 204874 190350 205494 207922
rect 204874 190294 204970 190350
rect 205026 190294 205094 190350
rect 205150 190294 205218 190350
rect 205274 190294 205342 190350
rect 205398 190294 205494 190350
rect 204874 190226 205494 190294
rect 204874 190170 204970 190226
rect 205026 190170 205094 190226
rect 205150 190170 205218 190226
rect 205274 190170 205342 190226
rect 205398 190170 205494 190226
rect 204874 190102 205494 190170
rect 204874 190046 204970 190102
rect 205026 190046 205094 190102
rect 205150 190046 205218 190102
rect 205274 190046 205342 190102
rect 205398 190046 205494 190102
rect 204874 189978 205494 190046
rect 204874 189922 204970 189978
rect 205026 189922 205094 189978
rect 205150 189922 205218 189978
rect 205274 189922 205342 189978
rect 205398 189922 205494 189978
rect 204874 172350 205494 189922
rect 204874 172294 204970 172350
rect 205026 172294 205094 172350
rect 205150 172294 205218 172350
rect 205274 172294 205342 172350
rect 205398 172294 205494 172350
rect 204874 172226 205494 172294
rect 204874 172170 204970 172226
rect 205026 172170 205094 172226
rect 205150 172170 205218 172226
rect 205274 172170 205342 172226
rect 205398 172170 205494 172226
rect 204874 172102 205494 172170
rect 204874 172046 204970 172102
rect 205026 172046 205094 172102
rect 205150 172046 205218 172102
rect 205274 172046 205342 172102
rect 205398 172046 205494 172102
rect 204874 171978 205494 172046
rect 204874 171922 204970 171978
rect 205026 171922 205094 171978
rect 205150 171922 205218 171978
rect 205274 171922 205342 171978
rect 205398 171922 205494 171978
rect 204874 154350 205494 171922
rect 204874 154294 204970 154350
rect 205026 154294 205094 154350
rect 205150 154294 205218 154350
rect 205274 154294 205342 154350
rect 205398 154294 205494 154350
rect 204874 154226 205494 154294
rect 204874 154170 204970 154226
rect 205026 154170 205094 154226
rect 205150 154170 205218 154226
rect 205274 154170 205342 154226
rect 205398 154170 205494 154226
rect 204874 154102 205494 154170
rect 204874 154046 204970 154102
rect 205026 154046 205094 154102
rect 205150 154046 205218 154102
rect 205274 154046 205342 154102
rect 205398 154046 205494 154102
rect 204874 153978 205494 154046
rect 211708 156884 211764 156894
rect 204874 153922 204970 153978
rect 205026 153922 205094 153978
rect 205150 153922 205218 153978
rect 205274 153922 205342 153978
rect 205398 153922 205494 153978
rect 204874 136350 205494 153922
rect 205660 153972 205716 153982
rect 205660 152852 205716 153916
rect 211708 153972 211764 156828
rect 211708 153906 211764 153916
rect 205660 152786 205716 152796
rect 219154 148422 219774 158858
rect 219154 148366 219250 148422
rect 219306 148366 219374 148422
rect 219430 148366 219498 148422
rect 219554 148366 219622 148422
rect 219678 148366 219774 148422
rect 219154 148342 219774 148366
rect 222874 154350 223494 158858
rect 222874 154294 222970 154350
rect 223026 154294 223094 154350
rect 223150 154294 223218 154350
rect 223274 154294 223342 154350
rect 223398 154294 223494 154350
rect 222874 154226 223494 154294
rect 222874 154170 222970 154226
rect 223026 154170 223094 154226
rect 223150 154170 223218 154226
rect 223274 154170 223342 154226
rect 223398 154170 223494 154226
rect 222874 154102 223494 154170
rect 222874 154046 222970 154102
rect 223026 154046 223094 154102
rect 223150 154046 223218 154102
rect 223274 154046 223342 154102
rect 223398 154046 223494 154102
rect 222874 153978 223494 154046
rect 222874 153922 222970 153978
rect 223026 153922 223094 153978
rect 223150 153922 223218 153978
rect 223274 153922 223342 153978
rect 223398 153922 223494 153978
rect 222874 148342 223494 153922
rect 237154 148422 237774 158858
rect 237154 148366 237250 148422
rect 237306 148366 237374 148422
rect 237430 148366 237498 148422
rect 237554 148366 237622 148422
rect 237678 148366 237774 148422
rect 237154 148342 237774 148366
rect 240874 154350 241494 158858
rect 240874 154294 240970 154350
rect 241026 154294 241094 154350
rect 241150 154294 241218 154350
rect 241274 154294 241342 154350
rect 241398 154294 241494 154350
rect 240874 154226 241494 154294
rect 240874 154170 240970 154226
rect 241026 154170 241094 154226
rect 241150 154170 241218 154226
rect 241274 154170 241342 154226
rect 241398 154170 241494 154226
rect 240874 154102 241494 154170
rect 240874 154046 240970 154102
rect 241026 154046 241094 154102
rect 241150 154046 241218 154102
rect 241274 154046 241342 154102
rect 241398 154046 241494 154102
rect 240874 153978 241494 154046
rect 240874 153922 240970 153978
rect 241026 153922 241094 153978
rect 241150 153922 241218 153978
rect 241274 153922 241342 153978
rect 241398 153922 241494 153978
rect 240874 148342 241494 153922
rect 255154 148422 255774 158858
rect 255154 148366 255250 148422
rect 255306 148366 255374 148422
rect 255430 148366 255498 148422
rect 255554 148366 255622 148422
rect 255678 148366 255774 148422
rect 255154 148342 255774 148366
rect 258874 154350 259494 158858
rect 258874 154294 258970 154350
rect 259026 154294 259094 154350
rect 259150 154294 259218 154350
rect 259274 154294 259342 154350
rect 259398 154294 259494 154350
rect 258874 154226 259494 154294
rect 258874 154170 258970 154226
rect 259026 154170 259094 154226
rect 259150 154170 259218 154226
rect 259274 154170 259342 154226
rect 259398 154170 259494 154226
rect 258874 154102 259494 154170
rect 258874 154046 258970 154102
rect 259026 154046 259094 154102
rect 259150 154046 259218 154102
rect 259274 154046 259342 154102
rect 259398 154046 259494 154102
rect 258874 153978 259494 154046
rect 258874 153922 258970 153978
rect 259026 153922 259094 153978
rect 259150 153922 259218 153978
rect 259274 153922 259342 153978
rect 259398 153922 259494 153978
rect 258874 148342 259494 153922
rect 273154 148422 273774 158858
rect 273154 148366 273250 148422
rect 273306 148366 273374 148422
rect 273430 148366 273498 148422
rect 273554 148366 273622 148422
rect 273678 148366 273774 148422
rect 273154 148342 273774 148366
rect 276874 154350 277494 158858
rect 276874 154294 276970 154350
rect 277026 154294 277094 154350
rect 277150 154294 277218 154350
rect 277274 154294 277342 154350
rect 277398 154294 277494 154350
rect 276874 154226 277494 154294
rect 276874 154170 276970 154226
rect 277026 154170 277094 154226
rect 277150 154170 277218 154226
rect 277274 154170 277342 154226
rect 277398 154170 277494 154226
rect 276874 154102 277494 154170
rect 276874 154046 276970 154102
rect 277026 154046 277094 154102
rect 277150 154046 277218 154102
rect 277274 154046 277342 154102
rect 277398 154046 277494 154102
rect 276874 153978 277494 154046
rect 276874 153922 276970 153978
rect 277026 153922 277094 153978
rect 277150 153922 277218 153978
rect 277274 153922 277342 153978
rect 277398 153922 277494 153978
rect 276874 148342 277494 153922
rect 291154 148422 291774 158858
rect 291154 148366 291250 148422
rect 291306 148366 291374 148422
rect 291430 148366 291498 148422
rect 291554 148366 291622 148422
rect 291678 148366 291774 148422
rect 291154 148342 291774 148366
rect 294874 154350 295494 158858
rect 294874 154294 294970 154350
rect 295026 154294 295094 154350
rect 295150 154294 295218 154350
rect 295274 154294 295342 154350
rect 295398 154294 295494 154350
rect 294874 154226 295494 154294
rect 294874 154170 294970 154226
rect 295026 154170 295094 154226
rect 295150 154170 295218 154226
rect 295274 154170 295342 154226
rect 295398 154170 295494 154226
rect 294874 154102 295494 154170
rect 294874 154046 294970 154102
rect 295026 154046 295094 154102
rect 295150 154046 295218 154102
rect 295274 154046 295342 154102
rect 295398 154046 295494 154102
rect 294874 153978 295494 154046
rect 294874 153922 294970 153978
rect 295026 153922 295094 153978
rect 295150 153922 295218 153978
rect 295274 153922 295342 153978
rect 295398 153922 295494 153978
rect 294874 148342 295494 153922
rect 309154 148422 309774 158858
rect 309154 148366 309250 148422
rect 309306 148366 309374 148422
rect 309430 148366 309498 148422
rect 309554 148366 309622 148422
rect 309678 148366 309774 148422
rect 309154 148342 309774 148366
rect 312874 154350 313494 158858
rect 312874 154294 312970 154350
rect 313026 154294 313094 154350
rect 313150 154294 313218 154350
rect 313274 154294 313342 154350
rect 313398 154294 313494 154350
rect 312874 154226 313494 154294
rect 312874 154170 312970 154226
rect 313026 154170 313094 154226
rect 313150 154170 313218 154226
rect 313274 154170 313342 154226
rect 313398 154170 313494 154226
rect 312874 154102 313494 154170
rect 312874 154046 312970 154102
rect 313026 154046 313094 154102
rect 313150 154046 313218 154102
rect 313274 154046 313342 154102
rect 313398 154046 313494 154102
rect 312874 153978 313494 154046
rect 312874 153922 312970 153978
rect 313026 153922 313094 153978
rect 313150 153922 313218 153978
rect 313274 153922 313342 153978
rect 313398 153922 313494 153978
rect 312874 148342 313494 153922
rect 327154 148422 327774 158858
rect 327154 148366 327250 148422
rect 327306 148366 327374 148422
rect 327430 148366 327498 148422
rect 327554 148366 327622 148422
rect 327678 148366 327774 148422
rect 327154 148342 327774 148366
rect 330874 154350 331494 158858
rect 330874 154294 330970 154350
rect 331026 154294 331094 154350
rect 331150 154294 331218 154350
rect 331274 154294 331342 154350
rect 331398 154294 331494 154350
rect 330874 154226 331494 154294
rect 330874 154170 330970 154226
rect 331026 154170 331094 154226
rect 331150 154170 331218 154226
rect 331274 154170 331342 154226
rect 331398 154170 331494 154226
rect 330874 154102 331494 154170
rect 330874 154046 330970 154102
rect 331026 154046 331094 154102
rect 331150 154046 331218 154102
rect 331274 154046 331342 154102
rect 331398 154046 331494 154102
rect 330874 153978 331494 154046
rect 330874 153922 330970 153978
rect 331026 153922 331094 153978
rect 331150 153922 331218 153978
rect 331274 153922 331342 153978
rect 331398 153922 331494 153978
rect 330874 148342 331494 153922
rect 345154 148422 345774 158858
rect 345154 148366 345250 148422
rect 345306 148366 345374 148422
rect 345430 148366 345498 148422
rect 345554 148366 345622 148422
rect 345678 148366 345774 148422
rect 345154 148342 345774 148366
rect 348874 154350 349494 158858
rect 348874 154294 348970 154350
rect 349026 154294 349094 154350
rect 349150 154294 349218 154350
rect 349274 154294 349342 154350
rect 349398 154294 349494 154350
rect 348874 154226 349494 154294
rect 348874 154170 348970 154226
rect 349026 154170 349094 154226
rect 349150 154170 349218 154226
rect 349274 154170 349342 154226
rect 349398 154170 349494 154226
rect 348874 154102 349494 154170
rect 348874 154046 348970 154102
rect 349026 154046 349094 154102
rect 349150 154046 349218 154102
rect 349274 154046 349342 154102
rect 349398 154046 349494 154102
rect 348874 153978 349494 154046
rect 348874 153922 348970 153978
rect 349026 153922 349094 153978
rect 349150 153922 349218 153978
rect 349274 153922 349342 153978
rect 349398 153922 349494 153978
rect 348874 148342 349494 153922
rect 363154 148422 363774 158858
rect 363154 148366 363250 148422
rect 363306 148366 363374 148422
rect 363430 148366 363498 148422
rect 363554 148366 363622 148422
rect 363678 148366 363774 148422
rect 363154 148342 363774 148366
rect 366874 154350 367494 158858
rect 366874 154294 366970 154350
rect 367026 154294 367094 154350
rect 367150 154294 367218 154350
rect 367274 154294 367342 154350
rect 367398 154294 367494 154350
rect 366874 154226 367494 154294
rect 366874 154170 366970 154226
rect 367026 154170 367094 154226
rect 367150 154170 367218 154226
rect 367274 154170 367342 154226
rect 367398 154170 367494 154226
rect 366874 154102 367494 154170
rect 366874 154046 366970 154102
rect 367026 154046 367094 154102
rect 367150 154046 367218 154102
rect 367274 154046 367342 154102
rect 367398 154046 367494 154102
rect 366874 153978 367494 154046
rect 366874 153922 366970 153978
rect 367026 153922 367094 153978
rect 367150 153922 367218 153978
rect 367274 153922 367342 153978
rect 367398 153922 367494 153978
rect 366874 148342 367494 153922
rect 376348 156324 376404 309932
rect 381154 309978 381774 310046
rect 381154 309922 381250 309978
rect 381306 309922 381374 309978
rect 381430 309922 381498 309978
rect 381554 309922 381622 309978
rect 381678 309922 381774 309978
rect 381154 292350 381774 309922
rect 381154 292294 381250 292350
rect 381306 292294 381374 292350
rect 381430 292294 381498 292350
rect 381554 292294 381622 292350
rect 381678 292294 381774 292350
rect 381154 292226 381774 292294
rect 381154 292170 381250 292226
rect 381306 292170 381374 292226
rect 381430 292170 381498 292226
rect 381554 292170 381622 292226
rect 381678 292170 381774 292226
rect 381154 292102 381774 292170
rect 381154 292046 381250 292102
rect 381306 292046 381374 292102
rect 381430 292046 381498 292102
rect 381554 292046 381622 292102
rect 381678 292046 381774 292102
rect 381154 291978 381774 292046
rect 381154 291922 381250 291978
rect 381306 291922 381374 291978
rect 381430 291922 381498 291978
rect 381554 291922 381622 291978
rect 381678 291922 381774 291978
rect 381154 274350 381774 291922
rect 381154 274294 381250 274350
rect 381306 274294 381374 274350
rect 381430 274294 381498 274350
rect 381554 274294 381622 274350
rect 381678 274294 381774 274350
rect 381154 274226 381774 274294
rect 381154 274170 381250 274226
rect 381306 274170 381374 274226
rect 381430 274170 381498 274226
rect 381554 274170 381622 274226
rect 381678 274170 381774 274226
rect 381154 274102 381774 274170
rect 381154 274046 381250 274102
rect 381306 274046 381374 274102
rect 381430 274046 381498 274102
rect 381554 274046 381622 274102
rect 381678 274046 381774 274102
rect 381154 273978 381774 274046
rect 381154 273922 381250 273978
rect 381306 273922 381374 273978
rect 381430 273922 381498 273978
rect 381554 273922 381622 273978
rect 381678 273922 381774 273978
rect 381154 256350 381774 273922
rect 381154 256294 381250 256350
rect 381306 256294 381374 256350
rect 381430 256294 381498 256350
rect 381554 256294 381622 256350
rect 381678 256294 381774 256350
rect 381154 256226 381774 256294
rect 381154 256170 381250 256226
rect 381306 256170 381374 256226
rect 381430 256170 381498 256226
rect 381554 256170 381622 256226
rect 381678 256170 381774 256226
rect 381154 256102 381774 256170
rect 381154 256046 381250 256102
rect 381306 256046 381374 256102
rect 381430 256046 381498 256102
rect 381554 256046 381622 256102
rect 381678 256046 381774 256102
rect 381154 255978 381774 256046
rect 381154 255922 381250 255978
rect 381306 255922 381374 255978
rect 381430 255922 381498 255978
rect 381554 255922 381622 255978
rect 381678 255922 381774 255978
rect 381154 238350 381774 255922
rect 381154 238294 381250 238350
rect 381306 238294 381374 238350
rect 381430 238294 381498 238350
rect 381554 238294 381622 238350
rect 381678 238294 381774 238350
rect 381154 238226 381774 238294
rect 381154 238170 381250 238226
rect 381306 238170 381374 238226
rect 381430 238170 381498 238226
rect 381554 238170 381622 238226
rect 381678 238170 381774 238226
rect 381154 238102 381774 238170
rect 381154 238046 381250 238102
rect 381306 238046 381374 238102
rect 381430 238046 381498 238102
rect 381554 238046 381622 238102
rect 381678 238046 381774 238102
rect 381154 237978 381774 238046
rect 381154 237922 381250 237978
rect 381306 237922 381374 237978
rect 381430 237922 381498 237978
rect 381554 237922 381622 237978
rect 381678 237922 381774 237978
rect 381154 220350 381774 237922
rect 381154 220294 381250 220350
rect 381306 220294 381374 220350
rect 381430 220294 381498 220350
rect 381554 220294 381622 220350
rect 381678 220294 381774 220350
rect 381154 220226 381774 220294
rect 381154 220170 381250 220226
rect 381306 220170 381374 220226
rect 381430 220170 381498 220226
rect 381554 220170 381622 220226
rect 381678 220170 381774 220226
rect 381154 220102 381774 220170
rect 381154 220046 381250 220102
rect 381306 220046 381374 220102
rect 381430 220046 381498 220102
rect 381554 220046 381622 220102
rect 381678 220046 381774 220102
rect 381154 219978 381774 220046
rect 381154 219922 381250 219978
rect 381306 219922 381374 219978
rect 381430 219922 381498 219978
rect 381554 219922 381622 219978
rect 381678 219922 381774 219978
rect 381154 202350 381774 219922
rect 381154 202294 381250 202350
rect 381306 202294 381374 202350
rect 381430 202294 381498 202350
rect 381554 202294 381622 202350
rect 381678 202294 381774 202350
rect 381154 202226 381774 202294
rect 381154 202170 381250 202226
rect 381306 202170 381374 202226
rect 381430 202170 381498 202226
rect 381554 202170 381622 202226
rect 381678 202170 381774 202226
rect 381154 202102 381774 202170
rect 381154 202046 381250 202102
rect 381306 202046 381374 202102
rect 381430 202046 381498 202102
rect 381554 202046 381622 202102
rect 381678 202046 381774 202102
rect 381154 201978 381774 202046
rect 381154 201922 381250 201978
rect 381306 201922 381374 201978
rect 381430 201922 381498 201978
rect 381554 201922 381622 201978
rect 381678 201922 381774 201978
rect 381154 184350 381774 201922
rect 381154 184294 381250 184350
rect 381306 184294 381374 184350
rect 381430 184294 381498 184350
rect 381554 184294 381622 184350
rect 381678 184294 381774 184350
rect 381154 184226 381774 184294
rect 381154 184170 381250 184226
rect 381306 184170 381374 184226
rect 381430 184170 381498 184226
rect 381554 184170 381622 184226
rect 381678 184170 381774 184226
rect 381154 184102 381774 184170
rect 381154 184046 381250 184102
rect 381306 184046 381374 184102
rect 381430 184046 381498 184102
rect 381554 184046 381622 184102
rect 381678 184046 381774 184102
rect 381154 183978 381774 184046
rect 381154 183922 381250 183978
rect 381306 183922 381374 183978
rect 381430 183922 381498 183978
rect 381554 183922 381622 183978
rect 381678 183922 381774 183978
rect 381154 166350 381774 183922
rect 381154 166294 381250 166350
rect 381306 166294 381374 166350
rect 381430 166294 381498 166350
rect 381554 166294 381622 166350
rect 381678 166294 381774 166350
rect 381154 166226 381774 166294
rect 381154 166170 381250 166226
rect 381306 166170 381374 166226
rect 381430 166170 381498 166226
rect 381554 166170 381622 166226
rect 381678 166170 381774 166226
rect 381154 166102 381774 166170
rect 381154 166046 381250 166102
rect 381306 166046 381374 166102
rect 381430 166046 381498 166102
rect 381554 166046 381622 166102
rect 381678 166046 381774 166102
rect 381154 165978 381774 166046
rect 381154 165922 381250 165978
rect 381306 165922 381374 165978
rect 381430 165922 381498 165978
rect 381554 165922 381622 165978
rect 381678 165922 381774 165978
rect 204874 136294 204970 136350
rect 205026 136294 205094 136350
rect 205150 136294 205218 136350
rect 205274 136294 205342 136350
rect 205398 136294 205494 136350
rect 204874 136226 205494 136294
rect 204874 136170 204970 136226
rect 205026 136170 205094 136226
rect 205150 136170 205218 136226
rect 205274 136170 205342 136226
rect 205398 136170 205494 136226
rect 204874 136102 205494 136170
rect 204874 136046 204970 136102
rect 205026 136046 205094 136102
rect 205150 136046 205218 136102
rect 205274 136046 205342 136102
rect 205398 136046 205494 136102
rect 204874 135978 205494 136046
rect 204874 135922 204970 135978
rect 205026 135922 205094 135978
rect 205150 135922 205218 135978
rect 205274 135922 205342 135978
rect 205398 135922 205494 135978
rect 204874 118350 205494 135922
rect 204874 118294 204970 118350
rect 205026 118294 205094 118350
rect 205150 118294 205218 118350
rect 205274 118294 205342 118350
rect 205398 118294 205494 118350
rect 204874 118226 205494 118294
rect 204874 118170 204970 118226
rect 205026 118170 205094 118226
rect 205150 118170 205218 118226
rect 205274 118170 205342 118226
rect 205398 118170 205494 118226
rect 204874 118102 205494 118170
rect 204874 118046 204970 118102
rect 205026 118046 205094 118102
rect 205150 118046 205218 118102
rect 205274 118046 205342 118102
rect 205398 118046 205494 118102
rect 204874 117978 205494 118046
rect 204874 117922 204970 117978
rect 205026 117922 205094 117978
rect 205150 117922 205218 117978
rect 205274 117922 205342 117978
rect 205398 117922 205494 117978
rect 204874 100350 205494 117922
rect 204874 100294 204970 100350
rect 205026 100294 205094 100350
rect 205150 100294 205218 100350
rect 205274 100294 205342 100350
rect 205398 100294 205494 100350
rect 204874 100226 205494 100294
rect 204874 100170 204970 100226
rect 205026 100170 205094 100226
rect 205150 100170 205218 100226
rect 205274 100170 205342 100226
rect 205398 100170 205494 100226
rect 204874 100102 205494 100170
rect 204874 100046 204970 100102
rect 205026 100046 205094 100102
rect 205150 100046 205218 100102
rect 205274 100046 205342 100102
rect 205398 100046 205494 100102
rect 204874 99978 205494 100046
rect 204874 99922 204970 99978
rect 205026 99922 205094 99978
rect 205150 99922 205218 99978
rect 205274 99922 205342 99978
rect 205398 99922 205494 99978
rect 204874 82350 205494 99922
rect 204874 82294 204970 82350
rect 205026 82294 205094 82350
rect 205150 82294 205218 82350
rect 205274 82294 205342 82350
rect 205398 82294 205494 82350
rect 204874 82226 205494 82294
rect 204874 82170 204970 82226
rect 205026 82170 205094 82226
rect 205150 82170 205218 82226
rect 205274 82170 205342 82226
rect 205398 82170 205494 82226
rect 204874 82102 205494 82170
rect 204874 82046 204970 82102
rect 205026 82046 205094 82102
rect 205150 82046 205218 82102
rect 205274 82046 205342 82102
rect 205398 82046 205494 82102
rect 204874 81978 205494 82046
rect 204874 81922 204970 81978
rect 205026 81922 205094 81978
rect 205150 81922 205218 81978
rect 205274 81922 205342 81978
rect 205398 81922 205494 81978
rect 204874 64350 205494 81922
rect 204874 64294 204970 64350
rect 205026 64294 205094 64350
rect 205150 64294 205218 64350
rect 205274 64294 205342 64350
rect 205398 64294 205494 64350
rect 204874 64226 205494 64294
rect 204874 64170 204970 64226
rect 205026 64170 205094 64226
rect 205150 64170 205218 64226
rect 205274 64170 205342 64226
rect 205398 64170 205494 64226
rect 204874 64102 205494 64170
rect 204874 64046 204970 64102
rect 205026 64046 205094 64102
rect 205150 64046 205218 64102
rect 205274 64046 205342 64102
rect 205398 64046 205494 64102
rect 204874 63978 205494 64046
rect 204874 63922 204970 63978
rect 205026 63922 205094 63978
rect 205150 63922 205218 63978
rect 205274 63922 205342 63978
rect 205398 63922 205494 63978
rect 204874 46350 205494 63922
rect 204874 46294 204970 46350
rect 205026 46294 205094 46350
rect 205150 46294 205218 46350
rect 205274 46294 205342 46350
rect 205398 46294 205494 46350
rect 204874 46226 205494 46294
rect 204874 46170 204970 46226
rect 205026 46170 205094 46226
rect 205150 46170 205218 46226
rect 205274 46170 205342 46226
rect 205398 46170 205494 46226
rect 204874 46102 205494 46170
rect 204874 46046 204970 46102
rect 205026 46046 205094 46102
rect 205150 46046 205218 46102
rect 205274 46046 205342 46102
rect 205398 46046 205494 46102
rect 204874 45978 205494 46046
rect 204874 45922 204970 45978
rect 205026 45922 205094 45978
rect 205150 45922 205218 45978
rect 205274 45922 205342 45978
rect 205398 45922 205494 45978
rect 204874 28350 205494 45922
rect 204874 28294 204970 28350
rect 205026 28294 205094 28350
rect 205150 28294 205218 28350
rect 205274 28294 205342 28350
rect 205398 28294 205494 28350
rect 204874 28226 205494 28294
rect 204874 28170 204970 28226
rect 205026 28170 205094 28226
rect 205150 28170 205218 28226
rect 205274 28170 205342 28226
rect 205398 28170 205494 28226
rect 204874 28102 205494 28170
rect 204874 28046 204970 28102
rect 205026 28046 205094 28102
rect 205150 28046 205218 28102
rect 205274 28046 205342 28102
rect 205398 28046 205494 28102
rect 204874 27978 205494 28046
rect 204874 27922 204970 27978
rect 205026 27922 205094 27978
rect 205150 27922 205218 27978
rect 205274 27922 205342 27978
rect 205398 27922 205494 27978
rect 204874 10350 205494 27922
rect 204874 10294 204970 10350
rect 205026 10294 205094 10350
rect 205150 10294 205218 10350
rect 205274 10294 205342 10350
rect 205398 10294 205494 10350
rect 204874 10226 205494 10294
rect 204874 10170 204970 10226
rect 205026 10170 205094 10226
rect 205150 10170 205218 10226
rect 205274 10170 205342 10226
rect 205398 10170 205494 10226
rect 204874 10102 205494 10170
rect 204874 10046 204970 10102
rect 205026 10046 205094 10102
rect 205150 10046 205218 10102
rect 205274 10046 205342 10102
rect 205398 10046 205494 10102
rect 204874 9978 205494 10046
rect 204874 9922 204970 9978
rect 205026 9922 205094 9978
rect 205150 9922 205218 9978
rect 205274 9922 205342 9978
rect 205398 9922 205494 9978
rect 204874 -1120 205494 9922
rect 204874 -1176 204970 -1120
rect 205026 -1176 205094 -1120
rect 205150 -1176 205218 -1120
rect 205274 -1176 205342 -1120
rect 205398 -1176 205494 -1120
rect 204874 -1244 205494 -1176
rect 204874 -1300 204970 -1244
rect 205026 -1300 205094 -1244
rect 205150 -1300 205218 -1244
rect 205274 -1300 205342 -1244
rect 205398 -1300 205494 -1244
rect 204874 -1368 205494 -1300
rect 204874 -1424 204970 -1368
rect 205026 -1424 205094 -1368
rect 205150 -1424 205218 -1368
rect 205274 -1424 205342 -1368
rect 205398 -1424 205494 -1368
rect 204874 -1492 205494 -1424
rect 204874 -1548 204970 -1492
rect 205026 -1548 205094 -1492
rect 205150 -1548 205218 -1492
rect 205274 -1548 205342 -1492
rect 205398 -1548 205494 -1492
rect 204874 -1644 205494 -1548
rect 219154 4350 219774 8858
rect 219154 4294 219250 4350
rect 219306 4294 219374 4350
rect 219430 4294 219498 4350
rect 219554 4294 219622 4350
rect 219678 4294 219774 4350
rect 219154 4226 219774 4294
rect 219154 4170 219250 4226
rect 219306 4170 219374 4226
rect 219430 4170 219498 4226
rect 219554 4170 219622 4226
rect 219678 4170 219774 4226
rect 219154 4102 219774 4170
rect 219154 4046 219250 4102
rect 219306 4046 219374 4102
rect 219430 4046 219498 4102
rect 219554 4046 219622 4102
rect 219678 4046 219774 4102
rect 219154 3978 219774 4046
rect 219154 3922 219250 3978
rect 219306 3922 219374 3978
rect 219430 3922 219498 3978
rect 219554 3922 219622 3978
rect 219678 3922 219774 3978
rect 219154 -160 219774 3922
rect 219154 -216 219250 -160
rect 219306 -216 219374 -160
rect 219430 -216 219498 -160
rect 219554 -216 219622 -160
rect 219678 -216 219774 -160
rect 219154 -284 219774 -216
rect 219154 -340 219250 -284
rect 219306 -340 219374 -284
rect 219430 -340 219498 -284
rect 219554 -340 219622 -284
rect 219678 -340 219774 -284
rect 219154 -408 219774 -340
rect 219154 -464 219250 -408
rect 219306 -464 219374 -408
rect 219430 -464 219498 -408
rect 219554 -464 219622 -408
rect 219678 -464 219774 -408
rect 219154 -532 219774 -464
rect 219154 -588 219250 -532
rect 219306 -588 219374 -532
rect 219430 -588 219498 -532
rect 219554 -588 219622 -532
rect 219678 -588 219774 -532
rect 219154 -1644 219774 -588
rect 237154 4350 237774 8858
rect 237154 4294 237250 4350
rect 237306 4294 237374 4350
rect 237430 4294 237498 4350
rect 237554 4294 237622 4350
rect 237678 4294 237774 4350
rect 237154 4226 237774 4294
rect 237154 4170 237250 4226
rect 237306 4170 237374 4226
rect 237430 4170 237498 4226
rect 237554 4170 237622 4226
rect 237678 4170 237774 4226
rect 237154 4102 237774 4170
rect 237154 4046 237250 4102
rect 237306 4046 237374 4102
rect 237430 4046 237498 4102
rect 237554 4046 237622 4102
rect 237678 4046 237774 4102
rect 237154 3978 237774 4046
rect 237154 3922 237250 3978
rect 237306 3922 237374 3978
rect 237430 3922 237498 3978
rect 237554 3922 237622 3978
rect 237678 3922 237774 3978
rect 237154 -160 237774 3922
rect 237154 -216 237250 -160
rect 237306 -216 237374 -160
rect 237430 -216 237498 -160
rect 237554 -216 237622 -160
rect 237678 -216 237774 -160
rect 237154 -284 237774 -216
rect 237154 -340 237250 -284
rect 237306 -340 237374 -284
rect 237430 -340 237498 -284
rect 237554 -340 237622 -284
rect 237678 -340 237774 -284
rect 237154 -408 237774 -340
rect 237154 -464 237250 -408
rect 237306 -464 237374 -408
rect 237430 -464 237498 -408
rect 237554 -464 237622 -408
rect 237678 -464 237774 -408
rect 237154 -532 237774 -464
rect 237154 -588 237250 -532
rect 237306 -588 237374 -532
rect 237430 -588 237498 -532
rect 237554 -588 237622 -532
rect 237678 -588 237774 -532
rect 237154 -1644 237774 -588
rect 255154 4350 255774 8858
rect 255154 4294 255250 4350
rect 255306 4294 255374 4350
rect 255430 4294 255498 4350
rect 255554 4294 255622 4350
rect 255678 4294 255774 4350
rect 255154 4226 255774 4294
rect 255154 4170 255250 4226
rect 255306 4170 255374 4226
rect 255430 4170 255498 4226
rect 255554 4170 255622 4226
rect 255678 4170 255774 4226
rect 255154 4102 255774 4170
rect 255154 4046 255250 4102
rect 255306 4046 255374 4102
rect 255430 4046 255498 4102
rect 255554 4046 255622 4102
rect 255678 4046 255774 4102
rect 255154 3978 255774 4046
rect 255154 3922 255250 3978
rect 255306 3922 255374 3978
rect 255430 3922 255498 3978
rect 255554 3922 255622 3978
rect 255678 3922 255774 3978
rect 255154 -160 255774 3922
rect 255154 -216 255250 -160
rect 255306 -216 255374 -160
rect 255430 -216 255498 -160
rect 255554 -216 255622 -160
rect 255678 -216 255774 -160
rect 255154 -284 255774 -216
rect 255154 -340 255250 -284
rect 255306 -340 255374 -284
rect 255430 -340 255498 -284
rect 255554 -340 255622 -284
rect 255678 -340 255774 -284
rect 255154 -408 255774 -340
rect 255154 -464 255250 -408
rect 255306 -464 255374 -408
rect 255430 -464 255498 -408
rect 255554 -464 255622 -408
rect 255678 -464 255774 -408
rect 255154 -532 255774 -464
rect 255154 -588 255250 -532
rect 255306 -588 255374 -532
rect 255430 -588 255498 -532
rect 255554 -588 255622 -532
rect 255678 -588 255774 -532
rect 255154 -1644 255774 -588
rect 273154 4350 273774 8858
rect 273154 4294 273250 4350
rect 273306 4294 273374 4350
rect 273430 4294 273498 4350
rect 273554 4294 273622 4350
rect 273678 4294 273774 4350
rect 273154 4226 273774 4294
rect 273154 4170 273250 4226
rect 273306 4170 273374 4226
rect 273430 4170 273498 4226
rect 273554 4170 273622 4226
rect 273678 4170 273774 4226
rect 273154 4102 273774 4170
rect 273154 4046 273250 4102
rect 273306 4046 273374 4102
rect 273430 4046 273498 4102
rect 273554 4046 273622 4102
rect 273678 4046 273774 4102
rect 273154 3978 273774 4046
rect 273154 3922 273250 3978
rect 273306 3922 273374 3978
rect 273430 3922 273498 3978
rect 273554 3922 273622 3978
rect 273678 3922 273774 3978
rect 273154 -160 273774 3922
rect 273154 -216 273250 -160
rect 273306 -216 273374 -160
rect 273430 -216 273498 -160
rect 273554 -216 273622 -160
rect 273678 -216 273774 -160
rect 273154 -284 273774 -216
rect 273154 -340 273250 -284
rect 273306 -340 273374 -284
rect 273430 -340 273498 -284
rect 273554 -340 273622 -284
rect 273678 -340 273774 -284
rect 273154 -408 273774 -340
rect 273154 -464 273250 -408
rect 273306 -464 273374 -408
rect 273430 -464 273498 -408
rect 273554 -464 273622 -408
rect 273678 -464 273774 -408
rect 273154 -532 273774 -464
rect 273154 -588 273250 -532
rect 273306 -588 273374 -532
rect 273430 -588 273498 -532
rect 273554 -588 273622 -532
rect 273678 -588 273774 -532
rect 273154 -1644 273774 -588
rect 291154 4350 291774 8858
rect 291154 4294 291250 4350
rect 291306 4294 291374 4350
rect 291430 4294 291498 4350
rect 291554 4294 291622 4350
rect 291678 4294 291774 4350
rect 291154 4226 291774 4294
rect 291154 4170 291250 4226
rect 291306 4170 291374 4226
rect 291430 4170 291498 4226
rect 291554 4170 291622 4226
rect 291678 4170 291774 4226
rect 291154 4102 291774 4170
rect 291154 4046 291250 4102
rect 291306 4046 291374 4102
rect 291430 4046 291498 4102
rect 291554 4046 291622 4102
rect 291678 4046 291774 4102
rect 291154 3978 291774 4046
rect 291154 3922 291250 3978
rect 291306 3922 291374 3978
rect 291430 3922 291498 3978
rect 291554 3922 291622 3978
rect 291678 3922 291774 3978
rect 291154 -160 291774 3922
rect 291154 -216 291250 -160
rect 291306 -216 291374 -160
rect 291430 -216 291498 -160
rect 291554 -216 291622 -160
rect 291678 -216 291774 -160
rect 291154 -284 291774 -216
rect 291154 -340 291250 -284
rect 291306 -340 291374 -284
rect 291430 -340 291498 -284
rect 291554 -340 291622 -284
rect 291678 -340 291774 -284
rect 291154 -408 291774 -340
rect 291154 -464 291250 -408
rect 291306 -464 291374 -408
rect 291430 -464 291498 -408
rect 291554 -464 291622 -408
rect 291678 -464 291774 -408
rect 291154 -532 291774 -464
rect 291154 -588 291250 -532
rect 291306 -588 291374 -532
rect 291430 -588 291498 -532
rect 291554 -588 291622 -532
rect 291678 -588 291774 -532
rect 291154 -1644 291774 -588
rect 309154 4350 309774 8858
rect 309154 4294 309250 4350
rect 309306 4294 309374 4350
rect 309430 4294 309498 4350
rect 309554 4294 309622 4350
rect 309678 4294 309774 4350
rect 309154 4226 309774 4294
rect 309154 4170 309250 4226
rect 309306 4170 309374 4226
rect 309430 4170 309498 4226
rect 309554 4170 309622 4226
rect 309678 4170 309774 4226
rect 309154 4102 309774 4170
rect 309154 4046 309250 4102
rect 309306 4046 309374 4102
rect 309430 4046 309498 4102
rect 309554 4046 309622 4102
rect 309678 4046 309774 4102
rect 309154 3978 309774 4046
rect 309154 3922 309250 3978
rect 309306 3922 309374 3978
rect 309430 3922 309498 3978
rect 309554 3922 309622 3978
rect 309678 3922 309774 3978
rect 309154 -160 309774 3922
rect 309154 -216 309250 -160
rect 309306 -216 309374 -160
rect 309430 -216 309498 -160
rect 309554 -216 309622 -160
rect 309678 -216 309774 -160
rect 309154 -284 309774 -216
rect 309154 -340 309250 -284
rect 309306 -340 309374 -284
rect 309430 -340 309498 -284
rect 309554 -340 309622 -284
rect 309678 -340 309774 -284
rect 309154 -408 309774 -340
rect 309154 -464 309250 -408
rect 309306 -464 309374 -408
rect 309430 -464 309498 -408
rect 309554 -464 309622 -408
rect 309678 -464 309774 -408
rect 309154 -532 309774 -464
rect 309154 -588 309250 -532
rect 309306 -588 309374 -532
rect 309430 -588 309498 -532
rect 309554 -588 309622 -532
rect 309678 -588 309774 -532
rect 309154 -1644 309774 -588
rect 327154 4350 327774 8858
rect 327154 4294 327250 4350
rect 327306 4294 327374 4350
rect 327430 4294 327498 4350
rect 327554 4294 327622 4350
rect 327678 4294 327774 4350
rect 327154 4226 327774 4294
rect 327154 4170 327250 4226
rect 327306 4170 327374 4226
rect 327430 4170 327498 4226
rect 327554 4170 327622 4226
rect 327678 4170 327774 4226
rect 327154 4102 327774 4170
rect 327154 4046 327250 4102
rect 327306 4046 327374 4102
rect 327430 4046 327498 4102
rect 327554 4046 327622 4102
rect 327678 4046 327774 4102
rect 327154 3978 327774 4046
rect 327154 3922 327250 3978
rect 327306 3922 327374 3978
rect 327430 3922 327498 3978
rect 327554 3922 327622 3978
rect 327678 3922 327774 3978
rect 327154 -160 327774 3922
rect 327154 -216 327250 -160
rect 327306 -216 327374 -160
rect 327430 -216 327498 -160
rect 327554 -216 327622 -160
rect 327678 -216 327774 -160
rect 327154 -284 327774 -216
rect 327154 -340 327250 -284
rect 327306 -340 327374 -284
rect 327430 -340 327498 -284
rect 327554 -340 327622 -284
rect 327678 -340 327774 -284
rect 327154 -408 327774 -340
rect 327154 -464 327250 -408
rect 327306 -464 327374 -408
rect 327430 -464 327498 -408
rect 327554 -464 327622 -408
rect 327678 -464 327774 -408
rect 327154 -532 327774 -464
rect 327154 -588 327250 -532
rect 327306 -588 327374 -532
rect 327430 -588 327498 -532
rect 327554 -588 327622 -532
rect 327678 -588 327774 -532
rect 327154 -1644 327774 -588
rect 345154 4350 345774 8858
rect 345154 4294 345250 4350
rect 345306 4294 345374 4350
rect 345430 4294 345498 4350
rect 345554 4294 345622 4350
rect 345678 4294 345774 4350
rect 345154 4226 345774 4294
rect 345154 4170 345250 4226
rect 345306 4170 345374 4226
rect 345430 4170 345498 4226
rect 345554 4170 345622 4226
rect 345678 4170 345774 4226
rect 345154 4102 345774 4170
rect 345154 4046 345250 4102
rect 345306 4046 345374 4102
rect 345430 4046 345498 4102
rect 345554 4046 345622 4102
rect 345678 4046 345774 4102
rect 345154 3978 345774 4046
rect 345154 3922 345250 3978
rect 345306 3922 345374 3978
rect 345430 3922 345498 3978
rect 345554 3922 345622 3978
rect 345678 3922 345774 3978
rect 345154 -160 345774 3922
rect 345154 -216 345250 -160
rect 345306 -216 345374 -160
rect 345430 -216 345498 -160
rect 345554 -216 345622 -160
rect 345678 -216 345774 -160
rect 345154 -284 345774 -216
rect 345154 -340 345250 -284
rect 345306 -340 345374 -284
rect 345430 -340 345498 -284
rect 345554 -340 345622 -284
rect 345678 -340 345774 -284
rect 345154 -408 345774 -340
rect 345154 -464 345250 -408
rect 345306 -464 345374 -408
rect 345430 -464 345498 -408
rect 345554 -464 345622 -408
rect 345678 -464 345774 -408
rect 345154 -532 345774 -464
rect 345154 -588 345250 -532
rect 345306 -588 345374 -532
rect 345430 -588 345498 -532
rect 345554 -588 345622 -532
rect 345678 -588 345774 -532
rect 345154 -1644 345774 -588
rect 363154 4350 363774 8858
rect 376348 6356 376404 156268
rect 376348 6290 376404 6300
rect 378028 160916 378084 160926
rect 378028 159908 378084 160860
rect 378028 4676 378084 159852
rect 378028 4610 378084 4620
rect 378140 155876 378196 155886
rect 363154 4294 363250 4350
rect 363306 4294 363374 4350
rect 363430 4294 363498 4350
rect 363554 4294 363622 4350
rect 363678 4294 363774 4350
rect 363154 4226 363774 4294
rect 363154 4170 363250 4226
rect 363306 4170 363374 4226
rect 363430 4170 363498 4226
rect 363554 4170 363622 4226
rect 363678 4170 363774 4226
rect 363154 4102 363774 4170
rect 363154 4046 363250 4102
rect 363306 4046 363374 4102
rect 363430 4046 363498 4102
rect 363554 4046 363622 4102
rect 363678 4046 363774 4102
rect 363154 3978 363774 4046
rect 363154 3922 363250 3978
rect 363306 3922 363374 3978
rect 363430 3922 363498 3978
rect 363554 3922 363622 3978
rect 363678 3922 363774 3978
rect 363154 -160 363774 3922
rect 378140 2996 378196 155820
rect 378140 2930 378196 2940
rect 381154 148350 381774 165922
rect 381154 148294 381250 148350
rect 381306 148294 381374 148350
rect 381430 148294 381498 148350
rect 381554 148294 381622 148350
rect 381678 148294 381774 148350
rect 381154 148226 381774 148294
rect 381154 148170 381250 148226
rect 381306 148170 381374 148226
rect 381430 148170 381498 148226
rect 381554 148170 381622 148226
rect 381678 148170 381774 148226
rect 381154 148102 381774 148170
rect 381154 148046 381250 148102
rect 381306 148046 381374 148102
rect 381430 148046 381498 148102
rect 381554 148046 381622 148102
rect 381678 148046 381774 148102
rect 381154 147978 381774 148046
rect 381154 147922 381250 147978
rect 381306 147922 381374 147978
rect 381430 147922 381498 147978
rect 381554 147922 381622 147978
rect 381678 147922 381774 147978
rect 381154 130350 381774 147922
rect 381154 130294 381250 130350
rect 381306 130294 381374 130350
rect 381430 130294 381498 130350
rect 381554 130294 381622 130350
rect 381678 130294 381774 130350
rect 381154 130226 381774 130294
rect 381154 130170 381250 130226
rect 381306 130170 381374 130226
rect 381430 130170 381498 130226
rect 381554 130170 381622 130226
rect 381678 130170 381774 130226
rect 381154 130102 381774 130170
rect 381154 130046 381250 130102
rect 381306 130046 381374 130102
rect 381430 130046 381498 130102
rect 381554 130046 381622 130102
rect 381678 130046 381774 130102
rect 381154 129978 381774 130046
rect 381154 129922 381250 129978
rect 381306 129922 381374 129978
rect 381430 129922 381498 129978
rect 381554 129922 381622 129978
rect 381678 129922 381774 129978
rect 381154 112350 381774 129922
rect 381154 112294 381250 112350
rect 381306 112294 381374 112350
rect 381430 112294 381498 112350
rect 381554 112294 381622 112350
rect 381678 112294 381774 112350
rect 381154 112226 381774 112294
rect 381154 112170 381250 112226
rect 381306 112170 381374 112226
rect 381430 112170 381498 112226
rect 381554 112170 381622 112226
rect 381678 112170 381774 112226
rect 381154 112102 381774 112170
rect 381154 112046 381250 112102
rect 381306 112046 381374 112102
rect 381430 112046 381498 112102
rect 381554 112046 381622 112102
rect 381678 112046 381774 112102
rect 381154 111978 381774 112046
rect 381154 111922 381250 111978
rect 381306 111922 381374 111978
rect 381430 111922 381498 111978
rect 381554 111922 381622 111978
rect 381678 111922 381774 111978
rect 381154 94350 381774 111922
rect 381154 94294 381250 94350
rect 381306 94294 381374 94350
rect 381430 94294 381498 94350
rect 381554 94294 381622 94350
rect 381678 94294 381774 94350
rect 381154 94226 381774 94294
rect 381154 94170 381250 94226
rect 381306 94170 381374 94226
rect 381430 94170 381498 94226
rect 381554 94170 381622 94226
rect 381678 94170 381774 94226
rect 381154 94102 381774 94170
rect 381154 94046 381250 94102
rect 381306 94046 381374 94102
rect 381430 94046 381498 94102
rect 381554 94046 381622 94102
rect 381678 94046 381774 94102
rect 381154 93978 381774 94046
rect 381154 93922 381250 93978
rect 381306 93922 381374 93978
rect 381430 93922 381498 93978
rect 381554 93922 381622 93978
rect 381678 93922 381774 93978
rect 381154 76350 381774 93922
rect 381154 76294 381250 76350
rect 381306 76294 381374 76350
rect 381430 76294 381498 76350
rect 381554 76294 381622 76350
rect 381678 76294 381774 76350
rect 381154 76226 381774 76294
rect 381154 76170 381250 76226
rect 381306 76170 381374 76226
rect 381430 76170 381498 76226
rect 381554 76170 381622 76226
rect 381678 76170 381774 76226
rect 381154 76102 381774 76170
rect 381154 76046 381250 76102
rect 381306 76046 381374 76102
rect 381430 76046 381498 76102
rect 381554 76046 381622 76102
rect 381678 76046 381774 76102
rect 381154 75978 381774 76046
rect 381154 75922 381250 75978
rect 381306 75922 381374 75978
rect 381430 75922 381498 75978
rect 381554 75922 381622 75978
rect 381678 75922 381774 75978
rect 381154 58350 381774 75922
rect 381154 58294 381250 58350
rect 381306 58294 381374 58350
rect 381430 58294 381498 58350
rect 381554 58294 381622 58350
rect 381678 58294 381774 58350
rect 381154 58226 381774 58294
rect 381154 58170 381250 58226
rect 381306 58170 381374 58226
rect 381430 58170 381498 58226
rect 381554 58170 381622 58226
rect 381678 58170 381774 58226
rect 381154 58102 381774 58170
rect 381154 58046 381250 58102
rect 381306 58046 381374 58102
rect 381430 58046 381498 58102
rect 381554 58046 381622 58102
rect 381678 58046 381774 58102
rect 381154 57978 381774 58046
rect 381154 57922 381250 57978
rect 381306 57922 381374 57978
rect 381430 57922 381498 57978
rect 381554 57922 381622 57978
rect 381678 57922 381774 57978
rect 381154 40350 381774 57922
rect 381154 40294 381250 40350
rect 381306 40294 381374 40350
rect 381430 40294 381498 40350
rect 381554 40294 381622 40350
rect 381678 40294 381774 40350
rect 381154 40226 381774 40294
rect 381154 40170 381250 40226
rect 381306 40170 381374 40226
rect 381430 40170 381498 40226
rect 381554 40170 381622 40226
rect 381678 40170 381774 40226
rect 381154 40102 381774 40170
rect 381154 40046 381250 40102
rect 381306 40046 381374 40102
rect 381430 40046 381498 40102
rect 381554 40046 381622 40102
rect 381678 40046 381774 40102
rect 381154 39978 381774 40046
rect 381154 39922 381250 39978
rect 381306 39922 381374 39978
rect 381430 39922 381498 39978
rect 381554 39922 381622 39978
rect 381678 39922 381774 39978
rect 381154 22350 381774 39922
rect 381154 22294 381250 22350
rect 381306 22294 381374 22350
rect 381430 22294 381498 22350
rect 381554 22294 381622 22350
rect 381678 22294 381774 22350
rect 381154 22226 381774 22294
rect 381154 22170 381250 22226
rect 381306 22170 381374 22226
rect 381430 22170 381498 22226
rect 381554 22170 381622 22226
rect 381678 22170 381774 22226
rect 381154 22102 381774 22170
rect 381154 22046 381250 22102
rect 381306 22046 381374 22102
rect 381430 22046 381498 22102
rect 381554 22046 381622 22102
rect 381678 22046 381774 22102
rect 381154 21978 381774 22046
rect 381154 21922 381250 21978
rect 381306 21922 381374 21978
rect 381430 21922 381498 21978
rect 381554 21922 381622 21978
rect 381678 21922 381774 21978
rect 381154 4350 381774 21922
rect 381154 4294 381250 4350
rect 381306 4294 381374 4350
rect 381430 4294 381498 4350
rect 381554 4294 381622 4350
rect 381678 4294 381774 4350
rect 381154 4226 381774 4294
rect 381154 4170 381250 4226
rect 381306 4170 381374 4226
rect 381430 4170 381498 4226
rect 381554 4170 381622 4226
rect 381678 4170 381774 4226
rect 381154 4102 381774 4170
rect 381154 4046 381250 4102
rect 381306 4046 381374 4102
rect 381430 4046 381498 4102
rect 381554 4046 381622 4102
rect 381678 4046 381774 4102
rect 381154 3978 381774 4046
rect 381154 3922 381250 3978
rect 381306 3922 381374 3978
rect 381430 3922 381498 3978
rect 381554 3922 381622 3978
rect 381678 3922 381774 3978
rect 363154 -216 363250 -160
rect 363306 -216 363374 -160
rect 363430 -216 363498 -160
rect 363554 -216 363622 -160
rect 363678 -216 363774 -160
rect 363154 -284 363774 -216
rect 363154 -340 363250 -284
rect 363306 -340 363374 -284
rect 363430 -340 363498 -284
rect 363554 -340 363622 -284
rect 363678 -340 363774 -284
rect 363154 -408 363774 -340
rect 363154 -464 363250 -408
rect 363306 -464 363374 -408
rect 363430 -464 363498 -408
rect 363554 -464 363622 -408
rect 363678 -464 363774 -408
rect 363154 -532 363774 -464
rect 363154 -588 363250 -532
rect 363306 -588 363374 -532
rect 363430 -588 363498 -532
rect 363554 -588 363622 -532
rect 363678 -588 363774 -532
rect 363154 -1644 363774 -588
rect 381154 -160 381774 3922
rect 381154 -216 381250 -160
rect 381306 -216 381374 -160
rect 381430 -216 381498 -160
rect 381554 -216 381622 -160
rect 381678 -216 381774 -160
rect 381154 -284 381774 -216
rect 381154 -340 381250 -284
rect 381306 -340 381374 -284
rect 381430 -340 381498 -284
rect 381554 -340 381622 -284
rect 381678 -340 381774 -284
rect 381154 -408 381774 -340
rect 381154 -464 381250 -408
rect 381306 -464 381374 -408
rect 381430 -464 381498 -408
rect 381554 -464 381622 -408
rect 381678 -464 381774 -408
rect 381154 -532 381774 -464
rect 381154 -588 381250 -532
rect 381306 -588 381374 -532
rect 381430 -588 381498 -532
rect 381554 -588 381622 -532
rect 381678 -588 381774 -532
rect 381154 -1644 381774 -588
rect 384874 598172 385494 598268
rect 384874 598116 384970 598172
rect 385026 598116 385094 598172
rect 385150 598116 385218 598172
rect 385274 598116 385342 598172
rect 385398 598116 385494 598172
rect 384874 598048 385494 598116
rect 384874 597992 384970 598048
rect 385026 597992 385094 598048
rect 385150 597992 385218 598048
rect 385274 597992 385342 598048
rect 385398 597992 385494 598048
rect 384874 597924 385494 597992
rect 384874 597868 384970 597924
rect 385026 597868 385094 597924
rect 385150 597868 385218 597924
rect 385274 597868 385342 597924
rect 385398 597868 385494 597924
rect 384874 597800 385494 597868
rect 384874 597744 384970 597800
rect 385026 597744 385094 597800
rect 385150 597744 385218 597800
rect 385274 597744 385342 597800
rect 385398 597744 385494 597800
rect 384874 586350 385494 597744
rect 384874 586294 384970 586350
rect 385026 586294 385094 586350
rect 385150 586294 385218 586350
rect 385274 586294 385342 586350
rect 385398 586294 385494 586350
rect 384874 586226 385494 586294
rect 384874 586170 384970 586226
rect 385026 586170 385094 586226
rect 385150 586170 385218 586226
rect 385274 586170 385342 586226
rect 385398 586170 385494 586226
rect 384874 586102 385494 586170
rect 384874 586046 384970 586102
rect 385026 586046 385094 586102
rect 385150 586046 385218 586102
rect 385274 586046 385342 586102
rect 385398 586046 385494 586102
rect 384874 585978 385494 586046
rect 384874 585922 384970 585978
rect 385026 585922 385094 585978
rect 385150 585922 385218 585978
rect 385274 585922 385342 585978
rect 385398 585922 385494 585978
rect 384874 568350 385494 585922
rect 384874 568294 384970 568350
rect 385026 568294 385094 568350
rect 385150 568294 385218 568350
rect 385274 568294 385342 568350
rect 385398 568294 385494 568350
rect 384874 568226 385494 568294
rect 384874 568170 384970 568226
rect 385026 568170 385094 568226
rect 385150 568170 385218 568226
rect 385274 568170 385342 568226
rect 385398 568170 385494 568226
rect 384874 568102 385494 568170
rect 384874 568046 384970 568102
rect 385026 568046 385094 568102
rect 385150 568046 385218 568102
rect 385274 568046 385342 568102
rect 385398 568046 385494 568102
rect 384874 567978 385494 568046
rect 384874 567922 384970 567978
rect 385026 567922 385094 567978
rect 385150 567922 385218 567978
rect 385274 567922 385342 567978
rect 385398 567922 385494 567978
rect 384874 550350 385494 567922
rect 384874 550294 384970 550350
rect 385026 550294 385094 550350
rect 385150 550294 385218 550350
rect 385274 550294 385342 550350
rect 385398 550294 385494 550350
rect 384874 550226 385494 550294
rect 384874 550170 384970 550226
rect 385026 550170 385094 550226
rect 385150 550170 385218 550226
rect 385274 550170 385342 550226
rect 385398 550170 385494 550226
rect 384874 550102 385494 550170
rect 384874 550046 384970 550102
rect 385026 550046 385094 550102
rect 385150 550046 385218 550102
rect 385274 550046 385342 550102
rect 385398 550046 385494 550102
rect 384874 549978 385494 550046
rect 384874 549922 384970 549978
rect 385026 549922 385094 549978
rect 385150 549922 385218 549978
rect 385274 549922 385342 549978
rect 385398 549922 385494 549978
rect 384874 532350 385494 549922
rect 384874 532294 384970 532350
rect 385026 532294 385094 532350
rect 385150 532294 385218 532350
rect 385274 532294 385342 532350
rect 385398 532294 385494 532350
rect 384874 532226 385494 532294
rect 384874 532170 384970 532226
rect 385026 532170 385094 532226
rect 385150 532170 385218 532226
rect 385274 532170 385342 532226
rect 385398 532170 385494 532226
rect 384874 532102 385494 532170
rect 384874 532046 384970 532102
rect 385026 532046 385094 532102
rect 385150 532046 385218 532102
rect 385274 532046 385342 532102
rect 385398 532046 385494 532102
rect 384874 531978 385494 532046
rect 384874 531922 384970 531978
rect 385026 531922 385094 531978
rect 385150 531922 385218 531978
rect 385274 531922 385342 531978
rect 385398 531922 385494 531978
rect 384874 514350 385494 531922
rect 384874 514294 384970 514350
rect 385026 514294 385094 514350
rect 385150 514294 385218 514350
rect 385274 514294 385342 514350
rect 385398 514294 385494 514350
rect 384874 514226 385494 514294
rect 384874 514170 384970 514226
rect 385026 514170 385094 514226
rect 385150 514170 385218 514226
rect 385274 514170 385342 514226
rect 385398 514170 385494 514226
rect 384874 514102 385494 514170
rect 384874 514046 384970 514102
rect 385026 514046 385094 514102
rect 385150 514046 385218 514102
rect 385274 514046 385342 514102
rect 385398 514046 385494 514102
rect 384874 513978 385494 514046
rect 384874 513922 384970 513978
rect 385026 513922 385094 513978
rect 385150 513922 385218 513978
rect 385274 513922 385342 513978
rect 385398 513922 385494 513978
rect 384874 496350 385494 513922
rect 384874 496294 384970 496350
rect 385026 496294 385094 496350
rect 385150 496294 385218 496350
rect 385274 496294 385342 496350
rect 385398 496294 385494 496350
rect 384874 496226 385494 496294
rect 384874 496170 384970 496226
rect 385026 496170 385094 496226
rect 385150 496170 385218 496226
rect 385274 496170 385342 496226
rect 385398 496170 385494 496226
rect 384874 496102 385494 496170
rect 384874 496046 384970 496102
rect 385026 496046 385094 496102
rect 385150 496046 385218 496102
rect 385274 496046 385342 496102
rect 385398 496046 385494 496102
rect 384874 495978 385494 496046
rect 384874 495922 384970 495978
rect 385026 495922 385094 495978
rect 385150 495922 385218 495978
rect 385274 495922 385342 495978
rect 385398 495922 385494 495978
rect 384874 478350 385494 495922
rect 384874 478294 384970 478350
rect 385026 478294 385094 478350
rect 385150 478294 385218 478350
rect 385274 478294 385342 478350
rect 385398 478294 385494 478350
rect 384874 478226 385494 478294
rect 384874 478170 384970 478226
rect 385026 478170 385094 478226
rect 385150 478170 385218 478226
rect 385274 478170 385342 478226
rect 385398 478170 385494 478226
rect 384874 478102 385494 478170
rect 384874 478046 384970 478102
rect 385026 478046 385094 478102
rect 385150 478046 385218 478102
rect 385274 478046 385342 478102
rect 385398 478046 385494 478102
rect 384874 477978 385494 478046
rect 384874 477922 384970 477978
rect 385026 477922 385094 477978
rect 385150 477922 385218 477978
rect 385274 477922 385342 477978
rect 385398 477922 385494 477978
rect 384874 460350 385494 477922
rect 384874 460294 384970 460350
rect 385026 460294 385094 460350
rect 385150 460294 385218 460350
rect 385274 460294 385342 460350
rect 385398 460294 385494 460350
rect 384874 460226 385494 460294
rect 384874 460170 384970 460226
rect 385026 460170 385094 460226
rect 385150 460170 385218 460226
rect 385274 460170 385342 460226
rect 385398 460170 385494 460226
rect 384874 460102 385494 460170
rect 384874 460046 384970 460102
rect 385026 460046 385094 460102
rect 385150 460046 385218 460102
rect 385274 460046 385342 460102
rect 385398 460046 385494 460102
rect 384874 459978 385494 460046
rect 384874 459922 384970 459978
rect 385026 459922 385094 459978
rect 385150 459922 385218 459978
rect 385274 459922 385342 459978
rect 385398 459922 385494 459978
rect 384874 442350 385494 459922
rect 384874 442294 384970 442350
rect 385026 442294 385094 442350
rect 385150 442294 385218 442350
rect 385274 442294 385342 442350
rect 385398 442294 385494 442350
rect 384874 442226 385494 442294
rect 384874 442170 384970 442226
rect 385026 442170 385094 442226
rect 385150 442170 385218 442226
rect 385274 442170 385342 442226
rect 385398 442170 385494 442226
rect 384874 442102 385494 442170
rect 384874 442046 384970 442102
rect 385026 442046 385094 442102
rect 385150 442046 385218 442102
rect 385274 442046 385342 442102
rect 385398 442046 385494 442102
rect 384874 441978 385494 442046
rect 384874 441922 384970 441978
rect 385026 441922 385094 441978
rect 385150 441922 385218 441978
rect 385274 441922 385342 441978
rect 385398 441922 385494 441978
rect 384874 424350 385494 441922
rect 384874 424294 384970 424350
rect 385026 424294 385094 424350
rect 385150 424294 385218 424350
rect 385274 424294 385342 424350
rect 385398 424294 385494 424350
rect 384874 424226 385494 424294
rect 384874 424170 384970 424226
rect 385026 424170 385094 424226
rect 385150 424170 385218 424226
rect 385274 424170 385342 424226
rect 385398 424170 385494 424226
rect 384874 424102 385494 424170
rect 384874 424046 384970 424102
rect 385026 424046 385094 424102
rect 385150 424046 385218 424102
rect 385274 424046 385342 424102
rect 385398 424046 385494 424102
rect 384874 423978 385494 424046
rect 384874 423922 384970 423978
rect 385026 423922 385094 423978
rect 385150 423922 385218 423978
rect 385274 423922 385342 423978
rect 385398 423922 385494 423978
rect 384874 406350 385494 423922
rect 384874 406294 384970 406350
rect 385026 406294 385094 406350
rect 385150 406294 385218 406350
rect 385274 406294 385342 406350
rect 385398 406294 385494 406350
rect 384874 406226 385494 406294
rect 384874 406170 384970 406226
rect 385026 406170 385094 406226
rect 385150 406170 385218 406226
rect 385274 406170 385342 406226
rect 385398 406170 385494 406226
rect 384874 406102 385494 406170
rect 384874 406046 384970 406102
rect 385026 406046 385094 406102
rect 385150 406046 385218 406102
rect 385274 406046 385342 406102
rect 385398 406046 385494 406102
rect 384874 405978 385494 406046
rect 384874 405922 384970 405978
rect 385026 405922 385094 405978
rect 385150 405922 385218 405978
rect 385274 405922 385342 405978
rect 385398 405922 385494 405978
rect 384874 388350 385494 405922
rect 384874 388294 384970 388350
rect 385026 388294 385094 388350
rect 385150 388294 385218 388350
rect 385274 388294 385342 388350
rect 385398 388294 385494 388350
rect 384874 388226 385494 388294
rect 384874 388170 384970 388226
rect 385026 388170 385094 388226
rect 385150 388170 385218 388226
rect 385274 388170 385342 388226
rect 385398 388170 385494 388226
rect 384874 388102 385494 388170
rect 384874 388046 384970 388102
rect 385026 388046 385094 388102
rect 385150 388046 385218 388102
rect 385274 388046 385342 388102
rect 385398 388046 385494 388102
rect 384874 387978 385494 388046
rect 384874 387922 384970 387978
rect 385026 387922 385094 387978
rect 385150 387922 385218 387978
rect 385274 387922 385342 387978
rect 385398 387922 385494 387978
rect 384874 370350 385494 387922
rect 384874 370294 384970 370350
rect 385026 370294 385094 370350
rect 385150 370294 385218 370350
rect 385274 370294 385342 370350
rect 385398 370294 385494 370350
rect 384874 370226 385494 370294
rect 384874 370170 384970 370226
rect 385026 370170 385094 370226
rect 385150 370170 385218 370226
rect 385274 370170 385342 370226
rect 385398 370170 385494 370226
rect 384874 370102 385494 370170
rect 384874 370046 384970 370102
rect 385026 370046 385094 370102
rect 385150 370046 385218 370102
rect 385274 370046 385342 370102
rect 385398 370046 385494 370102
rect 384874 369978 385494 370046
rect 384874 369922 384970 369978
rect 385026 369922 385094 369978
rect 385150 369922 385218 369978
rect 385274 369922 385342 369978
rect 385398 369922 385494 369978
rect 384874 352350 385494 369922
rect 384874 352294 384970 352350
rect 385026 352294 385094 352350
rect 385150 352294 385218 352350
rect 385274 352294 385342 352350
rect 385398 352294 385494 352350
rect 384874 352226 385494 352294
rect 384874 352170 384970 352226
rect 385026 352170 385094 352226
rect 385150 352170 385218 352226
rect 385274 352170 385342 352226
rect 385398 352170 385494 352226
rect 384874 352102 385494 352170
rect 384874 352046 384970 352102
rect 385026 352046 385094 352102
rect 385150 352046 385218 352102
rect 385274 352046 385342 352102
rect 385398 352046 385494 352102
rect 384874 351978 385494 352046
rect 384874 351922 384970 351978
rect 385026 351922 385094 351978
rect 385150 351922 385218 351978
rect 385274 351922 385342 351978
rect 385398 351922 385494 351978
rect 384874 334350 385494 351922
rect 384874 334294 384970 334350
rect 385026 334294 385094 334350
rect 385150 334294 385218 334350
rect 385274 334294 385342 334350
rect 385398 334294 385494 334350
rect 384874 334226 385494 334294
rect 384874 334170 384970 334226
rect 385026 334170 385094 334226
rect 385150 334170 385218 334226
rect 385274 334170 385342 334226
rect 385398 334170 385494 334226
rect 384874 334102 385494 334170
rect 384874 334046 384970 334102
rect 385026 334046 385094 334102
rect 385150 334046 385218 334102
rect 385274 334046 385342 334102
rect 385398 334046 385494 334102
rect 384874 333978 385494 334046
rect 384874 333922 384970 333978
rect 385026 333922 385094 333978
rect 385150 333922 385218 333978
rect 385274 333922 385342 333978
rect 385398 333922 385494 333978
rect 384874 316350 385494 333922
rect 384874 316294 384970 316350
rect 385026 316294 385094 316350
rect 385150 316294 385218 316350
rect 385274 316294 385342 316350
rect 385398 316294 385494 316350
rect 384874 316226 385494 316294
rect 384874 316170 384970 316226
rect 385026 316170 385094 316226
rect 385150 316170 385218 316226
rect 385274 316170 385342 316226
rect 385398 316170 385494 316226
rect 384874 316102 385494 316170
rect 384874 316046 384970 316102
rect 385026 316046 385094 316102
rect 385150 316046 385218 316102
rect 385274 316046 385342 316102
rect 385398 316046 385494 316102
rect 384874 315978 385494 316046
rect 384874 315922 384970 315978
rect 385026 315922 385094 315978
rect 385150 315922 385218 315978
rect 385274 315922 385342 315978
rect 385398 315922 385494 315978
rect 384874 298350 385494 315922
rect 399154 597212 399774 598268
rect 399154 597156 399250 597212
rect 399306 597156 399374 597212
rect 399430 597156 399498 597212
rect 399554 597156 399622 597212
rect 399678 597156 399774 597212
rect 399154 597088 399774 597156
rect 399154 597032 399250 597088
rect 399306 597032 399374 597088
rect 399430 597032 399498 597088
rect 399554 597032 399622 597088
rect 399678 597032 399774 597088
rect 399154 596964 399774 597032
rect 399154 596908 399250 596964
rect 399306 596908 399374 596964
rect 399430 596908 399498 596964
rect 399554 596908 399622 596964
rect 399678 596908 399774 596964
rect 399154 596840 399774 596908
rect 399154 596784 399250 596840
rect 399306 596784 399374 596840
rect 399430 596784 399498 596840
rect 399554 596784 399622 596840
rect 399678 596784 399774 596840
rect 399154 580350 399774 596784
rect 399154 580294 399250 580350
rect 399306 580294 399374 580350
rect 399430 580294 399498 580350
rect 399554 580294 399622 580350
rect 399678 580294 399774 580350
rect 399154 580226 399774 580294
rect 399154 580170 399250 580226
rect 399306 580170 399374 580226
rect 399430 580170 399498 580226
rect 399554 580170 399622 580226
rect 399678 580170 399774 580226
rect 399154 580102 399774 580170
rect 399154 580046 399250 580102
rect 399306 580046 399374 580102
rect 399430 580046 399498 580102
rect 399554 580046 399622 580102
rect 399678 580046 399774 580102
rect 399154 579978 399774 580046
rect 399154 579922 399250 579978
rect 399306 579922 399374 579978
rect 399430 579922 399498 579978
rect 399554 579922 399622 579978
rect 399678 579922 399774 579978
rect 399154 562350 399774 579922
rect 399154 562294 399250 562350
rect 399306 562294 399374 562350
rect 399430 562294 399498 562350
rect 399554 562294 399622 562350
rect 399678 562294 399774 562350
rect 399154 562226 399774 562294
rect 399154 562170 399250 562226
rect 399306 562170 399374 562226
rect 399430 562170 399498 562226
rect 399554 562170 399622 562226
rect 399678 562170 399774 562226
rect 399154 562102 399774 562170
rect 399154 562046 399250 562102
rect 399306 562046 399374 562102
rect 399430 562046 399498 562102
rect 399554 562046 399622 562102
rect 399678 562046 399774 562102
rect 399154 561978 399774 562046
rect 399154 561922 399250 561978
rect 399306 561922 399374 561978
rect 399430 561922 399498 561978
rect 399554 561922 399622 561978
rect 399678 561922 399774 561978
rect 399154 544350 399774 561922
rect 399154 544294 399250 544350
rect 399306 544294 399374 544350
rect 399430 544294 399498 544350
rect 399554 544294 399622 544350
rect 399678 544294 399774 544350
rect 399154 544226 399774 544294
rect 399154 544170 399250 544226
rect 399306 544170 399374 544226
rect 399430 544170 399498 544226
rect 399554 544170 399622 544226
rect 399678 544170 399774 544226
rect 399154 544102 399774 544170
rect 399154 544046 399250 544102
rect 399306 544046 399374 544102
rect 399430 544046 399498 544102
rect 399554 544046 399622 544102
rect 399678 544046 399774 544102
rect 399154 543978 399774 544046
rect 399154 543922 399250 543978
rect 399306 543922 399374 543978
rect 399430 543922 399498 543978
rect 399554 543922 399622 543978
rect 399678 543922 399774 543978
rect 399154 526350 399774 543922
rect 399154 526294 399250 526350
rect 399306 526294 399374 526350
rect 399430 526294 399498 526350
rect 399554 526294 399622 526350
rect 399678 526294 399774 526350
rect 399154 526226 399774 526294
rect 399154 526170 399250 526226
rect 399306 526170 399374 526226
rect 399430 526170 399498 526226
rect 399554 526170 399622 526226
rect 399678 526170 399774 526226
rect 399154 526102 399774 526170
rect 399154 526046 399250 526102
rect 399306 526046 399374 526102
rect 399430 526046 399498 526102
rect 399554 526046 399622 526102
rect 399678 526046 399774 526102
rect 399154 525978 399774 526046
rect 399154 525922 399250 525978
rect 399306 525922 399374 525978
rect 399430 525922 399498 525978
rect 399554 525922 399622 525978
rect 399678 525922 399774 525978
rect 399154 508350 399774 525922
rect 399154 508294 399250 508350
rect 399306 508294 399374 508350
rect 399430 508294 399498 508350
rect 399554 508294 399622 508350
rect 399678 508294 399774 508350
rect 399154 508226 399774 508294
rect 399154 508170 399250 508226
rect 399306 508170 399374 508226
rect 399430 508170 399498 508226
rect 399554 508170 399622 508226
rect 399678 508170 399774 508226
rect 399154 508102 399774 508170
rect 399154 508046 399250 508102
rect 399306 508046 399374 508102
rect 399430 508046 399498 508102
rect 399554 508046 399622 508102
rect 399678 508046 399774 508102
rect 399154 507978 399774 508046
rect 399154 507922 399250 507978
rect 399306 507922 399374 507978
rect 399430 507922 399498 507978
rect 399554 507922 399622 507978
rect 399678 507922 399774 507978
rect 399154 490350 399774 507922
rect 399154 490294 399250 490350
rect 399306 490294 399374 490350
rect 399430 490294 399498 490350
rect 399554 490294 399622 490350
rect 399678 490294 399774 490350
rect 399154 490226 399774 490294
rect 399154 490170 399250 490226
rect 399306 490170 399374 490226
rect 399430 490170 399498 490226
rect 399554 490170 399622 490226
rect 399678 490170 399774 490226
rect 399154 490102 399774 490170
rect 399154 490046 399250 490102
rect 399306 490046 399374 490102
rect 399430 490046 399498 490102
rect 399554 490046 399622 490102
rect 399678 490046 399774 490102
rect 399154 489978 399774 490046
rect 399154 489922 399250 489978
rect 399306 489922 399374 489978
rect 399430 489922 399498 489978
rect 399554 489922 399622 489978
rect 399678 489922 399774 489978
rect 399154 472350 399774 489922
rect 399154 472294 399250 472350
rect 399306 472294 399374 472350
rect 399430 472294 399498 472350
rect 399554 472294 399622 472350
rect 399678 472294 399774 472350
rect 399154 472226 399774 472294
rect 399154 472170 399250 472226
rect 399306 472170 399374 472226
rect 399430 472170 399498 472226
rect 399554 472170 399622 472226
rect 399678 472170 399774 472226
rect 399154 472102 399774 472170
rect 399154 472046 399250 472102
rect 399306 472046 399374 472102
rect 399430 472046 399498 472102
rect 399554 472046 399622 472102
rect 399678 472046 399774 472102
rect 399154 471978 399774 472046
rect 399154 471922 399250 471978
rect 399306 471922 399374 471978
rect 399430 471922 399498 471978
rect 399554 471922 399622 471978
rect 399678 471922 399774 471978
rect 399154 454350 399774 471922
rect 399154 454294 399250 454350
rect 399306 454294 399374 454350
rect 399430 454294 399498 454350
rect 399554 454294 399622 454350
rect 399678 454294 399774 454350
rect 399154 454226 399774 454294
rect 399154 454170 399250 454226
rect 399306 454170 399374 454226
rect 399430 454170 399498 454226
rect 399554 454170 399622 454226
rect 399678 454170 399774 454226
rect 399154 454102 399774 454170
rect 399154 454046 399250 454102
rect 399306 454046 399374 454102
rect 399430 454046 399498 454102
rect 399554 454046 399622 454102
rect 399678 454046 399774 454102
rect 399154 453978 399774 454046
rect 399154 453922 399250 453978
rect 399306 453922 399374 453978
rect 399430 453922 399498 453978
rect 399554 453922 399622 453978
rect 399678 453922 399774 453978
rect 399154 436350 399774 453922
rect 399154 436294 399250 436350
rect 399306 436294 399374 436350
rect 399430 436294 399498 436350
rect 399554 436294 399622 436350
rect 399678 436294 399774 436350
rect 399154 436226 399774 436294
rect 399154 436170 399250 436226
rect 399306 436170 399374 436226
rect 399430 436170 399498 436226
rect 399554 436170 399622 436226
rect 399678 436170 399774 436226
rect 399154 436102 399774 436170
rect 399154 436046 399250 436102
rect 399306 436046 399374 436102
rect 399430 436046 399498 436102
rect 399554 436046 399622 436102
rect 399678 436046 399774 436102
rect 399154 435978 399774 436046
rect 399154 435922 399250 435978
rect 399306 435922 399374 435978
rect 399430 435922 399498 435978
rect 399554 435922 399622 435978
rect 399678 435922 399774 435978
rect 399154 418350 399774 435922
rect 399154 418294 399250 418350
rect 399306 418294 399374 418350
rect 399430 418294 399498 418350
rect 399554 418294 399622 418350
rect 399678 418294 399774 418350
rect 399154 418226 399774 418294
rect 399154 418170 399250 418226
rect 399306 418170 399374 418226
rect 399430 418170 399498 418226
rect 399554 418170 399622 418226
rect 399678 418170 399774 418226
rect 399154 418102 399774 418170
rect 399154 418046 399250 418102
rect 399306 418046 399374 418102
rect 399430 418046 399498 418102
rect 399554 418046 399622 418102
rect 399678 418046 399774 418102
rect 399154 417978 399774 418046
rect 399154 417922 399250 417978
rect 399306 417922 399374 417978
rect 399430 417922 399498 417978
rect 399554 417922 399622 417978
rect 399678 417922 399774 417978
rect 399154 400350 399774 417922
rect 399154 400294 399250 400350
rect 399306 400294 399374 400350
rect 399430 400294 399498 400350
rect 399554 400294 399622 400350
rect 399678 400294 399774 400350
rect 399154 400226 399774 400294
rect 399154 400170 399250 400226
rect 399306 400170 399374 400226
rect 399430 400170 399498 400226
rect 399554 400170 399622 400226
rect 399678 400170 399774 400226
rect 399154 400102 399774 400170
rect 399154 400046 399250 400102
rect 399306 400046 399374 400102
rect 399430 400046 399498 400102
rect 399554 400046 399622 400102
rect 399678 400046 399774 400102
rect 399154 399978 399774 400046
rect 399154 399922 399250 399978
rect 399306 399922 399374 399978
rect 399430 399922 399498 399978
rect 399554 399922 399622 399978
rect 399678 399922 399774 399978
rect 399154 382350 399774 399922
rect 399154 382294 399250 382350
rect 399306 382294 399374 382350
rect 399430 382294 399498 382350
rect 399554 382294 399622 382350
rect 399678 382294 399774 382350
rect 399154 382226 399774 382294
rect 399154 382170 399250 382226
rect 399306 382170 399374 382226
rect 399430 382170 399498 382226
rect 399554 382170 399622 382226
rect 399678 382170 399774 382226
rect 399154 382102 399774 382170
rect 399154 382046 399250 382102
rect 399306 382046 399374 382102
rect 399430 382046 399498 382102
rect 399554 382046 399622 382102
rect 399678 382046 399774 382102
rect 399154 381978 399774 382046
rect 399154 381922 399250 381978
rect 399306 381922 399374 381978
rect 399430 381922 399498 381978
rect 399554 381922 399622 381978
rect 399678 381922 399774 381978
rect 399154 364350 399774 381922
rect 399154 364294 399250 364350
rect 399306 364294 399374 364350
rect 399430 364294 399498 364350
rect 399554 364294 399622 364350
rect 399678 364294 399774 364350
rect 399154 364226 399774 364294
rect 399154 364170 399250 364226
rect 399306 364170 399374 364226
rect 399430 364170 399498 364226
rect 399554 364170 399622 364226
rect 399678 364170 399774 364226
rect 399154 364102 399774 364170
rect 399154 364046 399250 364102
rect 399306 364046 399374 364102
rect 399430 364046 399498 364102
rect 399554 364046 399622 364102
rect 399678 364046 399774 364102
rect 399154 363978 399774 364046
rect 399154 363922 399250 363978
rect 399306 363922 399374 363978
rect 399430 363922 399498 363978
rect 399554 363922 399622 363978
rect 399678 363922 399774 363978
rect 399154 346350 399774 363922
rect 399154 346294 399250 346350
rect 399306 346294 399374 346350
rect 399430 346294 399498 346350
rect 399554 346294 399622 346350
rect 399678 346294 399774 346350
rect 399154 346226 399774 346294
rect 399154 346170 399250 346226
rect 399306 346170 399374 346226
rect 399430 346170 399498 346226
rect 399554 346170 399622 346226
rect 399678 346170 399774 346226
rect 399154 346102 399774 346170
rect 399154 346046 399250 346102
rect 399306 346046 399374 346102
rect 399430 346046 399498 346102
rect 399554 346046 399622 346102
rect 399678 346046 399774 346102
rect 399154 345978 399774 346046
rect 399154 345922 399250 345978
rect 399306 345922 399374 345978
rect 399430 345922 399498 345978
rect 399554 345922 399622 345978
rect 399678 345922 399774 345978
rect 399154 328350 399774 345922
rect 399154 328294 399250 328350
rect 399306 328294 399374 328350
rect 399430 328294 399498 328350
rect 399554 328294 399622 328350
rect 399678 328294 399774 328350
rect 399154 328226 399774 328294
rect 399154 328170 399250 328226
rect 399306 328170 399374 328226
rect 399430 328170 399498 328226
rect 399554 328170 399622 328226
rect 399678 328170 399774 328226
rect 399154 328102 399774 328170
rect 399154 328046 399250 328102
rect 399306 328046 399374 328102
rect 399430 328046 399498 328102
rect 399554 328046 399622 328102
rect 399678 328046 399774 328102
rect 399154 327978 399774 328046
rect 399154 327922 399250 327978
rect 399306 327922 399374 327978
rect 399430 327922 399498 327978
rect 399554 327922 399622 327978
rect 399678 327922 399774 327978
rect 399154 310350 399774 327922
rect 399154 310294 399250 310350
rect 399306 310294 399374 310350
rect 399430 310294 399498 310350
rect 399554 310294 399622 310350
rect 399678 310294 399774 310350
rect 399154 310226 399774 310294
rect 399154 310170 399250 310226
rect 399306 310170 399374 310226
rect 399430 310170 399498 310226
rect 399554 310170 399622 310226
rect 399678 310170 399774 310226
rect 399154 310102 399774 310170
rect 399154 310046 399250 310102
rect 399306 310046 399374 310102
rect 399430 310046 399498 310102
rect 399554 310046 399622 310102
rect 399678 310046 399774 310102
rect 399154 309978 399774 310046
rect 399154 309922 399250 309978
rect 399306 309922 399374 309978
rect 399430 309922 399498 309978
rect 399554 309922 399622 309978
rect 399678 309922 399774 309978
rect 384874 298294 384970 298350
rect 385026 298294 385094 298350
rect 385150 298294 385218 298350
rect 385274 298294 385342 298350
rect 385398 298294 385494 298350
rect 384874 298226 385494 298294
rect 384874 298170 384970 298226
rect 385026 298170 385094 298226
rect 385150 298170 385218 298226
rect 385274 298170 385342 298226
rect 385398 298170 385494 298226
rect 384874 298102 385494 298170
rect 384874 298046 384970 298102
rect 385026 298046 385094 298102
rect 385150 298046 385218 298102
rect 385274 298046 385342 298102
rect 385398 298046 385494 298102
rect 384874 297978 385494 298046
rect 384874 297922 384970 297978
rect 385026 297922 385094 297978
rect 385150 297922 385218 297978
rect 385274 297922 385342 297978
rect 385398 297922 385494 297978
rect 384874 280350 385494 297922
rect 384874 280294 384970 280350
rect 385026 280294 385094 280350
rect 385150 280294 385218 280350
rect 385274 280294 385342 280350
rect 385398 280294 385494 280350
rect 384874 280226 385494 280294
rect 384874 280170 384970 280226
rect 385026 280170 385094 280226
rect 385150 280170 385218 280226
rect 385274 280170 385342 280226
rect 385398 280170 385494 280226
rect 384874 280102 385494 280170
rect 384874 280046 384970 280102
rect 385026 280046 385094 280102
rect 385150 280046 385218 280102
rect 385274 280046 385342 280102
rect 385398 280046 385494 280102
rect 384874 279978 385494 280046
rect 384874 279922 384970 279978
rect 385026 279922 385094 279978
rect 385150 279922 385218 279978
rect 385274 279922 385342 279978
rect 385398 279922 385494 279978
rect 384874 262350 385494 279922
rect 384874 262294 384970 262350
rect 385026 262294 385094 262350
rect 385150 262294 385218 262350
rect 385274 262294 385342 262350
rect 385398 262294 385494 262350
rect 384874 262226 385494 262294
rect 384874 262170 384970 262226
rect 385026 262170 385094 262226
rect 385150 262170 385218 262226
rect 385274 262170 385342 262226
rect 385398 262170 385494 262226
rect 384874 262102 385494 262170
rect 384874 262046 384970 262102
rect 385026 262046 385094 262102
rect 385150 262046 385218 262102
rect 385274 262046 385342 262102
rect 385398 262046 385494 262102
rect 384874 261978 385494 262046
rect 384874 261922 384970 261978
rect 385026 261922 385094 261978
rect 385150 261922 385218 261978
rect 385274 261922 385342 261978
rect 385398 261922 385494 261978
rect 384874 244350 385494 261922
rect 384874 244294 384970 244350
rect 385026 244294 385094 244350
rect 385150 244294 385218 244350
rect 385274 244294 385342 244350
rect 385398 244294 385494 244350
rect 384874 244226 385494 244294
rect 384874 244170 384970 244226
rect 385026 244170 385094 244226
rect 385150 244170 385218 244226
rect 385274 244170 385342 244226
rect 385398 244170 385494 244226
rect 384874 244102 385494 244170
rect 384874 244046 384970 244102
rect 385026 244046 385094 244102
rect 385150 244046 385218 244102
rect 385274 244046 385342 244102
rect 385398 244046 385494 244102
rect 384874 243978 385494 244046
rect 384874 243922 384970 243978
rect 385026 243922 385094 243978
rect 385150 243922 385218 243978
rect 385274 243922 385342 243978
rect 385398 243922 385494 243978
rect 384874 226350 385494 243922
rect 384874 226294 384970 226350
rect 385026 226294 385094 226350
rect 385150 226294 385218 226350
rect 385274 226294 385342 226350
rect 385398 226294 385494 226350
rect 384874 226226 385494 226294
rect 384874 226170 384970 226226
rect 385026 226170 385094 226226
rect 385150 226170 385218 226226
rect 385274 226170 385342 226226
rect 385398 226170 385494 226226
rect 384874 226102 385494 226170
rect 384874 226046 384970 226102
rect 385026 226046 385094 226102
rect 385150 226046 385218 226102
rect 385274 226046 385342 226102
rect 385398 226046 385494 226102
rect 384874 225978 385494 226046
rect 384874 225922 384970 225978
rect 385026 225922 385094 225978
rect 385150 225922 385218 225978
rect 385274 225922 385342 225978
rect 385398 225922 385494 225978
rect 384874 208350 385494 225922
rect 384874 208294 384970 208350
rect 385026 208294 385094 208350
rect 385150 208294 385218 208350
rect 385274 208294 385342 208350
rect 385398 208294 385494 208350
rect 384874 208226 385494 208294
rect 384874 208170 384970 208226
rect 385026 208170 385094 208226
rect 385150 208170 385218 208226
rect 385274 208170 385342 208226
rect 385398 208170 385494 208226
rect 384874 208102 385494 208170
rect 384874 208046 384970 208102
rect 385026 208046 385094 208102
rect 385150 208046 385218 208102
rect 385274 208046 385342 208102
rect 385398 208046 385494 208102
rect 384874 207978 385494 208046
rect 384874 207922 384970 207978
rect 385026 207922 385094 207978
rect 385150 207922 385218 207978
rect 385274 207922 385342 207978
rect 385398 207922 385494 207978
rect 384874 190350 385494 207922
rect 384874 190294 384970 190350
rect 385026 190294 385094 190350
rect 385150 190294 385218 190350
rect 385274 190294 385342 190350
rect 385398 190294 385494 190350
rect 384874 190226 385494 190294
rect 384874 190170 384970 190226
rect 385026 190170 385094 190226
rect 385150 190170 385218 190226
rect 385274 190170 385342 190226
rect 385398 190170 385494 190226
rect 384874 190102 385494 190170
rect 384874 190046 384970 190102
rect 385026 190046 385094 190102
rect 385150 190046 385218 190102
rect 385274 190046 385342 190102
rect 385398 190046 385494 190102
rect 384874 189978 385494 190046
rect 384874 189922 384970 189978
rect 385026 189922 385094 189978
rect 385150 189922 385218 189978
rect 385274 189922 385342 189978
rect 385398 189922 385494 189978
rect 384874 172350 385494 189922
rect 384874 172294 384970 172350
rect 385026 172294 385094 172350
rect 385150 172294 385218 172350
rect 385274 172294 385342 172350
rect 385398 172294 385494 172350
rect 384874 172226 385494 172294
rect 384874 172170 384970 172226
rect 385026 172170 385094 172226
rect 385150 172170 385218 172226
rect 385274 172170 385342 172226
rect 385398 172170 385494 172226
rect 384874 172102 385494 172170
rect 384874 172046 384970 172102
rect 385026 172046 385094 172102
rect 385150 172046 385218 172102
rect 385274 172046 385342 172102
rect 385398 172046 385494 172102
rect 384874 171978 385494 172046
rect 384874 171922 384970 171978
rect 385026 171922 385094 171978
rect 385150 171922 385218 171978
rect 385274 171922 385342 171978
rect 385398 171922 385494 171978
rect 384874 154350 385494 171922
rect 397628 303380 397684 303390
rect 397628 300804 397684 303324
rect 397628 159460 397684 300748
rect 397628 159394 397684 159404
rect 399154 292350 399774 309922
rect 399154 292294 399250 292350
rect 399306 292294 399374 292350
rect 399430 292294 399498 292350
rect 399554 292294 399622 292350
rect 399678 292294 399774 292350
rect 399154 292226 399774 292294
rect 399154 292170 399250 292226
rect 399306 292170 399374 292226
rect 399430 292170 399498 292226
rect 399554 292170 399622 292226
rect 399678 292170 399774 292226
rect 399154 292102 399774 292170
rect 399154 292046 399250 292102
rect 399306 292046 399374 292102
rect 399430 292046 399498 292102
rect 399554 292046 399622 292102
rect 399678 292046 399774 292102
rect 399154 291978 399774 292046
rect 399154 291922 399250 291978
rect 399306 291922 399374 291978
rect 399430 291922 399498 291978
rect 399554 291922 399622 291978
rect 399678 291922 399774 291978
rect 399154 274350 399774 291922
rect 399154 274294 399250 274350
rect 399306 274294 399374 274350
rect 399430 274294 399498 274350
rect 399554 274294 399622 274350
rect 399678 274294 399774 274350
rect 399154 274226 399774 274294
rect 399154 274170 399250 274226
rect 399306 274170 399374 274226
rect 399430 274170 399498 274226
rect 399554 274170 399622 274226
rect 399678 274170 399774 274226
rect 399154 274102 399774 274170
rect 399154 274046 399250 274102
rect 399306 274046 399374 274102
rect 399430 274046 399498 274102
rect 399554 274046 399622 274102
rect 399678 274046 399774 274102
rect 399154 273978 399774 274046
rect 399154 273922 399250 273978
rect 399306 273922 399374 273978
rect 399430 273922 399498 273978
rect 399554 273922 399622 273978
rect 399678 273922 399774 273978
rect 399154 256350 399774 273922
rect 399154 256294 399250 256350
rect 399306 256294 399374 256350
rect 399430 256294 399498 256350
rect 399554 256294 399622 256350
rect 399678 256294 399774 256350
rect 399154 256226 399774 256294
rect 399154 256170 399250 256226
rect 399306 256170 399374 256226
rect 399430 256170 399498 256226
rect 399554 256170 399622 256226
rect 399678 256170 399774 256226
rect 399154 256102 399774 256170
rect 399154 256046 399250 256102
rect 399306 256046 399374 256102
rect 399430 256046 399498 256102
rect 399554 256046 399622 256102
rect 399678 256046 399774 256102
rect 399154 255978 399774 256046
rect 399154 255922 399250 255978
rect 399306 255922 399374 255978
rect 399430 255922 399498 255978
rect 399554 255922 399622 255978
rect 399678 255922 399774 255978
rect 399154 238350 399774 255922
rect 399154 238294 399250 238350
rect 399306 238294 399374 238350
rect 399430 238294 399498 238350
rect 399554 238294 399622 238350
rect 399678 238294 399774 238350
rect 399154 238226 399774 238294
rect 399154 238170 399250 238226
rect 399306 238170 399374 238226
rect 399430 238170 399498 238226
rect 399554 238170 399622 238226
rect 399678 238170 399774 238226
rect 399154 238102 399774 238170
rect 399154 238046 399250 238102
rect 399306 238046 399374 238102
rect 399430 238046 399498 238102
rect 399554 238046 399622 238102
rect 399678 238046 399774 238102
rect 399154 237978 399774 238046
rect 399154 237922 399250 237978
rect 399306 237922 399374 237978
rect 399430 237922 399498 237978
rect 399554 237922 399622 237978
rect 399678 237922 399774 237978
rect 399154 220350 399774 237922
rect 399154 220294 399250 220350
rect 399306 220294 399374 220350
rect 399430 220294 399498 220350
rect 399554 220294 399622 220350
rect 399678 220294 399774 220350
rect 399154 220226 399774 220294
rect 399154 220170 399250 220226
rect 399306 220170 399374 220226
rect 399430 220170 399498 220226
rect 399554 220170 399622 220226
rect 399678 220170 399774 220226
rect 399154 220102 399774 220170
rect 399154 220046 399250 220102
rect 399306 220046 399374 220102
rect 399430 220046 399498 220102
rect 399554 220046 399622 220102
rect 399678 220046 399774 220102
rect 399154 219978 399774 220046
rect 399154 219922 399250 219978
rect 399306 219922 399374 219978
rect 399430 219922 399498 219978
rect 399554 219922 399622 219978
rect 399678 219922 399774 219978
rect 399154 202350 399774 219922
rect 399154 202294 399250 202350
rect 399306 202294 399374 202350
rect 399430 202294 399498 202350
rect 399554 202294 399622 202350
rect 399678 202294 399774 202350
rect 399154 202226 399774 202294
rect 399154 202170 399250 202226
rect 399306 202170 399374 202226
rect 399430 202170 399498 202226
rect 399554 202170 399622 202226
rect 399678 202170 399774 202226
rect 399154 202102 399774 202170
rect 399154 202046 399250 202102
rect 399306 202046 399374 202102
rect 399430 202046 399498 202102
rect 399554 202046 399622 202102
rect 399678 202046 399774 202102
rect 399154 201978 399774 202046
rect 399154 201922 399250 201978
rect 399306 201922 399374 201978
rect 399430 201922 399498 201978
rect 399554 201922 399622 201978
rect 399678 201922 399774 201978
rect 399154 184350 399774 201922
rect 399154 184294 399250 184350
rect 399306 184294 399374 184350
rect 399430 184294 399498 184350
rect 399554 184294 399622 184350
rect 399678 184294 399774 184350
rect 399154 184226 399774 184294
rect 399154 184170 399250 184226
rect 399306 184170 399374 184226
rect 399430 184170 399498 184226
rect 399554 184170 399622 184226
rect 399678 184170 399774 184226
rect 399154 184102 399774 184170
rect 399154 184046 399250 184102
rect 399306 184046 399374 184102
rect 399430 184046 399498 184102
rect 399554 184046 399622 184102
rect 399678 184046 399774 184102
rect 399154 183978 399774 184046
rect 399154 183922 399250 183978
rect 399306 183922 399374 183978
rect 399430 183922 399498 183978
rect 399554 183922 399622 183978
rect 399678 183922 399774 183978
rect 399154 166350 399774 183922
rect 399154 166294 399250 166350
rect 399306 166294 399374 166350
rect 399430 166294 399498 166350
rect 399554 166294 399622 166350
rect 399678 166294 399774 166350
rect 399154 166226 399774 166294
rect 399154 166170 399250 166226
rect 399306 166170 399374 166226
rect 399430 166170 399498 166226
rect 399554 166170 399622 166226
rect 399678 166170 399774 166226
rect 399154 166102 399774 166170
rect 399154 166046 399250 166102
rect 399306 166046 399374 166102
rect 399430 166046 399498 166102
rect 399554 166046 399622 166102
rect 399678 166046 399774 166102
rect 399154 165978 399774 166046
rect 399154 165922 399250 165978
rect 399306 165922 399374 165978
rect 399430 165922 399498 165978
rect 399554 165922 399622 165978
rect 399678 165922 399774 165978
rect 384874 154294 384970 154350
rect 385026 154294 385094 154350
rect 385150 154294 385218 154350
rect 385274 154294 385342 154350
rect 385398 154294 385494 154350
rect 384874 154226 385494 154294
rect 384874 154170 384970 154226
rect 385026 154170 385094 154226
rect 385150 154170 385218 154226
rect 385274 154170 385342 154226
rect 385398 154170 385494 154226
rect 384874 154102 385494 154170
rect 384874 154046 384970 154102
rect 385026 154046 385094 154102
rect 385150 154046 385218 154102
rect 385274 154046 385342 154102
rect 385398 154046 385494 154102
rect 384874 153978 385494 154046
rect 384874 153922 384970 153978
rect 385026 153922 385094 153978
rect 385150 153922 385218 153978
rect 385274 153922 385342 153978
rect 385398 153922 385494 153978
rect 384874 136350 385494 153922
rect 384874 136294 384970 136350
rect 385026 136294 385094 136350
rect 385150 136294 385218 136350
rect 385274 136294 385342 136350
rect 385398 136294 385494 136350
rect 384874 136226 385494 136294
rect 384874 136170 384970 136226
rect 385026 136170 385094 136226
rect 385150 136170 385218 136226
rect 385274 136170 385342 136226
rect 385398 136170 385494 136226
rect 384874 136102 385494 136170
rect 384874 136046 384970 136102
rect 385026 136046 385094 136102
rect 385150 136046 385218 136102
rect 385274 136046 385342 136102
rect 385398 136046 385494 136102
rect 384874 135978 385494 136046
rect 384874 135922 384970 135978
rect 385026 135922 385094 135978
rect 385150 135922 385218 135978
rect 385274 135922 385342 135978
rect 385398 135922 385494 135978
rect 384874 118350 385494 135922
rect 384874 118294 384970 118350
rect 385026 118294 385094 118350
rect 385150 118294 385218 118350
rect 385274 118294 385342 118350
rect 385398 118294 385494 118350
rect 384874 118226 385494 118294
rect 384874 118170 384970 118226
rect 385026 118170 385094 118226
rect 385150 118170 385218 118226
rect 385274 118170 385342 118226
rect 385398 118170 385494 118226
rect 384874 118102 385494 118170
rect 384874 118046 384970 118102
rect 385026 118046 385094 118102
rect 385150 118046 385218 118102
rect 385274 118046 385342 118102
rect 385398 118046 385494 118102
rect 384874 117978 385494 118046
rect 384874 117922 384970 117978
rect 385026 117922 385094 117978
rect 385150 117922 385218 117978
rect 385274 117922 385342 117978
rect 385398 117922 385494 117978
rect 384874 100350 385494 117922
rect 384874 100294 384970 100350
rect 385026 100294 385094 100350
rect 385150 100294 385218 100350
rect 385274 100294 385342 100350
rect 385398 100294 385494 100350
rect 384874 100226 385494 100294
rect 384874 100170 384970 100226
rect 385026 100170 385094 100226
rect 385150 100170 385218 100226
rect 385274 100170 385342 100226
rect 385398 100170 385494 100226
rect 384874 100102 385494 100170
rect 384874 100046 384970 100102
rect 385026 100046 385094 100102
rect 385150 100046 385218 100102
rect 385274 100046 385342 100102
rect 385398 100046 385494 100102
rect 384874 99978 385494 100046
rect 384874 99922 384970 99978
rect 385026 99922 385094 99978
rect 385150 99922 385218 99978
rect 385274 99922 385342 99978
rect 385398 99922 385494 99978
rect 384874 82350 385494 99922
rect 384874 82294 384970 82350
rect 385026 82294 385094 82350
rect 385150 82294 385218 82350
rect 385274 82294 385342 82350
rect 385398 82294 385494 82350
rect 384874 82226 385494 82294
rect 384874 82170 384970 82226
rect 385026 82170 385094 82226
rect 385150 82170 385218 82226
rect 385274 82170 385342 82226
rect 385398 82170 385494 82226
rect 384874 82102 385494 82170
rect 384874 82046 384970 82102
rect 385026 82046 385094 82102
rect 385150 82046 385218 82102
rect 385274 82046 385342 82102
rect 385398 82046 385494 82102
rect 384874 81978 385494 82046
rect 384874 81922 384970 81978
rect 385026 81922 385094 81978
rect 385150 81922 385218 81978
rect 385274 81922 385342 81978
rect 385398 81922 385494 81978
rect 384874 64350 385494 81922
rect 384874 64294 384970 64350
rect 385026 64294 385094 64350
rect 385150 64294 385218 64350
rect 385274 64294 385342 64350
rect 385398 64294 385494 64350
rect 384874 64226 385494 64294
rect 384874 64170 384970 64226
rect 385026 64170 385094 64226
rect 385150 64170 385218 64226
rect 385274 64170 385342 64226
rect 385398 64170 385494 64226
rect 384874 64102 385494 64170
rect 384874 64046 384970 64102
rect 385026 64046 385094 64102
rect 385150 64046 385218 64102
rect 385274 64046 385342 64102
rect 385398 64046 385494 64102
rect 384874 63978 385494 64046
rect 384874 63922 384970 63978
rect 385026 63922 385094 63978
rect 385150 63922 385218 63978
rect 385274 63922 385342 63978
rect 385398 63922 385494 63978
rect 384874 46350 385494 63922
rect 384874 46294 384970 46350
rect 385026 46294 385094 46350
rect 385150 46294 385218 46350
rect 385274 46294 385342 46350
rect 385398 46294 385494 46350
rect 384874 46226 385494 46294
rect 384874 46170 384970 46226
rect 385026 46170 385094 46226
rect 385150 46170 385218 46226
rect 385274 46170 385342 46226
rect 385398 46170 385494 46226
rect 384874 46102 385494 46170
rect 384874 46046 384970 46102
rect 385026 46046 385094 46102
rect 385150 46046 385218 46102
rect 385274 46046 385342 46102
rect 385398 46046 385494 46102
rect 384874 45978 385494 46046
rect 384874 45922 384970 45978
rect 385026 45922 385094 45978
rect 385150 45922 385218 45978
rect 385274 45922 385342 45978
rect 385398 45922 385494 45978
rect 384874 28350 385494 45922
rect 384874 28294 384970 28350
rect 385026 28294 385094 28350
rect 385150 28294 385218 28350
rect 385274 28294 385342 28350
rect 385398 28294 385494 28350
rect 384874 28226 385494 28294
rect 384874 28170 384970 28226
rect 385026 28170 385094 28226
rect 385150 28170 385218 28226
rect 385274 28170 385342 28226
rect 385398 28170 385494 28226
rect 384874 28102 385494 28170
rect 384874 28046 384970 28102
rect 385026 28046 385094 28102
rect 385150 28046 385218 28102
rect 385274 28046 385342 28102
rect 385398 28046 385494 28102
rect 384874 27978 385494 28046
rect 384874 27922 384970 27978
rect 385026 27922 385094 27978
rect 385150 27922 385218 27978
rect 385274 27922 385342 27978
rect 385398 27922 385494 27978
rect 384874 10350 385494 27922
rect 384874 10294 384970 10350
rect 385026 10294 385094 10350
rect 385150 10294 385218 10350
rect 385274 10294 385342 10350
rect 385398 10294 385494 10350
rect 384874 10226 385494 10294
rect 384874 10170 384970 10226
rect 385026 10170 385094 10226
rect 385150 10170 385218 10226
rect 385274 10170 385342 10226
rect 385398 10170 385494 10226
rect 384874 10102 385494 10170
rect 384874 10046 384970 10102
rect 385026 10046 385094 10102
rect 385150 10046 385218 10102
rect 385274 10046 385342 10102
rect 385398 10046 385494 10102
rect 384874 9978 385494 10046
rect 384874 9922 384970 9978
rect 385026 9922 385094 9978
rect 385150 9922 385218 9978
rect 385274 9922 385342 9978
rect 385398 9922 385494 9978
rect 384874 -1120 385494 9922
rect 384874 -1176 384970 -1120
rect 385026 -1176 385094 -1120
rect 385150 -1176 385218 -1120
rect 385274 -1176 385342 -1120
rect 385398 -1176 385494 -1120
rect 384874 -1244 385494 -1176
rect 384874 -1300 384970 -1244
rect 385026 -1300 385094 -1244
rect 385150 -1300 385218 -1244
rect 385274 -1300 385342 -1244
rect 385398 -1300 385494 -1244
rect 384874 -1368 385494 -1300
rect 384874 -1424 384970 -1368
rect 385026 -1424 385094 -1368
rect 385150 -1424 385218 -1368
rect 385274 -1424 385342 -1368
rect 385398 -1424 385494 -1368
rect 384874 -1492 385494 -1424
rect 384874 -1548 384970 -1492
rect 385026 -1548 385094 -1492
rect 385150 -1548 385218 -1492
rect 385274 -1548 385342 -1492
rect 385398 -1548 385494 -1492
rect 384874 -1644 385494 -1548
rect 399154 148350 399774 165922
rect 399154 148294 399250 148350
rect 399306 148294 399374 148350
rect 399430 148294 399498 148350
rect 399554 148294 399622 148350
rect 399678 148294 399774 148350
rect 399154 148226 399774 148294
rect 399154 148170 399250 148226
rect 399306 148170 399374 148226
rect 399430 148170 399498 148226
rect 399554 148170 399622 148226
rect 399678 148170 399774 148226
rect 399154 148102 399774 148170
rect 399154 148046 399250 148102
rect 399306 148046 399374 148102
rect 399430 148046 399498 148102
rect 399554 148046 399622 148102
rect 399678 148046 399774 148102
rect 399154 147978 399774 148046
rect 399154 147922 399250 147978
rect 399306 147922 399374 147978
rect 399430 147922 399498 147978
rect 399554 147922 399622 147978
rect 399678 147922 399774 147978
rect 399154 130350 399774 147922
rect 399154 130294 399250 130350
rect 399306 130294 399374 130350
rect 399430 130294 399498 130350
rect 399554 130294 399622 130350
rect 399678 130294 399774 130350
rect 399154 130226 399774 130294
rect 399154 130170 399250 130226
rect 399306 130170 399374 130226
rect 399430 130170 399498 130226
rect 399554 130170 399622 130226
rect 399678 130170 399774 130226
rect 399154 130102 399774 130170
rect 399154 130046 399250 130102
rect 399306 130046 399374 130102
rect 399430 130046 399498 130102
rect 399554 130046 399622 130102
rect 399678 130046 399774 130102
rect 399154 129978 399774 130046
rect 399154 129922 399250 129978
rect 399306 129922 399374 129978
rect 399430 129922 399498 129978
rect 399554 129922 399622 129978
rect 399678 129922 399774 129978
rect 399154 112350 399774 129922
rect 399154 112294 399250 112350
rect 399306 112294 399374 112350
rect 399430 112294 399498 112350
rect 399554 112294 399622 112350
rect 399678 112294 399774 112350
rect 399154 112226 399774 112294
rect 399154 112170 399250 112226
rect 399306 112170 399374 112226
rect 399430 112170 399498 112226
rect 399554 112170 399622 112226
rect 399678 112170 399774 112226
rect 399154 112102 399774 112170
rect 399154 112046 399250 112102
rect 399306 112046 399374 112102
rect 399430 112046 399498 112102
rect 399554 112046 399622 112102
rect 399678 112046 399774 112102
rect 399154 111978 399774 112046
rect 399154 111922 399250 111978
rect 399306 111922 399374 111978
rect 399430 111922 399498 111978
rect 399554 111922 399622 111978
rect 399678 111922 399774 111978
rect 399154 94350 399774 111922
rect 399154 94294 399250 94350
rect 399306 94294 399374 94350
rect 399430 94294 399498 94350
rect 399554 94294 399622 94350
rect 399678 94294 399774 94350
rect 399154 94226 399774 94294
rect 399154 94170 399250 94226
rect 399306 94170 399374 94226
rect 399430 94170 399498 94226
rect 399554 94170 399622 94226
rect 399678 94170 399774 94226
rect 399154 94102 399774 94170
rect 399154 94046 399250 94102
rect 399306 94046 399374 94102
rect 399430 94046 399498 94102
rect 399554 94046 399622 94102
rect 399678 94046 399774 94102
rect 399154 93978 399774 94046
rect 399154 93922 399250 93978
rect 399306 93922 399374 93978
rect 399430 93922 399498 93978
rect 399554 93922 399622 93978
rect 399678 93922 399774 93978
rect 399154 76350 399774 93922
rect 399154 76294 399250 76350
rect 399306 76294 399374 76350
rect 399430 76294 399498 76350
rect 399554 76294 399622 76350
rect 399678 76294 399774 76350
rect 399154 76226 399774 76294
rect 399154 76170 399250 76226
rect 399306 76170 399374 76226
rect 399430 76170 399498 76226
rect 399554 76170 399622 76226
rect 399678 76170 399774 76226
rect 399154 76102 399774 76170
rect 399154 76046 399250 76102
rect 399306 76046 399374 76102
rect 399430 76046 399498 76102
rect 399554 76046 399622 76102
rect 399678 76046 399774 76102
rect 399154 75978 399774 76046
rect 399154 75922 399250 75978
rect 399306 75922 399374 75978
rect 399430 75922 399498 75978
rect 399554 75922 399622 75978
rect 399678 75922 399774 75978
rect 399154 58350 399774 75922
rect 399154 58294 399250 58350
rect 399306 58294 399374 58350
rect 399430 58294 399498 58350
rect 399554 58294 399622 58350
rect 399678 58294 399774 58350
rect 399154 58226 399774 58294
rect 399154 58170 399250 58226
rect 399306 58170 399374 58226
rect 399430 58170 399498 58226
rect 399554 58170 399622 58226
rect 399678 58170 399774 58226
rect 399154 58102 399774 58170
rect 399154 58046 399250 58102
rect 399306 58046 399374 58102
rect 399430 58046 399498 58102
rect 399554 58046 399622 58102
rect 399678 58046 399774 58102
rect 399154 57978 399774 58046
rect 399154 57922 399250 57978
rect 399306 57922 399374 57978
rect 399430 57922 399498 57978
rect 399554 57922 399622 57978
rect 399678 57922 399774 57978
rect 399154 40350 399774 57922
rect 399154 40294 399250 40350
rect 399306 40294 399374 40350
rect 399430 40294 399498 40350
rect 399554 40294 399622 40350
rect 399678 40294 399774 40350
rect 399154 40226 399774 40294
rect 399154 40170 399250 40226
rect 399306 40170 399374 40226
rect 399430 40170 399498 40226
rect 399554 40170 399622 40226
rect 399678 40170 399774 40226
rect 399154 40102 399774 40170
rect 399154 40046 399250 40102
rect 399306 40046 399374 40102
rect 399430 40046 399498 40102
rect 399554 40046 399622 40102
rect 399678 40046 399774 40102
rect 399154 39978 399774 40046
rect 399154 39922 399250 39978
rect 399306 39922 399374 39978
rect 399430 39922 399498 39978
rect 399554 39922 399622 39978
rect 399678 39922 399774 39978
rect 399154 22350 399774 39922
rect 399154 22294 399250 22350
rect 399306 22294 399374 22350
rect 399430 22294 399498 22350
rect 399554 22294 399622 22350
rect 399678 22294 399774 22350
rect 399154 22226 399774 22294
rect 399154 22170 399250 22226
rect 399306 22170 399374 22226
rect 399430 22170 399498 22226
rect 399554 22170 399622 22226
rect 399678 22170 399774 22226
rect 399154 22102 399774 22170
rect 399154 22046 399250 22102
rect 399306 22046 399374 22102
rect 399430 22046 399498 22102
rect 399554 22046 399622 22102
rect 399678 22046 399774 22102
rect 399154 21978 399774 22046
rect 399154 21922 399250 21978
rect 399306 21922 399374 21978
rect 399430 21922 399498 21978
rect 399554 21922 399622 21978
rect 399678 21922 399774 21978
rect 399154 4350 399774 21922
rect 399154 4294 399250 4350
rect 399306 4294 399374 4350
rect 399430 4294 399498 4350
rect 399554 4294 399622 4350
rect 399678 4294 399774 4350
rect 399154 4226 399774 4294
rect 399154 4170 399250 4226
rect 399306 4170 399374 4226
rect 399430 4170 399498 4226
rect 399554 4170 399622 4226
rect 399678 4170 399774 4226
rect 399154 4102 399774 4170
rect 399154 4046 399250 4102
rect 399306 4046 399374 4102
rect 399430 4046 399498 4102
rect 399554 4046 399622 4102
rect 399678 4046 399774 4102
rect 399154 3978 399774 4046
rect 399154 3922 399250 3978
rect 399306 3922 399374 3978
rect 399430 3922 399498 3978
rect 399554 3922 399622 3978
rect 399678 3922 399774 3978
rect 399154 -160 399774 3922
rect 399154 -216 399250 -160
rect 399306 -216 399374 -160
rect 399430 -216 399498 -160
rect 399554 -216 399622 -160
rect 399678 -216 399774 -160
rect 399154 -284 399774 -216
rect 399154 -340 399250 -284
rect 399306 -340 399374 -284
rect 399430 -340 399498 -284
rect 399554 -340 399622 -284
rect 399678 -340 399774 -284
rect 399154 -408 399774 -340
rect 399154 -464 399250 -408
rect 399306 -464 399374 -408
rect 399430 -464 399498 -408
rect 399554 -464 399622 -408
rect 399678 -464 399774 -408
rect 399154 -532 399774 -464
rect 399154 -588 399250 -532
rect 399306 -588 399374 -532
rect 399430 -588 399498 -532
rect 399554 -588 399622 -532
rect 399678 -588 399774 -532
rect 399154 -1644 399774 -588
rect 402874 598172 403494 598268
rect 402874 598116 402970 598172
rect 403026 598116 403094 598172
rect 403150 598116 403218 598172
rect 403274 598116 403342 598172
rect 403398 598116 403494 598172
rect 402874 598048 403494 598116
rect 402874 597992 402970 598048
rect 403026 597992 403094 598048
rect 403150 597992 403218 598048
rect 403274 597992 403342 598048
rect 403398 597992 403494 598048
rect 402874 597924 403494 597992
rect 402874 597868 402970 597924
rect 403026 597868 403094 597924
rect 403150 597868 403218 597924
rect 403274 597868 403342 597924
rect 403398 597868 403494 597924
rect 402874 597800 403494 597868
rect 402874 597744 402970 597800
rect 403026 597744 403094 597800
rect 403150 597744 403218 597800
rect 403274 597744 403342 597800
rect 403398 597744 403494 597800
rect 402874 586350 403494 597744
rect 402874 586294 402970 586350
rect 403026 586294 403094 586350
rect 403150 586294 403218 586350
rect 403274 586294 403342 586350
rect 403398 586294 403494 586350
rect 402874 586226 403494 586294
rect 402874 586170 402970 586226
rect 403026 586170 403094 586226
rect 403150 586170 403218 586226
rect 403274 586170 403342 586226
rect 403398 586170 403494 586226
rect 402874 586102 403494 586170
rect 402874 586046 402970 586102
rect 403026 586046 403094 586102
rect 403150 586046 403218 586102
rect 403274 586046 403342 586102
rect 403398 586046 403494 586102
rect 402874 585978 403494 586046
rect 402874 585922 402970 585978
rect 403026 585922 403094 585978
rect 403150 585922 403218 585978
rect 403274 585922 403342 585978
rect 403398 585922 403494 585978
rect 402874 568350 403494 585922
rect 402874 568294 402970 568350
rect 403026 568294 403094 568350
rect 403150 568294 403218 568350
rect 403274 568294 403342 568350
rect 403398 568294 403494 568350
rect 402874 568226 403494 568294
rect 402874 568170 402970 568226
rect 403026 568170 403094 568226
rect 403150 568170 403218 568226
rect 403274 568170 403342 568226
rect 403398 568170 403494 568226
rect 402874 568102 403494 568170
rect 402874 568046 402970 568102
rect 403026 568046 403094 568102
rect 403150 568046 403218 568102
rect 403274 568046 403342 568102
rect 403398 568046 403494 568102
rect 402874 567978 403494 568046
rect 402874 567922 402970 567978
rect 403026 567922 403094 567978
rect 403150 567922 403218 567978
rect 403274 567922 403342 567978
rect 403398 567922 403494 567978
rect 402874 550350 403494 567922
rect 402874 550294 402970 550350
rect 403026 550294 403094 550350
rect 403150 550294 403218 550350
rect 403274 550294 403342 550350
rect 403398 550294 403494 550350
rect 402874 550226 403494 550294
rect 402874 550170 402970 550226
rect 403026 550170 403094 550226
rect 403150 550170 403218 550226
rect 403274 550170 403342 550226
rect 403398 550170 403494 550226
rect 402874 550102 403494 550170
rect 402874 550046 402970 550102
rect 403026 550046 403094 550102
rect 403150 550046 403218 550102
rect 403274 550046 403342 550102
rect 403398 550046 403494 550102
rect 402874 549978 403494 550046
rect 402874 549922 402970 549978
rect 403026 549922 403094 549978
rect 403150 549922 403218 549978
rect 403274 549922 403342 549978
rect 403398 549922 403494 549978
rect 402874 532350 403494 549922
rect 402874 532294 402970 532350
rect 403026 532294 403094 532350
rect 403150 532294 403218 532350
rect 403274 532294 403342 532350
rect 403398 532294 403494 532350
rect 402874 532226 403494 532294
rect 402874 532170 402970 532226
rect 403026 532170 403094 532226
rect 403150 532170 403218 532226
rect 403274 532170 403342 532226
rect 403398 532170 403494 532226
rect 402874 532102 403494 532170
rect 402874 532046 402970 532102
rect 403026 532046 403094 532102
rect 403150 532046 403218 532102
rect 403274 532046 403342 532102
rect 403398 532046 403494 532102
rect 402874 531978 403494 532046
rect 402874 531922 402970 531978
rect 403026 531922 403094 531978
rect 403150 531922 403218 531978
rect 403274 531922 403342 531978
rect 403398 531922 403494 531978
rect 402874 514350 403494 531922
rect 402874 514294 402970 514350
rect 403026 514294 403094 514350
rect 403150 514294 403218 514350
rect 403274 514294 403342 514350
rect 403398 514294 403494 514350
rect 402874 514226 403494 514294
rect 402874 514170 402970 514226
rect 403026 514170 403094 514226
rect 403150 514170 403218 514226
rect 403274 514170 403342 514226
rect 403398 514170 403494 514226
rect 402874 514102 403494 514170
rect 402874 514046 402970 514102
rect 403026 514046 403094 514102
rect 403150 514046 403218 514102
rect 403274 514046 403342 514102
rect 403398 514046 403494 514102
rect 402874 513978 403494 514046
rect 402874 513922 402970 513978
rect 403026 513922 403094 513978
rect 403150 513922 403218 513978
rect 403274 513922 403342 513978
rect 403398 513922 403494 513978
rect 402874 496350 403494 513922
rect 402874 496294 402970 496350
rect 403026 496294 403094 496350
rect 403150 496294 403218 496350
rect 403274 496294 403342 496350
rect 403398 496294 403494 496350
rect 402874 496226 403494 496294
rect 402874 496170 402970 496226
rect 403026 496170 403094 496226
rect 403150 496170 403218 496226
rect 403274 496170 403342 496226
rect 403398 496170 403494 496226
rect 402874 496102 403494 496170
rect 402874 496046 402970 496102
rect 403026 496046 403094 496102
rect 403150 496046 403218 496102
rect 403274 496046 403342 496102
rect 403398 496046 403494 496102
rect 402874 495978 403494 496046
rect 402874 495922 402970 495978
rect 403026 495922 403094 495978
rect 403150 495922 403218 495978
rect 403274 495922 403342 495978
rect 403398 495922 403494 495978
rect 402874 478350 403494 495922
rect 402874 478294 402970 478350
rect 403026 478294 403094 478350
rect 403150 478294 403218 478350
rect 403274 478294 403342 478350
rect 403398 478294 403494 478350
rect 402874 478226 403494 478294
rect 402874 478170 402970 478226
rect 403026 478170 403094 478226
rect 403150 478170 403218 478226
rect 403274 478170 403342 478226
rect 403398 478170 403494 478226
rect 402874 478102 403494 478170
rect 402874 478046 402970 478102
rect 403026 478046 403094 478102
rect 403150 478046 403218 478102
rect 403274 478046 403342 478102
rect 403398 478046 403494 478102
rect 402874 477978 403494 478046
rect 402874 477922 402970 477978
rect 403026 477922 403094 477978
rect 403150 477922 403218 477978
rect 403274 477922 403342 477978
rect 403398 477922 403494 477978
rect 402874 460350 403494 477922
rect 402874 460294 402970 460350
rect 403026 460294 403094 460350
rect 403150 460294 403218 460350
rect 403274 460294 403342 460350
rect 403398 460294 403494 460350
rect 402874 460226 403494 460294
rect 402874 460170 402970 460226
rect 403026 460170 403094 460226
rect 403150 460170 403218 460226
rect 403274 460170 403342 460226
rect 403398 460170 403494 460226
rect 402874 460102 403494 460170
rect 402874 460046 402970 460102
rect 403026 460046 403094 460102
rect 403150 460046 403218 460102
rect 403274 460046 403342 460102
rect 403398 460046 403494 460102
rect 402874 459978 403494 460046
rect 402874 459922 402970 459978
rect 403026 459922 403094 459978
rect 403150 459922 403218 459978
rect 403274 459922 403342 459978
rect 403398 459922 403494 459978
rect 402874 442350 403494 459922
rect 417154 597212 417774 598268
rect 417154 597156 417250 597212
rect 417306 597156 417374 597212
rect 417430 597156 417498 597212
rect 417554 597156 417622 597212
rect 417678 597156 417774 597212
rect 417154 597088 417774 597156
rect 417154 597032 417250 597088
rect 417306 597032 417374 597088
rect 417430 597032 417498 597088
rect 417554 597032 417622 597088
rect 417678 597032 417774 597088
rect 417154 596964 417774 597032
rect 417154 596908 417250 596964
rect 417306 596908 417374 596964
rect 417430 596908 417498 596964
rect 417554 596908 417622 596964
rect 417678 596908 417774 596964
rect 417154 596840 417774 596908
rect 417154 596784 417250 596840
rect 417306 596784 417374 596840
rect 417430 596784 417498 596840
rect 417554 596784 417622 596840
rect 417678 596784 417774 596840
rect 417154 580350 417774 596784
rect 417154 580294 417250 580350
rect 417306 580294 417374 580350
rect 417430 580294 417498 580350
rect 417554 580294 417622 580350
rect 417678 580294 417774 580350
rect 417154 580226 417774 580294
rect 417154 580170 417250 580226
rect 417306 580170 417374 580226
rect 417430 580170 417498 580226
rect 417554 580170 417622 580226
rect 417678 580170 417774 580226
rect 417154 580102 417774 580170
rect 417154 580046 417250 580102
rect 417306 580046 417374 580102
rect 417430 580046 417498 580102
rect 417554 580046 417622 580102
rect 417678 580046 417774 580102
rect 417154 579978 417774 580046
rect 417154 579922 417250 579978
rect 417306 579922 417374 579978
rect 417430 579922 417498 579978
rect 417554 579922 417622 579978
rect 417678 579922 417774 579978
rect 417154 562350 417774 579922
rect 417154 562294 417250 562350
rect 417306 562294 417374 562350
rect 417430 562294 417498 562350
rect 417554 562294 417622 562350
rect 417678 562294 417774 562350
rect 417154 562226 417774 562294
rect 417154 562170 417250 562226
rect 417306 562170 417374 562226
rect 417430 562170 417498 562226
rect 417554 562170 417622 562226
rect 417678 562170 417774 562226
rect 417154 562102 417774 562170
rect 417154 562046 417250 562102
rect 417306 562046 417374 562102
rect 417430 562046 417498 562102
rect 417554 562046 417622 562102
rect 417678 562046 417774 562102
rect 417154 561978 417774 562046
rect 417154 561922 417250 561978
rect 417306 561922 417374 561978
rect 417430 561922 417498 561978
rect 417554 561922 417622 561978
rect 417678 561922 417774 561978
rect 417154 544350 417774 561922
rect 417154 544294 417250 544350
rect 417306 544294 417374 544350
rect 417430 544294 417498 544350
rect 417554 544294 417622 544350
rect 417678 544294 417774 544350
rect 417154 544226 417774 544294
rect 417154 544170 417250 544226
rect 417306 544170 417374 544226
rect 417430 544170 417498 544226
rect 417554 544170 417622 544226
rect 417678 544170 417774 544226
rect 417154 544102 417774 544170
rect 417154 544046 417250 544102
rect 417306 544046 417374 544102
rect 417430 544046 417498 544102
rect 417554 544046 417622 544102
rect 417678 544046 417774 544102
rect 417154 543978 417774 544046
rect 417154 543922 417250 543978
rect 417306 543922 417374 543978
rect 417430 543922 417498 543978
rect 417554 543922 417622 543978
rect 417678 543922 417774 543978
rect 417154 526350 417774 543922
rect 417154 526294 417250 526350
rect 417306 526294 417374 526350
rect 417430 526294 417498 526350
rect 417554 526294 417622 526350
rect 417678 526294 417774 526350
rect 417154 526226 417774 526294
rect 417154 526170 417250 526226
rect 417306 526170 417374 526226
rect 417430 526170 417498 526226
rect 417554 526170 417622 526226
rect 417678 526170 417774 526226
rect 417154 526102 417774 526170
rect 417154 526046 417250 526102
rect 417306 526046 417374 526102
rect 417430 526046 417498 526102
rect 417554 526046 417622 526102
rect 417678 526046 417774 526102
rect 417154 525978 417774 526046
rect 417154 525922 417250 525978
rect 417306 525922 417374 525978
rect 417430 525922 417498 525978
rect 417554 525922 417622 525978
rect 417678 525922 417774 525978
rect 417154 508350 417774 525922
rect 417154 508294 417250 508350
rect 417306 508294 417374 508350
rect 417430 508294 417498 508350
rect 417554 508294 417622 508350
rect 417678 508294 417774 508350
rect 417154 508226 417774 508294
rect 417154 508170 417250 508226
rect 417306 508170 417374 508226
rect 417430 508170 417498 508226
rect 417554 508170 417622 508226
rect 417678 508170 417774 508226
rect 417154 508102 417774 508170
rect 417154 508046 417250 508102
rect 417306 508046 417374 508102
rect 417430 508046 417498 508102
rect 417554 508046 417622 508102
rect 417678 508046 417774 508102
rect 417154 507978 417774 508046
rect 417154 507922 417250 507978
rect 417306 507922 417374 507978
rect 417430 507922 417498 507978
rect 417554 507922 417622 507978
rect 417678 507922 417774 507978
rect 417154 490350 417774 507922
rect 417154 490294 417250 490350
rect 417306 490294 417374 490350
rect 417430 490294 417498 490350
rect 417554 490294 417622 490350
rect 417678 490294 417774 490350
rect 417154 490226 417774 490294
rect 417154 490170 417250 490226
rect 417306 490170 417374 490226
rect 417430 490170 417498 490226
rect 417554 490170 417622 490226
rect 417678 490170 417774 490226
rect 417154 490102 417774 490170
rect 417154 490046 417250 490102
rect 417306 490046 417374 490102
rect 417430 490046 417498 490102
rect 417554 490046 417622 490102
rect 417678 490046 417774 490102
rect 417154 489978 417774 490046
rect 417154 489922 417250 489978
rect 417306 489922 417374 489978
rect 417430 489922 417498 489978
rect 417554 489922 417622 489978
rect 417678 489922 417774 489978
rect 417154 472350 417774 489922
rect 417154 472294 417250 472350
rect 417306 472294 417374 472350
rect 417430 472294 417498 472350
rect 417554 472294 417622 472350
rect 417678 472294 417774 472350
rect 417154 472226 417774 472294
rect 417154 472170 417250 472226
rect 417306 472170 417374 472226
rect 417430 472170 417498 472226
rect 417554 472170 417622 472226
rect 417678 472170 417774 472226
rect 417154 472102 417774 472170
rect 417154 472046 417250 472102
rect 417306 472046 417374 472102
rect 417430 472046 417498 472102
rect 417554 472046 417622 472102
rect 417678 472046 417774 472102
rect 417154 471978 417774 472046
rect 417154 471922 417250 471978
rect 417306 471922 417374 471978
rect 417430 471922 417498 471978
rect 417554 471922 417622 471978
rect 417678 471922 417774 471978
rect 417154 458342 417774 471922
rect 420874 598172 421494 598268
rect 420874 598116 420970 598172
rect 421026 598116 421094 598172
rect 421150 598116 421218 598172
rect 421274 598116 421342 598172
rect 421398 598116 421494 598172
rect 420874 598048 421494 598116
rect 420874 597992 420970 598048
rect 421026 597992 421094 598048
rect 421150 597992 421218 598048
rect 421274 597992 421342 598048
rect 421398 597992 421494 598048
rect 420874 597924 421494 597992
rect 420874 597868 420970 597924
rect 421026 597868 421094 597924
rect 421150 597868 421218 597924
rect 421274 597868 421342 597924
rect 421398 597868 421494 597924
rect 420874 597800 421494 597868
rect 420874 597744 420970 597800
rect 421026 597744 421094 597800
rect 421150 597744 421218 597800
rect 421274 597744 421342 597800
rect 421398 597744 421494 597800
rect 420874 586350 421494 597744
rect 420874 586294 420970 586350
rect 421026 586294 421094 586350
rect 421150 586294 421218 586350
rect 421274 586294 421342 586350
rect 421398 586294 421494 586350
rect 420874 586226 421494 586294
rect 420874 586170 420970 586226
rect 421026 586170 421094 586226
rect 421150 586170 421218 586226
rect 421274 586170 421342 586226
rect 421398 586170 421494 586226
rect 420874 586102 421494 586170
rect 420874 586046 420970 586102
rect 421026 586046 421094 586102
rect 421150 586046 421218 586102
rect 421274 586046 421342 586102
rect 421398 586046 421494 586102
rect 420874 585978 421494 586046
rect 420874 585922 420970 585978
rect 421026 585922 421094 585978
rect 421150 585922 421218 585978
rect 421274 585922 421342 585978
rect 421398 585922 421494 585978
rect 420874 568350 421494 585922
rect 420874 568294 420970 568350
rect 421026 568294 421094 568350
rect 421150 568294 421218 568350
rect 421274 568294 421342 568350
rect 421398 568294 421494 568350
rect 420874 568226 421494 568294
rect 420874 568170 420970 568226
rect 421026 568170 421094 568226
rect 421150 568170 421218 568226
rect 421274 568170 421342 568226
rect 421398 568170 421494 568226
rect 420874 568102 421494 568170
rect 420874 568046 420970 568102
rect 421026 568046 421094 568102
rect 421150 568046 421218 568102
rect 421274 568046 421342 568102
rect 421398 568046 421494 568102
rect 420874 567978 421494 568046
rect 420874 567922 420970 567978
rect 421026 567922 421094 567978
rect 421150 567922 421218 567978
rect 421274 567922 421342 567978
rect 421398 567922 421494 567978
rect 420874 550350 421494 567922
rect 420874 550294 420970 550350
rect 421026 550294 421094 550350
rect 421150 550294 421218 550350
rect 421274 550294 421342 550350
rect 421398 550294 421494 550350
rect 420874 550226 421494 550294
rect 420874 550170 420970 550226
rect 421026 550170 421094 550226
rect 421150 550170 421218 550226
rect 421274 550170 421342 550226
rect 421398 550170 421494 550226
rect 420874 550102 421494 550170
rect 420874 550046 420970 550102
rect 421026 550046 421094 550102
rect 421150 550046 421218 550102
rect 421274 550046 421342 550102
rect 421398 550046 421494 550102
rect 420874 549978 421494 550046
rect 420874 549922 420970 549978
rect 421026 549922 421094 549978
rect 421150 549922 421218 549978
rect 421274 549922 421342 549978
rect 421398 549922 421494 549978
rect 420874 532350 421494 549922
rect 420874 532294 420970 532350
rect 421026 532294 421094 532350
rect 421150 532294 421218 532350
rect 421274 532294 421342 532350
rect 421398 532294 421494 532350
rect 420874 532226 421494 532294
rect 420874 532170 420970 532226
rect 421026 532170 421094 532226
rect 421150 532170 421218 532226
rect 421274 532170 421342 532226
rect 421398 532170 421494 532226
rect 420874 532102 421494 532170
rect 420874 532046 420970 532102
rect 421026 532046 421094 532102
rect 421150 532046 421218 532102
rect 421274 532046 421342 532102
rect 421398 532046 421494 532102
rect 420874 531978 421494 532046
rect 420874 531922 420970 531978
rect 421026 531922 421094 531978
rect 421150 531922 421218 531978
rect 421274 531922 421342 531978
rect 421398 531922 421494 531978
rect 420874 514350 421494 531922
rect 420874 514294 420970 514350
rect 421026 514294 421094 514350
rect 421150 514294 421218 514350
rect 421274 514294 421342 514350
rect 421398 514294 421494 514350
rect 420874 514226 421494 514294
rect 420874 514170 420970 514226
rect 421026 514170 421094 514226
rect 421150 514170 421218 514226
rect 421274 514170 421342 514226
rect 421398 514170 421494 514226
rect 420874 514102 421494 514170
rect 420874 514046 420970 514102
rect 421026 514046 421094 514102
rect 421150 514046 421218 514102
rect 421274 514046 421342 514102
rect 421398 514046 421494 514102
rect 420874 513978 421494 514046
rect 420874 513922 420970 513978
rect 421026 513922 421094 513978
rect 421150 513922 421218 513978
rect 421274 513922 421342 513978
rect 421398 513922 421494 513978
rect 420874 496350 421494 513922
rect 420874 496294 420970 496350
rect 421026 496294 421094 496350
rect 421150 496294 421218 496350
rect 421274 496294 421342 496350
rect 421398 496294 421494 496350
rect 420874 496226 421494 496294
rect 420874 496170 420970 496226
rect 421026 496170 421094 496226
rect 421150 496170 421218 496226
rect 421274 496170 421342 496226
rect 421398 496170 421494 496226
rect 420874 496102 421494 496170
rect 420874 496046 420970 496102
rect 421026 496046 421094 496102
rect 421150 496046 421218 496102
rect 421274 496046 421342 496102
rect 421398 496046 421494 496102
rect 420874 495978 421494 496046
rect 420874 495922 420970 495978
rect 421026 495922 421094 495978
rect 421150 495922 421218 495978
rect 421274 495922 421342 495978
rect 421398 495922 421494 495978
rect 420874 478350 421494 495922
rect 420874 478294 420970 478350
rect 421026 478294 421094 478350
rect 421150 478294 421218 478350
rect 421274 478294 421342 478350
rect 421398 478294 421494 478350
rect 420874 478226 421494 478294
rect 420874 478170 420970 478226
rect 421026 478170 421094 478226
rect 421150 478170 421218 478226
rect 421274 478170 421342 478226
rect 421398 478170 421494 478226
rect 420874 478102 421494 478170
rect 420874 478046 420970 478102
rect 421026 478046 421094 478102
rect 421150 478046 421218 478102
rect 421274 478046 421342 478102
rect 421398 478046 421494 478102
rect 420874 477978 421494 478046
rect 420874 477922 420970 477978
rect 421026 477922 421094 477978
rect 421150 477922 421218 477978
rect 421274 477922 421342 477978
rect 421398 477922 421494 477978
rect 420874 460350 421494 477922
rect 420874 460294 420970 460350
rect 421026 460294 421094 460350
rect 421150 460294 421218 460350
rect 421274 460294 421342 460350
rect 421398 460294 421494 460350
rect 420874 460226 421494 460294
rect 420874 460170 420970 460226
rect 421026 460170 421094 460226
rect 421150 460170 421218 460226
rect 421274 460170 421342 460226
rect 421398 460170 421494 460226
rect 420874 460102 421494 460170
rect 420874 460046 420970 460102
rect 421026 460046 421094 460102
rect 421150 460046 421218 460102
rect 421274 460046 421342 460102
rect 421398 460046 421494 460102
rect 420874 459978 421494 460046
rect 420874 459922 420970 459978
rect 421026 459922 421094 459978
rect 421150 459922 421218 459978
rect 421274 459922 421342 459978
rect 421398 459922 421494 459978
rect 420874 458342 421494 459922
rect 435154 597212 435774 598268
rect 435154 597156 435250 597212
rect 435306 597156 435374 597212
rect 435430 597156 435498 597212
rect 435554 597156 435622 597212
rect 435678 597156 435774 597212
rect 435154 597088 435774 597156
rect 435154 597032 435250 597088
rect 435306 597032 435374 597088
rect 435430 597032 435498 597088
rect 435554 597032 435622 597088
rect 435678 597032 435774 597088
rect 435154 596964 435774 597032
rect 435154 596908 435250 596964
rect 435306 596908 435374 596964
rect 435430 596908 435498 596964
rect 435554 596908 435622 596964
rect 435678 596908 435774 596964
rect 435154 596840 435774 596908
rect 435154 596784 435250 596840
rect 435306 596784 435374 596840
rect 435430 596784 435498 596840
rect 435554 596784 435622 596840
rect 435678 596784 435774 596840
rect 435154 580350 435774 596784
rect 435154 580294 435250 580350
rect 435306 580294 435374 580350
rect 435430 580294 435498 580350
rect 435554 580294 435622 580350
rect 435678 580294 435774 580350
rect 435154 580226 435774 580294
rect 435154 580170 435250 580226
rect 435306 580170 435374 580226
rect 435430 580170 435498 580226
rect 435554 580170 435622 580226
rect 435678 580170 435774 580226
rect 435154 580102 435774 580170
rect 435154 580046 435250 580102
rect 435306 580046 435374 580102
rect 435430 580046 435498 580102
rect 435554 580046 435622 580102
rect 435678 580046 435774 580102
rect 435154 579978 435774 580046
rect 435154 579922 435250 579978
rect 435306 579922 435374 579978
rect 435430 579922 435498 579978
rect 435554 579922 435622 579978
rect 435678 579922 435774 579978
rect 435154 562350 435774 579922
rect 435154 562294 435250 562350
rect 435306 562294 435374 562350
rect 435430 562294 435498 562350
rect 435554 562294 435622 562350
rect 435678 562294 435774 562350
rect 435154 562226 435774 562294
rect 435154 562170 435250 562226
rect 435306 562170 435374 562226
rect 435430 562170 435498 562226
rect 435554 562170 435622 562226
rect 435678 562170 435774 562226
rect 435154 562102 435774 562170
rect 435154 562046 435250 562102
rect 435306 562046 435374 562102
rect 435430 562046 435498 562102
rect 435554 562046 435622 562102
rect 435678 562046 435774 562102
rect 435154 561978 435774 562046
rect 435154 561922 435250 561978
rect 435306 561922 435374 561978
rect 435430 561922 435498 561978
rect 435554 561922 435622 561978
rect 435678 561922 435774 561978
rect 435154 544350 435774 561922
rect 435154 544294 435250 544350
rect 435306 544294 435374 544350
rect 435430 544294 435498 544350
rect 435554 544294 435622 544350
rect 435678 544294 435774 544350
rect 435154 544226 435774 544294
rect 435154 544170 435250 544226
rect 435306 544170 435374 544226
rect 435430 544170 435498 544226
rect 435554 544170 435622 544226
rect 435678 544170 435774 544226
rect 435154 544102 435774 544170
rect 435154 544046 435250 544102
rect 435306 544046 435374 544102
rect 435430 544046 435498 544102
rect 435554 544046 435622 544102
rect 435678 544046 435774 544102
rect 435154 543978 435774 544046
rect 435154 543922 435250 543978
rect 435306 543922 435374 543978
rect 435430 543922 435498 543978
rect 435554 543922 435622 543978
rect 435678 543922 435774 543978
rect 435154 526350 435774 543922
rect 435154 526294 435250 526350
rect 435306 526294 435374 526350
rect 435430 526294 435498 526350
rect 435554 526294 435622 526350
rect 435678 526294 435774 526350
rect 435154 526226 435774 526294
rect 435154 526170 435250 526226
rect 435306 526170 435374 526226
rect 435430 526170 435498 526226
rect 435554 526170 435622 526226
rect 435678 526170 435774 526226
rect 435154 526102 435774 526170
rect 435154 526046 435250 526102
rect 435306 526046 435374 526102
rect 435430 526046 435498 526102
rect 435554 526046 435622 526102
rect 435678 526046 435774 526102
rect 435154 525978 435774 526046
rect 435154 525922 435250 525978
rect 435306 525922 435374 525978
rect 435430 525922 435498 525978
rect 435554 525922 435622 525978
rect 435678 525922 435774 525978
rect 435154 508350 435774 525922
rect 435154 508294 435250 508350
rect 435306 508294 435374 508350
rect 435430 508294 435498 508350
rect 435554 508294 435622 508350
rect 435678 508294 435774 508350
rect 435154 508226 435774 508294
rect 435154 508170 435250 508226
rect 435306 508170 435374 508226
rect 435430 508170 435498 508226
rect 435554 508170 435622 508226
rect 435678 508170 435774 508226
rect 435154 508102 435774 508170
rect 435154 508046 435250 508102
rect 435306 508046 435374 508102
rect 435430 508046 435498 508102
rect 435554 508046 435622 508102
rect 435678 508046 435774 508102
rect 435154 507978 435774 508046
rect 435154 507922 435250 507978
rect 435306 507922 435374 507978
rect 435430 507922 435498 507978
rect 435554 507922 435622 507978
rect 435678 507922 435774 507978
rect 435154 490350 435774 507922
rect 435154 490294 435250 490350
rect 435306 490294 435374 490350
rect 435430 490294 435498 490350
rect 435554 490294 435622 490350
rect 435678 490294 435774 490350
rect 435154 490226 435774 490294
rect 435154 490170 435250 490226
rect 435306 490170 435374 490226
rect 435430 490170 435498 490226
rect 435554 490170 435622 490226
rect 435678 490170 435774 490226
rect 435154 490102 435774 490170
rect 435154 490046 435250 490102
rect 435306 490046 435374 490102
rect 435430 490046 435498 490102
rect 435554 490046 435622 490102
rect 435678 490046 435774 490102
rect 435154 489978 435774 490046
rect 435154 489922 435250 489978
rect 435306 489922 435374 489978
rect 435430 489922 435498 489978
rect 435554 489922 435622 489978
rect 435678 489922 435774 489978
rect 435154 472350 435774 489922
rect 435154 472294 435250 472350
rect 435306 472294 435374 472350
rect 435430 472294 435498 472350
rect 435554 472294 435622 472350
rect 435678 472294 435774 472350
rect 435154 472226 435774 472294
rect 435154 472170 435250 472226
rect 435306 472170 435374 472226
rect 435430 472170 435498 472226
rect 435554 472170 435622 472226
rect 435678 472170 435774 472226
rect 435154 472102 435774 472170
rect 435154 472046 435250 472102
rect 435306 472046 435374 472102
rect 435430 472046 435498 472102
rect 435554 472046 435622 472102
rect 435678 472046 435774 472102
rect 435154 471978 435774 472046
rect 435154 471922 435250 471978
rect 435306 471922 435374 471978
rect 435430 471922 435498 471978
rect 435554 471922 435622 471978
rect 435678 471922 435774 471978
rect 435154 458342 435774 471922
rect 438874 598172 439494 598268
rect 438874 598116 438970 598172
rect 439026 598116 439094 598172
rect 439150 598116 439218 598172
rect 439274 598116 439342 598172
rect 439398 598116 439494 598172
rect 438874 598048 439494 598116
rect 438874 597992 438970 598048
rect 439026 597992 439094 598048
rect 439150 597992 439218 598048
rect 439274 597992 439342 598048
rect 439398 597992 439494 598048
rect 438874 597924 439494 597992
rect 438874 597868 438970 597924
rect 439026 597868 439094 597924
rect 439150 597868 439218 597924
rect 439274 597868 439342 597924
rect 439398 597868 439494 597924
rect 438874 597800 439494 597868
rect 438874 597744 438970 597800
rect 439026 597744 439094 597800
rect 439150 597744 439218 597800
rect 439274 597744 439342 597800
rect 439398 597744 439494 597800
rect 438874 586350 439494 597744
rect 438874 586294 438970 586350
rect 439026 586294 439094 586350
rect 439150 586294 439218 586350
rect 439274 586294 439342 586350
rect 439398 586294 439494 586350
rect 438874 586226 439494 586294
rect 438874 586170 438970 586226
rect 439026 586170 439094 586226
rect 439150 586170 439218 586226
rect 439274 586170 439342 586226
rect 439398 586170 439494 586226
rect 438874 586102 439494 586170
rect 438874 586046 438970 586102
rect 439026 586046 439094 586102
rect 439150 586046 439218 586102
rect 439274 586046 439342 586102
rect 439398 586046 439494 586102
rect 438874 585978 439494 586046
rect 438874 585922 438970 585978
rect 439026 585922 439094 585978
rect 439150 585922 439218 585978
rect 439274 585922 439342 585978
rect 439398 585922 439494 585978
rect 438874 568350 439494 585922
rect 438874 568294 438970 568350
rect 439026 568294 439094 568350
rect 439150 568294 439218 568350
rect 439274 568294 439342 568350
rect 439398 568294 439494 568350
rect 438874 568226 439494 568294
rect 438874 568170 438970 568226
rect 439026 568170 439094 568226
rect 439150 568170 439218 568226
rect 439274 568170 439342 568226
rect 439398 568170 439494 568226
rect 438874 568102 439494 568170
rect 438874 568046 438970 568102
rect 439026 568046 439094 568102
rect 439150 568046 439218 568102
rect 439274 568046 439342 568102
rect 439398 568046 439494 568102
rect 438874 567978 439494 568046
rect 438874 567922 438970 567978
rect 439026 567922 439094 567978
rect 439150 567922 439218 567978
rect 439274 567922 439342 567978
rect 439398 567922 439494 567978
rect 438874 550350 439494 567922
rect 438874 550294 438970 550350
rect 439026 550294 439094 550350
rect 439150 550294 439218 550350
rect 439274 550294 439342 550350
rect 439398 550294 439494 550350
rect 438874 550226 439494 550294
rect 438874 550170 438970 550226
rect 439026 550170 439094 550226
rect 439150 550170 439218 550226
rect 439274 550170 439342 550226
rect 439398 550170 439494 550226
rect 438874 550102 439494 550170
rect 438874 550046 438970 550102
rect 439026 550046 439094 550102
rect 439150 550046 439218 550102
rect 439274 550046 439342 550102
rect 439398 550046 439494 550102
rect 438874 549978 439494 550046
rect 438874 549922 438970 549978
rect 439026 549922 439094 549978
rect 439150 549922 439218 549978
rect 439274 549922 439342 549978
rect 439398 549922 439494 549978
rect 438874 532350 439494 549922
rect 438874 532294 438970 532350
rect 439026 532294 439094 532350
rect 439150 532294 439218 532350
rect 439274 532294 439342 532350
rect 439398 532294 439494 532350
rect 438874 532226 439494 532294
rect 438874 532170 438970 532226
rect 439026 532170 439094 532226
rect 439150 532170 439218 532226
rect 439274 532170 439342 532226
rect 439398 532170 439494 532226
rect 438874 532102 439494 532170
rect 438874 532046 438970 532102
rect 439026 532046 439094 532102
rect 439150 532046 439218 532102
rect 439274 532046 439342 532102
rect 439398 532046 439494 532102
rect 438874 531978 439494 532046
rect 438874 531922 438970 531978
rect 439026 531922 439094 531978
rect 439150 531922 439218 531978
rect 439274 531922 439342 531978
rect 439398 531922 439494 531978
rect 438874 514350 439494 531922
rect 438874 514294 438970 514350
rect 439026 514294 439094 514350
rect 439150 514294 439218 514350
rect 439274 514294 439342 514350
rect 439398 514294 439494 514350
rect 438874 514226 439494 514294
rect 438874 514170 438970 514226
rect 439026 514170 439094 514226
rect 439150 514170 439218 514226
rect 439274 514170 439342 514226
rect 439398 514170 439494 514226
rect 438874 514102 439494 514170
rect 438874 514046 438970 514102
rect 439026 514046 439094 514102
rect 439150 514046 439218 514102
rect 439274 514046 439342 514102
rect 439398 514046 439494 514102
rect 438874 513978 439494 514046
rect 438874 513922 438970 513978
rect 439026 513922 439094 513978
rect 439150 513922 439218 513978
rect 439274 513922 439342 513978
rect 439398 513922 439494 513978
rect 438874 496350 439494 513922
rect 438874 496294 438970 496350
rect 439026 496294 439094 496350
rect 439150 496294 439218 496350
rect 439274 496294 439342 496350
rect 439398 496294 439494 496350
rect 438874 496226 439494 496294
rect 438874 496170 438970 496226
rect 439026 496170 439094 496226
rect 439150 496170 439218 496226
rect 439274 496170 439342 496226
rect 439398 496170 439494 496226
rect 438874 496102 439494 496170
rect 438874 496046 438970 496102
rect 439026 496046 439094 496102
rect 439150 496046 439218 496102
rect 439274 496046 439342 496102
rect 439398 496046 439494 496102
rect 438874 495978 439494 496046
rect 438874 495922 438970 495978
rect 439026 495922 439094 495978
rect 439150 495922 439218 495978
rect 439274 495922 439342 495978
rect 439398 495922 439494 495978
rect 438874 478350 439494 495922
rect 438874 478294 438970 478350
rect 439026 478294 439094 478350
rect 439150 478294 439218 478350
rect 439274 478294 439342 478350
rect 439398 478294 439494 478350
rect 438874 478226 439494 478294
rect 438874 478170 438970 478226
rect 439026 478170 439094 478226
rect 439150 478170 439218 478226
rect 439274 478170 439342 478226
rect 439398 478170 439494 478226
rect 438874 478102 439494 478170
rect 438874 478046 438970 478102
rect 439026 478046 439094 478102
rect 439150 478046 439218 478102
rect 439274 478046 439342 478102
rect 439398 478046 439494 478102
rect 438874 477978 439494 478046
rect 438874 477922 438970 477978
rect 439026 477922 439094 477978
rect 439150 477922 439218 477978
rect 439274 477922 439342 477978
rect 439398 477922 439494 477978
rect 438874 460350 439494 477922
rect 438874 460294 438970 460350
rect 439026 460294 439094 460350
rect 439150 460294 439218 460350
rect 439274 460294 439342 460350
rect 439398 460294 439494 460350
rect 438874 460226 439494 460294
rect 438874 460170 438970 460226
rect 439026 460170 439094 460226
rect 439150 460170 439218 460226
rect 439274 460170 439342 460226
rect 439398 460170 439494 460226
rect 438874 460102 439494 460170
rect 438874 460046 438970 460102
rect 439026 460046 439094 460102
rect 439150 460046 439218 460102
rect 439274 460046 439342 460102
rect 439398 460046 439494 460102
rect 438874 459978 439494 460046
rect 438874 459922 438970 459978
rect 439026 459922 439094 459978
rect 439150 459922 439218 459978
rect 439274 459922 439342 459978
rect 439398 459922 439494 459978
rect 438874 458342 439494 459922
rect 453154 597212 453774 598268
rect 453154 597156 453250 597212
rect 453306 597156 453374 597212
rect 453430 597156 453498 597212
rect 453554 597156 453622 597212
rect 453678 597156 453774 597212
rect 453154 597088 453774 597156
rect 453154 597032 453250 597088
rect 453306 597032 453374 597088
rect 453430 597032 453498 597088
rect 453554 597032 453622 597088
rect 453678 597032 453774 597088
rect 453154 596964 453774 597032
rect 453154 596908 453250 596964
rect 453306 596908 453374 596964
rect 453430 596908 453498 596964
rect 453554 596908 453622 596964
rect 453678 596908 453774 596964
rect 453154 596840 453774 596908
rect 453154 596784 453250 596840
rect 453306 596784 453374 596840
rect 453430 596784 453498 596840
rect 453554 596784 453622 596840
rect 453678 596784 453774 596840
rect 453154 580350 453774 596784
rect 453154 580294 453250 580350
rect 453306 580294 453374 580350
rect 453430 580294 453498 580350
rect 453554 580294 453622 580350
rect 453678 580294 453774 580350
rect 453154 580226 453774 580294
rect 453154 580170 453250 580226
rect 453306 580170 453374 580226
rect 453430 580170 453498 580226
rect 453554 580170 453622 580226
rect 453678 580170 453774 580226
rect 453154 580102 453774 580170
rect 453154 580046 453250 580102
rect 453306 580046 453374 580102
rect 453430 580046 453498 580102
rect 453554 580046 453622 580102
rect 453678 580046 453774 580102
rect 453154 579978 453774 580046
rect 453154 579922 453250 579978
rect 453306 579922 453374 579978
rect 453430 579922 453498 579978
rect 453554 579922 453622 579978
rect 453678 579922 453774 579978
rect 453154 562350 453774 579922
rect 453154 562294 453250 562350
rect 453306 562294 453374 562350
rect 453430 562294 453498 562350
rect 453554 562294 453622 562350
rect 453678 562294 453774 562350
rect 453154 562226 453774 562294
rect 453154 562170 453250 562226
rect 453306 562170 453374 562226
rect 453430 562170 453498 562226
rect 453554 562170 453622 562226
rect 453678 562170 453774 562226
rect 453154 562102 453774 562170
rect 453154 562046 453250 562102
rect 453306 562046 453374 562102
rect 453430 562046 453498 562102
rect 453554 562046 453622 562102
rect 453678 562046 453774 562102
rect 453154 561978 453774 562046
rect 453154 561922 453250 561978
rect 453306 561922 453374 561978
rect 453430 561922 453498 561978
rect 453554 561922 453622 561978
rect 453678 561922 453774 561978
rect 453154 544350 453774 561922
rect 453154 544294 453250 544350
rect 453306 544294 453374 544350
rect 453430 544294 453498 544350
rect 453554 544294 453622 544350
rect 453678 544294 453774 544350
rect 453154 544226 453774 544294
rect 453154 544170 453250 544226
rect 453306 544170 453374 544226
rect 453430 544170 453498 544226
rect 453554 544170 453622 544226
rect 453678 544170 453774 544226
rect 453154 544102 453774 544170
rect 453154 544046 453250 544102
rect 453306 544046 453374 544102
rect 453430 544046 453498 544102
rect 453554 544046 453622 544102
rect 453678 544046 453774 544102
rect 453154 543978 453774 544046
rect 453154 543922 453250 543978
rect 453306 543922 453374 543978
rect 453430 543922 453498 543978
rect 453554 543922 453622 543978
rect 453678 543922 453774 543978
rect 453154 526350 453774 543922
rect 453154 526294 453250 526350
rect 453306 526294 453374 526350
rect 453430 526294 453498 526350
rect 453554 526294 453622 526350
rect 453678 526294 453774 526350
rect 453154 526226 453774 526294
rect 453154 526170 453250 526226
rect 453306 526170 453374 526226
rect 453430 526170 453498 526226
rect 453554 526170 453622 526226
rect 453678 526170 453774 526226
rect 453154 526102 453774 526170
rect 453154 526046 453250 526102
rect 453306 526046 453374 526102
rect 453430 526046 453498 526102
rect 453554 526046 453622 526102
rect 453678 526046 453774 526102
rect 453154 525978 453774 526046
rect 453154 525922 453250 525978
rect 453306 525922 453374 525978
rect 453430 525922 453498 525978
rect 453554 525922 453622 525978
rect 453678 525922 453774 525978
rect 453154 508350 453774 525922
rect 453154 508294 453250 508350
rect 453306 508294 453374 508350
rect 453430 508294 453498 508350
rect 453554 508294 453622 508350
rect 453678 508294 453774 508350
rect 453154 508226 453774 508294
rect 453154 508170 453250 508226
rect 453306 508170 453374 508226
rect 453430 508170 453498 508226
rect 453554 508170 453622 508226
rect 453678 508170 453774 508226
rect 453154 508102 453774 508170
rect 453154 508046 453250 508102
rect 453306 508046 453374 508102
rect 453430 508046 453498 508102
rect 453554 508046 453622 508102
rect 453678 508046 453774 508102
rect 453154 507978 453774 508046
rect 453154 507922 453250 507978
rect 453306 507922 453374 507978
rect 453430 507922 453498 507978
rect 453554 507922 453622 507978
rect 453678 507922 453774 507978
rect 453154 490350 453774 507922
rect 453154 490294 453250 490350
rect 453306 490294 453374 490350
rect 453430 490294 453498 490350
rect 453554 490294 453622 490350
rect 453678 490294 453774 490350
rect 453154 490226 453774 490294
rect 453154 490170 453250 490226
rect 453306 490170 453374 490226
rect 453430 490170 453498 490226
rect 453554 490170 453622 490226
rect 453678 490170 453774 490226
rect 453154 490102 453774 490170
rect 453154 490046 453250 490102
rect 453306 490046 453374 490102
rect 453430 490046 453498 490102
rect 453554 490046 453622 490102
rect 453678 490046 453774 490102
rect 453154 489978 453774 490046
rect 453154 489922 453250 489978
rect 453306 489922 453374 489978
rect 453430 489922 453498 489978
rect 453554 489922 453622 489978
rect 453678 489922 453774 489978
rect 453154 472350 453774 489922
rect 453154 472294 453250 472350
rect 453306 472294 453374 472350
rect 453430 472294 453498 472350
rect 453554 472294 453622 472350
rect 453678 472294 453774 472350
rect 453154 472226 453774 472294
rect 453154 472170 453250 472226
rect 453306 472170 453374 472226
rect 453430 472170 453498 472226
rect 453554 472170 453622 472226
rect 453678 472170 453774 472226
rect 453154 472102 453774 472170
rect 453154 472046 453250 472102
rect 453306 472046 453374 472102
rect 453430 472046 453498 472102
rect 453554 472046 453622 472102
rect 453678 472046 453774 472102
rect 453154 471978 453774 472046
rect 453154 471922 453250 471978
rect 453306 471922 453374 471978
rect 453430 471922 453498 471978
rect 453554 471922 453622 471978
rect 453678 471922 453774 471978
rect 453154 458342 453774 471922
rect 456874 598172 457494 598268
rect 456874 598116 456970 598172
rect 457026 598116 457094 598172
rect 457150 598116 457218 598172
rect 457274 598116 457342 598172
rect 457398 598116 457494 598172
rect 456874 598048 457494 598116
rect 456874 597992 456970 598048
rect 457026 597992 457094 598048
rect 457150 597992 457218 598048
rect 457274 597992 457342 598048
rect 457398 597992 457494 598048
rect 456874 597924 457494 597992
rect 456874 597868 456970 597924
rect 457026 597868 457094 597924
rect 457150 597868 457218 597924
rect 457274 597868 457342 597924
rect 457398 597868 457494 597924
rect 456874 597800 457494 597868
rect 456874 597744 456970 597800
rect 457026 597744 457094 597800
rect 457150 597744 457218 597800
rect 457274 597744 457342 597800
rect 457398 597744 457494 597800
rect 456874 586350 457494 597744
rect 456874 586294 456970 586350
rect 457026 586294 457094 586350
rect 457150 586294 457218 586350
rect 457274 586294 457342 586350
rect 457398 586294 457494 586350
rect 456874 586226 457494 586294
rect 456874 586170 456970 586226
rect 457026 586170 457094 586226
rect 457150 586170 457218 586226
rect 457274 586170 457342 586226
rect 457398 586170 457494 586226
rect 456874 586102 457494 586170
rect 456874 586046 456970 586102
rect 457026 586046 457094 586102
rect 457150 586046 457218 586102
rect 457274 586046 457342 586102
rect 457398 586046 457494 586102
rect 456874 585978 457494 586046
rect 456874 585922 456970 585978
rect 457026 585922 457094 585978
rect 457150 585922 457218 585978
rect 457274 585922 457342 585978
rect 457398 585922 457494 585978
rect 456874 568350 457494 585922
rect 456874 568294 456970 568350
rect 457026 568294 457094 568350
rect 457150 568294 457218 568350
rect 457274 568294 457342 568350
rect 457398 568294 457494 568350
rect 456874 568226 457494 568294
rect 456874 568170 456970 568226
rect 457026 568170 457094 568226
rect 457150 568170 457218 568226
rect 457274 568170 457342 568226
rect 457398 568170 457494 568226
rect 456874 568102 457494 568170
rect 456874 568046 456970 568102
rect 457026 568046 457094 568102
rect 457150 568046 457218 568102
rect 457274 568046 457342 568102
rect 457398 568046 457494 568102
rect 456874 567978 457494 568046
rect 456874 567922 456970 567978
rect 457026 567922 457094 567978
rect 457150 567922 457218 567978
rect 457274 567922 457342 567978
rect 457398 567922 457494 567978
rect 456874 550350 457494 567922
rect 456874 550294 456970 550350
rect 457026 550294 457094 550350
rect 457150 550294 457218 550350
rect 457274 550294 457342 550350
rect 457398 550294 457494 550350
rect 456874 550226 457494 550294
rect 456874 550170 456970 550226
rect 457026 550170 457094 550226
rect 457150 550170 457218 550226
rect 457274 550170 457342 550226
rect 457398 550170 457494 550226
rect 456874 550102 457494 550170
rect 456874 550046 456970 550102
rect 457026 550046 457094 550102
rect 457150 550046 457218 550102
rect 457274 550046 457342 550102
rect 457398 550046 457494 550102
rect 456874 549978 457494 550046
rect 456874 549922 456970 549978
rect 457026 549922 457094 549978
rect 457150 549922 457218 549978
rect 457274 549922 457342 549978
rect 457398 549922 457494 549978
rect 456874 532350 457494 549922
rect 456874 532294 456970 532350
rect 457026 532294 457094 532350
rect 457150 532294 457218 532350
rect 457274 532294 457342 532350
rect 457398 532294 457494 532350
rect 456874 532226 457494 532294
rect 456874 532170 456970 532226
rect 457026 532170 457094 532226
rect 457150 532170 457218 532226
rect 457274 532170 457342 532226
rect 457398 532170 457494 532226
rect 456874 532102 457494 532170
rect 456874 532046 456970 532102
rect 457026 532046 457094 532102
rect 457150 532046 457218 532102
rect 457274 532046 457342 532102
rect 457398 532046 457494 532102
rect 456874 531978 457494 532046
rect 456874 531922 456970 531978
rect 457026 531922 457094 531978
rect 457150 531922 457218 531978
rect 457274 531922 457342 531978
rect 457398 531922 457494 531978
rect 456874 514350 457494 531922
rect 456874 514294 456970 514350
rect 457026 514294 457094 514350
rect 457150 514294 457218 514350
rect 457274 514294 457342 514350
rect 457398 514294 457494 514350
rect 456874 514226 457494 514294
rect 456874 514170 456970 514226
rect 457026 514170 457094 514226
rect 457150 514170 457218 514226
rect 457274 514170 457342 514226
rect 457398 514170 457494 514226
rect 456874 514102 457494 514170
rect 456874 514046 456970 514102
rect 457026 514046 457094 514102
rect 457150 514046 457218 514102
rect 457274 514046 457342 514102
rect 457398 514046 457494 514102
rect 456874 513978 457494 514046
rect 456874 513922 456970 513978
rect 457026 513922 457094 513978
rect 457150 513922 457218 513978
rect 457274 513922 457342 513978
rect 457398 513922 457494 513978
rect 456874 496350 457494 513922
rect 456874 496294 456970 496350
rect 457026 496294 457094 496350
rect 457150 496294 457218 496350
rect 457274 496294 457342 496350
rect 457398 496294 457494 496350
rect 456874 496226 457494 496294
rect 456874 496170 456970 496226
rect 457026 496170 457094 496226
rect 457150 496170 457218 496226
rect 457274 496170 457342 496226
rect 457398 496170 457494 496226
rect 456874 496102 457494 496170
rect 456874 496046 456970 496102
rect 457026 496046 457094 496102
rect 457150 496046 457218 496102
rect 457274 496046 457342 496102
rect 457398 496046 457494 496102
rect 456874 495978 457494 496046
rect 456874 495922 456970 495978
rect 457026 495922 457094 495978
rect 457150 495922 457218 495978
rect 457274 495922 457342 495978
rect 457398 495922 457494 495978
rect 456874 478350 457494 495922
rect 456874 478294 456970 478350
rect 457026 478294 457094 478350
rect 457150 478294 457218 478350
rect 457274 478294 457342 478350
rect 457398 478294 457494 478350
rect 456874 478226 457494 478294
rect 456874 478170 456970 478226
rect 457026 478170 457094 478226
rect 457150 478170 457218 478226
rect 457274 478170 457342 478226
rect 457398 478170 457494 478226
rect 456874 478102 457494 478170
rect 456874 478046 456970 478102
rect 457026 478046 457094 478102
rect 457150 478046 457218 478102
rect 457274 478046 457342 478102
rect 457398 478046 457494 478102
rect 456874 477978 457494 478046
rect 456874 477922 456970 477978
rect 457026 477922 457094 477978
rect 457150 477922 457218 477978
rect 457274 477922 457342 477978
rect 457398 477922 457494 477978
rect 456874 460350 457494 477922
rect 456874 460294 456970 460350
rect 457026 460294 457094 460350
rect 457150 460294 457218 460350
rect 457274 460294 457342 460350
rect 457398 460294 457494 460350
rect 456874 460226 457494 460294
rect 456874 460170 456970 460226
rect 457026 460170 457094 460226
rect 457150 460170 457218 460226
rect 457274 460170 457342 460226
rect 457398 460170 457494 460226
rect 456874 460102 457494 460170
rect 456874 460046 456970 460102
rect 457026 460046 457094 460102
rect 457150 460046 457218 460102
rect 457274 460046 457342 460102
rect 457398 460046 457494 460102
rect 456874 459978 457494 460046
rect 456874 459922 456970 459978
rect 457026 459922 457094 459978
rect 457150 459922 457218 459978
rect 457274 459922 457342 459978
rect 457398 459922 457494 459978
rect 456874 458342 457494 459922
rect 471154 597212 471774 598268
rect 471154 597156 471250 597212
rect 471306 597156 471374 597212
rect 471430 597156 471498 597212
rect 471554 597156 471622 597212
rect 471678 597156 471774 597212
rect 471154 597088 471774 597156
rect 471154 597032 471250 597088
rect 471306 597032 471374 597088
rect 471430 597032 471498 597088
rect 471554 597032 471622 597088
rect 471678 597032 471774 597088
rect 471154 596964 471774 597032
rect 471154 596908 471250 596964
rect 471306 596908 471374 596964
rect 471430 596908 471498 596964
rect 471554 596908 471622 596964
rect 471678 596908 471774 596964
rect 471154 596840 471774 596908
rect 471154 596784 471250 596840
rect 471306 596784 471374 596840
rect 471430 596784 471498 596840
rect 471554 596784 471622 596840
rect 471678 596784 471774 596840
rect 471154 580350 471774 596784
rect 471154 580294 471250 580350
rect 471306 580294 471374 580350
rect 471430 580294 471498 580350
rect 471554 580294 471622 580350
rect 471678 580294 471774 580350
rect 471154 580226 471774 580294
rect 471154 580170 471250 580226
rect 471306 580170 471374 580226
rect 471430 580170 471498 580226
rect 471554 580170 471622 580226
rect 471678 580170 471774 580226
rect 471154 580102 471774 580170
rect 471154 580046 471250 580102
rect 471306 580046 471374 580102
rect 471430 580046 471498 580102
rect 471554 580046 471622 580102
rect 471678 580046 471774 580102
rect 471154 579978 471774 580046
rect 471154 579922 471250 579978
rect 471306 579922 471374 579978
rect 471430 579922 471498 579978
rect 471554 579922 471622 579978
rect 471678 579922 471774 579978
rect 471154 562350 471774 579922
rect 471154 562294 471250 562350
rect 471306 562294 471374 562350
rect 471430 562294 471498 562350
rect 471554 562294 471622 562350
rect 471678 562294 471774 562350
rect 471154 562226 471774 562294
rect 471154 562170 471250 562226
rect 471306 562170 471374 562226
rect 471430 562170 471498 562226
rect 471554 562170 471622 562226
rect 471678 562170 471774 562226
rect 471154 562102 471774 562170
rect 471154 562046 471250 562102
rect 471306 562046 471374 562102
rect 471430 562046 471498 562102
rect 471554 562046 471622 562102
rect 471678 562046 471774 562102
rect 471154 561978 471774 562046
rect 471154 561922 471250 561978
rect 471306 561922 471374 561978
rect 471430 561922 471498 561978
rect 471554 561922 471622 561978
rect 471678 561922 471774 561978
rect 471154 544350 471774 561922
rect 471154 544294 471250 544350
rect 471306 544294 471374 544350
rect 471430 544294 471498 544350
rect 471554 544294 471622 544350
rect 471678 544294 471774 544350
rect 471154 544226 471774 544294
rect 471154 544170 471250 544226
rect 471306 544170 471374 544226
rect 471430 544170 471498 544226
rect 471554 544170 471622 544226
rect 471678 544170 471774 544226
rect 471154 544102 471774 544170
rect 471154 544046 471250 544102
rect 471306 544046 471374 544102
rect 471430 544046 471498 544102
rect 471554 544046 471622 544102
rect 471678 544046 471774 544102
rect 471154 543978 471774 544046
rect 471154 543922 471250 543978
rect 471306 543922 471374 543978
rect 471430 543922 471498 543978
rect 471554 543922 471622 543978
rect 471678 543922 471774 543978
rect 471154 526350 471774 543922
rect 471154 526294 471250 526350
rect 471306 526294 471374 526350
rect 471430 526294 471498 526350
rect 471554 526294 471622 526350
rect 471678 526294 471774 526350
rect 471154 526226 471774 526294
rect 471154 526170 471250 526226
rect 471306 526170 471374 526226
rect 471430 526170 471498 526226
rect 471554 526170 471622 526226
rect 471678 526170 471774 526226
rect 471154 526102 471774 526170
rect 471154 526046 471250 526102
rect 471306 526046 471374 526102
rect 471430 526046 471498 526102
rect 471554 526046 471622 526102
rect 471678 526046 471774 526102
rect 471154 525978 471774 526046
rect 471154 525922 471250 525978
rect 471306 525922 471374 525978
rect 471430 525922 471498 525978
rect 471554 525922 471622 525978
rect 471678 525922 471774 525978
rect 471154 508350 471774 525922
rect 471154 508294 471250 508350
rect 471306 508294 471374 508350
rect 471430 508294 471498 508350
rect 471554 508294 471622 508350
rect 471678 508294 471774 508350
rect 471154 508226 471774 508294
rect 471154 508170 471250 508226
rect 471306 508170 471374 508226
rect 471430 508170 471498 508226
rect 471554 508170 471622 508226
rect 471678 508170 471774 508226
rect 471154 508102 471774 508170
rect 471154 508046 471250 508102
rect 471306 508046 471374 508102
rect 471430 508046 471498 508102
rect 471554 508046 471622 508102
rect 471678 508046 471774 508102
rect 471154 507978 471774 508046
rect 471154 507922 471250 507978
rect 471306 507922 471374 507978
rect 471430 507922 471498 507978
rect 471554 507922 471622 507978
rect 471678 507922 471774 507978
rect 471154 490350 471774 507922
rect 471154 490294 471250 490350
rect 471306 490294 471374 490350
rect 471430 490294 471498 490350
rect 471554 490294 471622 490350
rect 471678 490294 471774 490350
rect 471154 490226 471774 490294
rect 471154 490170 471250 490226
rect 471306 490170 471374 490226
rect 471430 490170 471498 490226
rect 471554 490170 471622 490226
rect 471678 490170 471774 490226
rect 471154 490102 471774 490170
rect 471154 490046 471250 490102
rect 471306 490046 471374 490102
rect 471430 490046 471498 490102
rect 471554 490046 471622 490102
rect 471678 490046 471774 490102
rect 471154 489978 471774 490046
rect 471154 489922 471250 489978
rect 471306 489922 471374 489978
rect 471430 489922 471498 489978
rect 471554 489922 471622 489978
rect 471678 489922 471774 489978
rect 471154 472350 471774 489922
rect 471154 472294 471250 472350
rect 471306 472294 471374 472350
rect 471430 472294 471498 472350
rect 471554 472294 471622 472350
rect 471678 472294 471774 472350
rect 471154 472226 471774 472294
rect 471154 472170 471250 472226
rect 471306 472170 471374 472226
rect 471430 472170 471498 472226
rect 471554 472170 471622 472226
rect 471678 472170 471774 472226
rect 471154 472102 471774 472170
rect 471154 472046 471250 472102
rect 471306 472046 471374 472102
rect 471430 472046 471498 472102
rect 471554 472046 471622 472102
rect 471678 472046 471774 472102
rect 471154 471978 471774 472046
rect 471154 471922 471250 471978
rect 471306 471922 471374 471978
rect 471430 471922 471498 471978
rect 471554 471922 471622 471978
rect 471678 471922 471774 471978
rect 471154 458342 471774 471922
rect 474874 598172 475494 598268
rect 474874 598116 474970 598172
rect 475026 598116 475094 598172
rect 475150 598116 475218 598172
rect 475274 598116 475342 598172
rect 475398 598116 475494 598172
rect 474874 598048 475494 598116
rect 474874 597992 474970 598048
rect 475026 597992 475094 598048
rect 475150 597992 475218 598048
rect 475274 597992 475342 598048
rect 475398 597992 475494 598048
rect 474874 597924 475494 597992
rect 474874 597868 474970 597924
rect 475026 597868 475094 597924
rect 475150 597868 475218 597924
rect 475274 597868 475342 597924
rect 475398 597868 475494 597924
rect 474874 597800 475494 597868
rect 474874 597744 474970 597800
rect 475026 597744 475094 597800
rect 475150 597744 475218 597800
rect 475274 597744 475342 597800
rect 475398 597744 475494 597800
rect 474874 586350 475494 597744
rect 474874 586294 474970 586350
rect 475026 586294 475094 586350
rect 475150 586294 475218 586350
rect 475274 586294 475342 586350
rect 475398 586294 475494 586350
rect 474874 586226 475494 586294
rect 474874 586170 474970 586226
rect 475026 586170 475094 586226
rect 475150 586170 475218 586226
rect 475274 586170 475342 586226
rect 475398 586170 475494 586226
rect 474874 586102 475494 586170
rect 474874 586046 474970 586102
rect 475026 586046 475094 586102
rect 475150 586046 475218 586102
rect 475274 586046 475342 586102
rect 475398 586046 475494 586102
rect 474874 585978 475494 586046
rect 474874 585922 474970 585978
rect 475026 585922 475094 585978
rect 475150 585922 475218 585978
rect 475274 585922 475342 585978
rect 475398 585922 475494 585978
rect 474874 568350 475494 585922
rect 474874 568294 474970 568350
rect 475026 568294 475094 568350
rect 475150 568294 475218 568350
rect 475274 568294 475342 568350
rect 475398 568294 475494 568350
rect 474874 568226 475494 568294
rect 474874 568170 474970 568226
rect 475026 568170 475094 568226
rect 475150 568170 475218 568226
rect 475274 568170 475342 568226
rect 475398 568170 475494 568226
rect 474874 568102 475494 568170
rect 474874 568046 474970 568102
rect 475026 568046 475094 568102
rect 475150 568046 475218 568102
rect 475274 568046 475342 568102
rect 475398 568046 475494 568102
rect 474874 567978 475494 568046
rect 474874 567922 474970 567978
rect 475026 567922 475094 567978
rect 475150 567922 475218 567978
rect 475274 567922 475342 567978
rect 475398 567922 475494 567978
rect 474874 550350 475494 567922
rect 474874 550294 474970 550350
rect 475026 550294 475094 550350
rect 475150 550294 475218 550350
rect 475274 550294 475342 550350
rect 475398 550294 475494 550350
rect 474874 550226 475494 550294
rect 474874 550170 474970 550226
rect 475026 550170 475094 550226
rect 475150 550170 475218 550226
rect 475274 550170 475342 550226
rect 475398 550170 475494 550226
rect 474874 550102 475494 550170
rect 474874 550046 474970 550102
rect 475026 550046 475094 550102
rect 475150 550046 475218 550102
rect 475274 550046 475342 550102
rect 475398 550046 475494 550102
rect 474874 549978 475494 550046
rect 474874 549922 474970 549978
rect 475026 549922 475094 549978
rect 475150 549922 475218 549978
rect 475274 549922 475342 549978
rect 475398 549922 475494 549978
rect 474874 532350 475494 549922
rect 474874 532294 474970 532350
rect 475026 532294 475094 532350
rect 475150 532294 475218 532350
rect 475274 532294 475342 532350
rect 475398 532294 475494 532350
rect 474874 532226 475494 532294
rect 474874 532170 474970 532226
rect 475026 532170 475094 532226
rect 475150 532170 475218 532226
rect 475274 532170 475342 532226
rect 475398 532170 475494 532226
rect 474874 532102 475494 532170
rect 474874 532046 474970 532102
rect 475026 532046 475094 532102
rect 475150 532046 475218 532102
rect 475274 532046 475342 532102
rect 475398 532046 475494 532102
rect 474874 531978 475494 532046
rect 474874 531922 474970 531978
rect 475026 531922 475094 531978
rect 475150 531922 475218 531978
rect 475274 531922 475342 531978
rect 475398 531922 475494 531978
rect 474874 514350 475494 531922
rect 474874 514294 474970 514350
rect 475026 514294 475094 514350
rect 475150 514294 475218 514350
rect 475274 514294 475342 514350
rect 475398 514294 475494 514350
rect 474874 514226 475494 514294
rect 474874 514170 474970 514226
rect 475026 514170 475094 514226
rect 475150 514170 475218 514226
rect 475274 514170 475342 514226
rect 475398 514170 475494 514226
rect 474874 514102 475494 514170
rect 474874 514046 474970 514102
rect 475026 514046 475094 514102
rect 475150 514046 475218 514102
rect 475274 514046 475342 514102
rect 475398 514046 475494 514102
rect 474874 513978 475494 514046
rect 474874 513922 474970 513978
rect 475026 513922 475094 513978
rect 475150 513922 475218 513978
rect 475274 513922 475342 513978
rect 475398 513922 475494 513978
rect 474874 496350 475494 513922
rect 474874 496294 474970 496350
rect 475026 496294 475094 496350
rect 475150 496294 475218 496350
rect 475274 496294 475342 496350
rect 475398 496294 475494 496350
rect 474874 496226 475494 496294
rect 474874 496170 474970 496226
rect 475026 496170 475094 496226
rect 475150 496170 475218 496226
rect 475274 496170 475342 496226
rect 475398 496170 475494 496226
rect 474874 496102 475494 496170
rect 474874 496046 474970 496102
rect 475026 496046 475094 496102
rect 475150 496046 475218 496102
rect 475274 496046 475342 496102
rect 475398 496046 475494 496102
rect 474874 495978 475494 496046
rect 474874 495922 474970 495978
rect 475026 495922 475094 495978
rect 475150 495922 475218 495978
rect 475274 495922 475342 495978
rect 475398 495922 475494 495978
rect 474874 478350 475494 495922
rect 474874 478294 474970 478350
rect 475026 478294 475094 478350
rect 475150 478294 475218 478350
rect 475274 478294 475342 478350
rect 475398 478294 475494 478350
rect 474874 478226 475494 478294
rect 474874 478170 474970 478226
rect 475026 478170 475094 478226
rect 475150 478170 475218 478226
rect 475274 478170 475342 478226
rect 475398 478170 475494 478226
rect 474874 478102 475494 478170
rect 474874 478046 474970 478102
rect 475026 478046 475094 478102
rect 475150 478046 475218 478102
rect 475274 478046 475342 478102
rect 475398 478046 475494 478102
rect 474874 477978 475494 478046
rect 474874 477922 474970 477978
rect 475026 477922 475094 477978
rect 475150 477922 475218 477978
rect 475274 477922 475342 477978
rect 475398 477922 475494 477978
rect 474874 460350 475494 477922
rect 474874 460294 474970 460350
rect 475026 460294 475094 460350
rect 475150 460294 475218 460350
rect 475274 460294 475342 460350
rect 475398 460294 475494 460350
rect 474874 460226 475494 460294
rect 474874 460170 474970 460226
rect 475026 460170 475094 460226
rect 475150 460170 475218 460226
rect 475274 460170 475342 460226
rect 475398 460170 475494 460226
rect 474874 460102 475494 460170
rect 474874 460046 474970 460102
rect 475026 460046 475094 460102
rect 475150 460046 475218 460102
rect 475274 460046 475342 460102
rect 475398 460046 475494 460102
rect 474874 459978 475494 460046
rect 474874 459922 474970 459978
rect 475026 459922 475094 459978
rect 475150 459922 475218 459978
rect 475274 459922 475342 459978
rect 475398 459922 475494 459978
rect 474874 458342 475494 459922
rect 489154 597212 489774 598268
rect 489154 597156 489250 597212
rect 489306 597156 489374 597212
rect 489430 597156 489498 597212
rect 489554 597156 489622 597212
rect 489678 597156 489774 597212
rect 489154 597088 489774 597156
rect 489154 597032 489250 597088
rect 489306 597032 489374 597088
rect 489430 597032 489498 597088
rect 489554 597032 489622 597088
rect 489678 597032 489774 597088
rect 489154 596964 489774 597032
rect 489154 596908 489250 596964
rect 489306 596908 489374 596964
rect 489430 596908 489498 596964
rect 489554 596908 489622 596964
rect 489678 596908 489774 596964
rect 489154 596840 489774 596908
rect 489154 596784 489250 596840
rect 489306 596784 489374 596840
rect 489430 596784 489498 596840
rect 489554 596784 489622 596840
rect 489678 596784 489774 596840
rect 489154 580350 489774 596784
rect 489154 580294 489250 580350
rect 489306 580294 489374 580350
rect 489430 580294 489498 580350
rect 489554 580294 489622 580350
rect 489678 580294 489774 580350
rect 489154 580226 489774 580294
rect 489154 580170 489250 580226
rect 489306 580170 489374 580226
rect 489430 580170 489498 580226
rect 489554 580170 489622 580226
rect 489678 580170 489774 580226
rect 489154 580102 489774 580170
rect 489154 580046 489250 580102
rect 489306 580046 489374 580102
rect 489430 580046 489498 580102
rect 489554 580046 489622 580102
rect 489678 580046 489774 580102
rect 489154 579978 489774 580046
rect 489154 579922 489250 579978
rect 489306 579922 489374 579978
rect 489430 579922 489498 579978
rect 489554 579922 489622 579978
rect 489678 579922 489774 579978
rect 489154 562350 489774 579922
rect 489154 562294 489250 562350
rect 489306 562294 489374 562350
rect 489430 562294 489498 562350
rect 489554 562294 489622 562350
rect 489678 562294 489774 562350
rect 489154 562226 489774 562294
rect 489154 562170 489250 562226
rect 489306 562170 489374 562226
rect 489430 562170 489498 562226
rect 489554 562170 489622 562226
rect 489678 562170 489774 562226
rect 489154 562102 489774 562170
rect 489154 562046 489250 562102
rect 489306 562046 489374 562102
rect 489430 562046 489498 562102
rect 489554 562046 489622 562102
rect 489678 562046 489774 562102
rect 489154 561978 489774 562046
rect 489154 561922 489250 561978
rect 489306 561922 489374 561978
rect 489430 561922 489498 561978
rect 489554 561922 489622 561978
rect 489678 561922 489774 561978
rect 489154 544350 489774 561922
rect 489154 544294 489250 544350
rect 489306 544294 489374 544350
rect 489430 544294 489498 544350
rect 489554 544294 489622 544350
rect 489678 544294 489774 544350
rect 489154 544226 489774 544294
rect 489154 544170 489250 544226
rect 489306 544170 489374 544226
rect 489430 544170 489498 544226
rect 489554 544170 489622 544226
rect 489678 544170 489774 544226
rect 489154 544102 489774 544170
rect 489154 544046 489250 544102
rect 489306 544046 489374 544102
rect 489430 544046 489498 544102
rect 489554 544046 489622 544102
rect 489678 544046 489774 544102
rect 489154 543978 489774 544046
rect 489154 543922 489250 543978
rect 489306 543922 489374 543978
rect 489430 543922 489498 543978
rect 489554 543922 489622 543978
rect 489678 543922 489774 543978
rect 489154 526350 489774 543922
rect 489154 526294 489250 526350
rect 489306 526294 489374 526350
rect 489430 526294 489498 526350
rect 489554 526294 489622 526350
rect 489678 526294 489774 526350
rect 489154 526226 489774 526294
rect 489154 526170 489250 526226
rect 489306 526170 489374 526226
rect 489430 526170 489498 526226
rect 489554 526170 489622 526226
rect 489678 526170 489774 526226
rect 489154 526102 489774 526170
rect 489154 526046 489250 526102
rect 489306 526046 489374 526102
rect 489430 526046 489498 526102
rect 489554 526046 489622 526102
rect 489678 526046 489774 526102
rect 489154 525978 489774 526046
rect 489154 525922 489250 525978
rect 489306 525922 489374 525978
rect 489430 525922 489498 525978
rect 489554 525922 489622 525978
rect 489678 525922 489774 525978
rect 489154 508350 489774 525922
rect 489154 508294 489250 508350
rect 489306 508294 489374 508350
rect 489430 508294 489498 508350
rect 489554 508294 489622 508350
rect 489678 508294 489774 508350
rect 489154 508226 489774 508294
rect 489154 508170 489250 508226
rect 489306 508170 489374 508226
rect 489430 508170 489498 508226
rect 489554 508170 489622 508226
rect 489678 508170 489774 508226
rect 489154 508102 489774 508170
rect 489154 508046 489250 508102
rect 489306 508046 489374 508102
rect 489430 508046 489498 508102
rect 489554 508046 489622 508102
rect 489678 508046 489774 508102
rect 489154 507978 489774 508046
rect 489154 507922 489250 507978
rect 489306 507922 489374 507978
rect 489430 507922 489498 507978
rect 489554 507922 489622 507978
rect 489678 507922 489774 507978
rect 489154 490350 489774 507922
rect 489154 490294 489250 490350
rect 489306 490294 489374 490350
rect 489430 490294 489498 490350
rect 489554 490294 489622 490350
rect 489678 490294 489774 490350
rect 489154 490226 489774 490294
rect 489154 490170 489250 490226
rect 489306 490170 489374 490226
rect 489430 490170 489498 490226
rect 489554 490170 489622 490226
rect 489678 490170 489774 490226
rect 489154 490102 489774 490170
rect 489154 490046 489250 490102
rect 489306 490046 489374 490102
rect 489430 490046 489498 490102
rect 489554 490046 489622 490102
rect 489678 490046 489774 490102
rect 489154 489978 489774 490046
rect 489154 489922 489250 489978
rect 489306 489922 489374 489978
rect 489430 489922 489498 489978
rect 489554 489922 489622 489978
rect 489678 489922 489774 489978
rect 489154 472350 489774 489922
rect 489154 472294 489250 472350
rect 489306 472294 489374 472350
rect 489430 472294 489498 472350
rect 489554 472294 489622 472350
rect 489678 472294 489774 472350
rect 489154 472226 489774 472294
rect 489154 472170 489250 472226
rect 489306 472170 489374 472226
rect 489430 472170 489498 472226
rect 489554 472170 489622 472226
rect 489678 472170 489774 472226
rect 489154 472102 489774 472170
rect 489154 472046 489250 472102
rect 489306 472046 489374 472102
rect 489430 472046 489498 472102
rect 489554 472046 489622 472102
rect 489678 472046 489774 472102
rect 489154 471978 489774 472046
rect 489154 471922 489250 471978
rect 489306 471922 489374 471978
rect 489430 471922 489498 471978
rect 489554 471922 489622 471978
rect 489678 471922 489774 471978
rect 489154 458342 489774 471922
rect 492874 598172 493494 598268
rect 492874 598116 492970 598172
rect 493026 598116 493094 598172
rect 493150 598116 493218 598172
rect 493274 598116 493342 598172
rect 493398 598116 493494 598172
rect 492874 598048 493494 598116
rect 492874 597992 492970 598048
rect 493026 597992 493094 598048
rect 493150 597992 493218 598048
rect 493274 597992 493342 598048
rect 493398 597992 493494 598048
rect 492874 597924 493494 597992
rect 492874 597868 492970 597924
rect 493026 597868 493094 597924
rect 493150 597868 493218 597924
rect 493274 597868 493342 597924
rect 493398 597868 493494 597924
rect 492874 597800 493494 597868
rect 492874 597744 492970 597800
rect 493026 597744 493094 597800
rect 493150 597744 493218 597800
rect 493274 597744 493342 597800
rect 493398 597744 493494 597800
rect 492874 586350 493494 597744
rect 492874 586294 492970 586350
rect 493026 586294 493094 586350
rect 493150 586294 493218 586350
rect 493274 586294 493342 586350
rect 493398 586294 493494 586350
rect 492874 586226 493494 586294
rect 492874 586170 492970 586226
rect 493026 586170 493094 586226
rect 493150 586170 493218 586226
rect 493274 586170 493342 586226
rect 493398 586170 493494 586226
rect 492874 586102 493494 586170
rect 492874 586046 492970 586102
rect 493026 586046 493094 586102
rect 493150 586046 493218 586102
rect 493274 586046 493342 586102
rect 493398 586046 493494 586102
rect 492874 585978 493494 586046
rect 492874 585922 492970 585978
rect 493026 585922 493094 585978
rect 493150 585922 493218 585978
rect 493274 585922 493342 585978
rect 493398 585922 493494 585978
rect 492874 568350 493494 585922
rect 492874 568294 492970 568350
rect 493026 568294 493094 568350
rect 493150 568294 493218 568350
rect 493274 568294 493342 568350
rect 493398 568294 493494 568350
rect 492874 568226 493494 568294
rect 492874 568170 492970 568226
rect 493026 568170 493094 568226
rect 493150 568170 493218 568226
rect 493274 568170 493342 568226
rect 493398 568170 493494 568226
rect 492874 568102 493494 568170
rect 492874 568046 492970 568102
rect 493026 568046 493094 568102
rect 493150 568046 493218 568102
rect 493274 568046 493342 568102
rect 493398 568046 493494 568102
rect 492874 567978 493494 568046
rect 492874 567922 492970 567978
rect 493026 567922 493094 567978
rect 493150 567922 493218 567978
rect 493274 567922 493342 567978
rect 493398 567922 493494 567978
rect 492874 550350 493494 567922
rect 492874 550294 492970 550350
rect 493026 550294 493094 550350
rect 493150 550294 493218 550350
rect 493274 550294 493342 550350
rect 493398 550294 493494 550350
rect 492874 550226 493494 550294
rect 492874 550170 492970 550226
rect 493026 550170 493094 550226
rect 493150 550170 493218 550226
rect 493274 550170 493342 550226
rect 493398 550170 493494 550226
rect 492874 550102 493494 550170
rect 492874 550046 492970 550102
rect 493026 550046 493094 550102
rect 493150 550046 493218 550102
rect 493274 550046 493342 550102
rect 493398 550046 493494 550102
rect 492874 549978 493494 550046
rect 492874 549922 492970 549978
rect 493026 549922 493094 549978
rect 493150 549922 493218 549978
rect 493274 549922 493342 549978
rect 493398 549922 493494 549978
rect 492874 532350 493494 549922
rect 492874 532294 492970 532350
rect 493026 532294 493094 532350
rect 493150 532294 493218 532350
rect 493274 532294 493342 532350
rect 493398 532294 493494 532350
rect 492874 532226 493494 532294
rect 492874 532170 492970 532226
rect 493026 532170 493094 532226
rect 493150 532170 493218 532226
rect 493274 532170 493342 532226
rect 493398 532170 493494 532226
rect 492874 532102 493494 532170
rect 492874 532046 492970 532102
rect 493026 532046 493094 532102
rect 493150 532046 493218 532102
rect 493274 532046 493342 532102
rect 493398 532046 493494 532102
rect 492874 531978 493494 532046
rect 492874 531922 492970 531978
rect 493026 531922 493094 531978
rect 493150 531922 493218 531978
rect 493274 531922 493342 531978
rect 493398 531922 493494 531978
rect 492874 514350 493494 531922
rect 492874 514294 492970 514350
rect 493026 514294 493094 514350
rect 493150 514294 493218 514350
rect 493274 514294 493342 514350
rect 493398 514294 493494 514350
rect 492874 514226 493494 514294
rect 492874 514170 492970 514226
rect 493026 514170 493094 514226
rect 493150 514170 493218 514226
rect 493274 514170 493342 514226
rect 493398 514170 493494 514226
rect 492874 514102 493494 514170
rect 492874 514046 492970 514102
rect 493026 514046 493094 514102
rect 493150 514046 493218 514102
rect 493274 514046 493342 514102
rect 493398 514046 493494 514102
rect 492874 513978 493494 514046
rect 492874 513922 492970 513978
rect 493026 513922 493094 513978
rect 493150 513922 493218 513978
rect 493274 513922 493342 513978
rect 493398 513922 493494 513978
rect 492874 496350 493494 513922
rect 492874 496294 492970 496350
rect 493026 496294 493094 496350
rect 493150 496294 493218 496350
rect 493274 496294 493342 496350
rect 493398 496294 493494 496350
rect 492874 496226 493494 496294
rect 492874 496170 492970 496226
rect 493026 496170 493094 496226
rect 493150 496170 493218 496226
rect 493274 496170 493342 496226
rect 493398 496170 493494 496226
rect 492874 496102 493494 496170
rect 492874 496046 492970 496102
rect 493026 496046 493094 496102
rect 493150 496046 493218 496102
rect 493274 496046 493342 496102
rect 493398 496046 493494 496102
rect 492874 495978 493494 496046
rect 492874 495922 492970 495978
rect 493026 495922 493094 495978
rect 493150 495922 493218 495978
rect 493274 495922 493342 495978
rect 493398 495922 493494 495978
rect 492874 478350 493494 495922
rect 492874 478294 492970 478350
rect 493026 478294 493094 478350
rect 493150 478294 493218 478350
rect 493274 478294 493342 478350
rect 493398 478294 493494 478350
rect 492874 478226 493494 478294
rect 492874 478170 492970 478226
rect 493026 478170 493094 478226
rect 493150 478170 493218 478226
rect 493274 478170 493342 478226
rect 493398 478170 493494 478226
rect 492874 478102 493494 478170
rect 492874 478046 492970 478102
rect 493026 478046 493094 478102
rect 493150 478046 493218 478102
rect 493274 478046 493342 478102
rect 493398 478046 493494 478102
rect 492874 477978 493494 478046
rect 492874 477922 492970 477978
rect 493026 477922 493094 477978
rect 493150 477922 493218 477978
rect 493274 477922 493342 477978
rect 493398 477922 493494 477978
rect 492874 460350 493494 477922
rect 492874 460294 492970 460350
rect 493026 460294 493094 460350
rect 493150 460294 493218 460350
rect 493274 460294 493342 460350
rect 493398 460294 493494 460350
rect 492874 460226 493494 460294
rect 492874 460170 492970 460226
rect 493026 460170 493094 460226
rect 493150 460170 493218 460226
rect 493274 460170 493342 460226
rect 493398 460170 493494 460226
rect 492874 460102 493494 460170
rect 492874 460046 492970 460102
rect 493026 460046 493094 460102
rect 493150 460046 493218 460102
rect 493274 460046 493342 460102
rect 493398 460046 493494 460102
rect 492874 459978 493494 460046
rect 492874 459922 492970 459978
rect 493026 459922 493094 459978
rect 493150 459922 493218 459978
rect 493274 459922 493342 459978
rect 493398 459922 493494 459978
rect 492874 458342 493494 459922
rect 507154 597212 507774 598268
rect 507154 597156 507250 597212
rect 507306 597156 507374 597212
rect 507430 597156 507498 597212
rect 507554 597156 507622 597212
rect 507678 597156 507774 597212
rect 507154 597088 507774 597156
rect 507154 597032 507250 597088
rect 507306 597032 507374 597088
rect 507430 597032 507498 597088
rect 507554 597032 507622 597088
rect 507678 597032 507774 597088
rect 507154 596964 507774 597032
rect 507154 596908 507250 596964
rect 507306 596908 507374 596964
rect 507430 596908 507498 596964
rect 507554 596908 507622 596964
rect 507678 596908 507774 596964
rect 507154 596840 507774 596908
rect 507154 596784 507250 596840
rect 507306 596784 507374 596840
rect 507430 596784 507498 596840
rect 507554 596784 507622 596840
rect 507678 596784 507774 596840
rect 507154 580350 507774 596784
rect 507154 580294 507250 580350
rect 507306 580294 507374 580350
rect 507430 580294 507498 580350
rect 507554 580294 507622 580350
rect 507678 580294 507774 580350
rect 507154 580226 507774 580294
rect 507154 580170 507250 580226
rect 507306 580170 507374 580226
rect 507430 580170 507498 580226
rect 507554 580170 507622 580226
rect 507678 580170 507774 580226
rect 507154 580102 507774 580170
rect 507154 580046 507250 580102
rect 507306 580046 507374 580102
rect 507430 580046 507498 580102
rect 507554 580046 507622 580102
rect 507678 580046 507774 580102
rect 507154 579978 507774 580046
rect 507154 579922 507250 579978
rect 507306 579922 507374 579978
rect 507430 579922 507498 579978
rect 507554 579922 507622 579978
rect 507678 579922 507774 579978
rect 507154 562350 507774 579922
rect 507154 562294 507250 562350
rect 507306 562294 507374 562350
rect 507430 562294 507498 562350
rect 507554 562294 507622 562350
rect 507678 562294 507774 562350
rect 507154 562226 507774 562294
rect 507154 562170 507250 562226
rect 507306 562170 507374 562226
rect 507430 562170 507498 562226
rect 507554 562170 507622 562226
rect 507678 562170 507774 562226
rect 507154 562102 507774 562170
rect 507154 562046 507250 562102
rect 507306 562046 507374 562102
rect 507430 562046 507498 562102
rect 507554 562046 507622 562102
rect 507678 562046 507774 562102
rect 507154 561978 507774 562046
rect 507154 561922 507250 561978
rect 507306 561922 507374 561978
rect 507430 561922 507498 561978
rect 507554 561922 507622 561978
rect 507678 561922 507774 561978
rect 507154 544350 507774 561922
rect 507154 544294 507250 544350
rect 507306 544294 507374 544350
rect 507430 544294 507498 544350
rect 507554 544294 507622 544350
rect 507678 544294 507774 544350
rect 507154 544226 507774 544294
rect 507154 544170 507250 544226
rect 507306 544170 507374 544226
rect 507430 544170 507498 544226
rect 507554 544170 507622 544226
rect 507678 544170 507774 544226
rect 507154 544102 507774 544170
rect 507154 544046 507250 544102
rect 507306 544046 507374 544102
rect 507430 544046 507498 544102
rect 507554 544046 507622 544102
rect 507678 544046 507774 544102
rect 507154 543978 507774 544046
rect 507154 543922 507250 543978
rect 507306 543922 507374 543978
rect 507430 543922 507498 543978
rect 507554 543922 507622 543978
rect 507678 543922 507774 543978
rect 507154 526350 507774 543922
rect 507154 526294 507250 526350
rect 507306 526294 507374 526350
rect 507430 526294 507498 526350
rect 507554 526294 507622 526350
rect 507678 526294 507774 526350
rect 507154 526226 507774 526294
rect 507154 526170 507250 526226
rect 507306 526170 507374 526226
rect 507430 526170 507498 526226
rect 507554 526170 507622 526226
rect 507678 526170 507774 526226
rect 507154 526102 507774 526170
rect 507154 526046 507250 526102
rect 507306 526046 507374 526102
rect 507430 526046 507498 526102
rect 507554 526046 507622 526102
rect 507678 526046 507774 526102
rect 507154 525978 507774 526046
rect 507154 525922 507250 525978
rect 507306 525922 507374 525978
rect 507430 525922 507498 525978
rect 507554 525922 507622 525978
rect 507678 525922 507774 525978
rect 507154 508350 507774 525922
rect 507154 508294 507250 508350
rect 507306 508294 507374 508350
rect 507430 508294 507498 508350
rect 507554 508294 507622 508350
rect 507678 508294 507774 508350
rect 507154 508226 507774 508294
rect 507154 508170 507250 508226
rect 507306 508170 507374 508226
rect 507430 508170 507498 508226
rect 507554 508170 507622 508226
rect 507678 508170 507774 508226
rect 507154 508102 507774 508170
rect 507154 508046 507250 508102
rect 507306 508046 507374 508102
rect 507430 508046 507498 508102
rect 507554 508046 507622 508102
rect 507678 508046 507774 508102
rect 507154 507978 507774 508046
rect 507154 507922 507250 507978
rect 507306 507922 507374 507978
rect 507430 507922 507498 507978
rect 507554 507922 507622 507978
rect 507678 507922 507774 507978
rect 507154 490350 507774 507922
rect 507154 490294 507250 490350
rect 507306 490294 507374 490350
rect 507430 490294 507498 490350
rect 507554 490294 507622 490350
rect 507678 490294 507774 490350
rect 507154 490226 507774 490294
rect 507154 490170 507250 490226
rect 507306 490170 507374 490226
rect 507430 490170 507498 490226
rect 507554 490170 507622 490226
rect 507678 490170 507774 490226
rect 507154 490102 507774 490170
rect 507154 490046 507250 490102
rect 507306 490046 507374 490102
rect 507430 490046 507498 490102
rect 507554 490046 507622 490102
rect 507678 490046 507774 490102
rect 507154 489978 507774 490046
rect 507154 489922 507250 489978
rect 507306 489922 507374 489978
rect 507430 489922 507498 489978
rect 507554 489922 507622 489978
rect 507678 489922 507774 489978
rect 507154 472350 507774 489922
rect 507154 472294 507250 472350
rect 507306 472294 507374 472350
rect 507430 472294 507498 472350
rect 507554 472294 507622 472350
rect 507678 472294 507774 472350
rect 507154 472226 507774 472294
rect 507154 472170 507250 472226
rect 507306 472170 507374 472226
rect 507430 472170 507498 472226
rect 507554 472170 507622 472226
rect 507678 472170 507774 472226
rect 507154 472102 507774 472170
rect 507154 472046 507250 472102
rect 507306 472046 507374 472102
rect 507430 472046 507498 472102
rect 507554 472046 507622 472102
rect 507678 472046 507774 472102
rect 507154 471978 507774 472046
rect 507154 471922 507250 471978
rect 507306 471922 507374 471978
rect 507430 471922 507498 471978
rect 507554 471922 507622 471978
rect 507678 471922 507774 471978
rect 507154 458342 507774 471922
rect 510874 598172 511494 598268
rect 510874 598116 510970 598172
rect 511026 598116 511094 598172
rect 511150 598116 511218 598172
rect 511274 598116 511342 598172
rect 511398 598116 511494 598172
rect 510874 598048 511494 598116
rect 510874 597992 510970 598048
rect 511026 597992 511094 598048
rect 511150 597992 511218 598048
rect 511274 597992 511342 598048
rect 511398 597992 511494 598048
rect 510874 597924 511494 597992
rect 510874 597868 510970 597924
rect 511026 597868 511094 597924
rect 511150 597868 511218 597924
rect 511274 597868 511342 597924
rect 511398 597868 511494 597924
rect 510874 597800 511494 597868
rect 510874 597744 510970 597800
rect 511026 597744 511094 597800
rect 511150 597744 511218 597800
rect 511274 597744 511342 597800
rect 511398 597744 511494 597800
rect 510874 586350 511494 597744
rect 510874 586294 510970 586350
rect 511026 586294 511094 586350
rect 511150 586294 511218 586350
rect 511274 586294 511342 586350
rect 511398 586294 511494 586350
rect 510874 586226 511494 586294
rect 510874 586170 510970 586226
rect 511026 586170 511094 586226
rect 511150 586170 511218 586226
rect 511274 586170 511342 586226
rect 511398 586170 511494 586226
rect 510874 586102 511494 586170
rect 510874 586046 510970 586102
rect 511026 586046 511094 586102
rect 511150 586046 511218 586102
rect 511274 586046 511342 586102
rect 511398 586046 511494 586102
rect 510874 585978 511494 586046
rect 510874 585922 510970 585978
rect 511026 585922 511094 585978
rect 511150 585922 511218 585978
rect 511274 585922 511342 585978
rect 511398 585922 511494 585978
rect 510874 568350 511494 585922
rect 510874 568294 510970 568350
rect 511026 568294 511094 568350
rect 511150 568294 511218 568350
rect 511274 568294 511342 568350
rect 511398 568294 511494 568350
rect 510874 568226 511494 568294
rect 510874 568170 510970 568226
rect 511026 568170 511094 568226
rect 511150 568170 511218 568226
rect 511274 568170 511342 568226
rect 511398 568170 511494 568226
rect 510874 568102 511494 568170
rect 510874 568046 510970 568102
rect 511026 568046 511094 568102
rect 511150 568046 511218 568102
rect 511274 568046 511342 568102
rect 511398 568046 511494 568102
rect 510874 567978 511494 568046
rect 510874 567922 510970 567978
rect 511026 567922 511094 567978
rect 511150 567922 511218 567978
rect 511274 567922 511342 567978
rect 511398 567922 511494 567978
rect 510874 550350 511494 567922
rect 510874 550294 510970 550350
rect 511026 550294 511094 550350
rect 511150 550294 511218 550350
rect 511274 550294 511342 550350
rect 511398 550294 511494 550350
rect 510874 550226 511494 550294
rect 510874 550170 510970 550226
rect 511026 550170 511094 550226
rect 511150 550170 511218 550226
rect 511274 550170 511342 550226
rect 511398 550170 511494 550226
rect 510874 550102 511494 550170
rect 510874 550046 510970 550102
rect 511026 550046 511094 550102
rect 511150 550046 511218 550102
rect 511274 550046 511342 550102
rect 511398 550046 511494 550102
rect 510874 549978 511494 550046
rect 510874 549922 510970 549978
rect 511026 549922 511094 549978
rect 511150 549922 511218 549978
rect 511274 549922 511342 549978
rect 511398 549922 511494 549978
rect 510874 532350 511494 549922
rect 510874 532294 510970 532350
rect 511026 532294 511094 532350
rect 511150 532294 511218 532350
rect 511274 532294 511342 532350
rect 511398 532294 511494 532350
rect 510874 532226 511494 532294
rect 510874 532170 510970 532226
rect 511026 532170 511094 532226
rect 511150 532170 511218 532226
rect 511274 532170 511342 532226
rect 511398 532170 511494 532226
rect 510874 532102 511494 532170
rect 510874 532046 510970 532102
rect 511026 532046 511094 532102
rect 511150 532046 511218 532102
rect 511274 532046 511342 532102
rect 511398 532046 511494 532102
rect 510874 531978 511494 532046
rect 510874 531922 510970 531978
rect 511026 531922 511094 531978
rect 511150 531922 511218 531978
rect 511274 531922 511342 531978
rect 511398 531922 511494 531978
rect 510874 514350 511494 531922
rect 510874 514294 510970 514350
rect 511026 514294 511094 514350
rect 511150 514294 511218 514350
rect 511274 514294 511342 514350
rect 511398 514294 511494 514350
rect 510874 514226 511494 514294
rect 510874 514170 510970 514226
rect 511026 514170 511094 514226
rect 511150 514170 511218 514226
rect 511274 514170 511342 514226
rect 511398 514170 511494 514226
rect 510874 514102 511494 514170
rect 510874 514046 510970 514102
rect 511026 514046 511094 514102
rect 511150 514046 511218 514102
rect 511274 514046 511342 514102
rect 511398 514046 511494 514102
rect 510874 513978 511494 514046
rect 510874 513922 510970 513978
rect 511026 513922 511094 513978
rect 511150 513922 511218 513978
rect 511274 513922 511342 513978
rect 511398 513922 511494 513978
rect 510874 496350 511494 513922
rect 510874 496294 510970 496350
rect 511026 496294 511094 496350
rect 511150 496294 511218 496350
rect 511274 496294 511342 496350
rect 511398 496294 511494 496350
rect 510874 496226 511494 496294
rect 510874 496170 510970 496226
rect 511026 496170 511094 496226
rect 511150 496170 511218 496226
rect 511274 496170 511342 496226
rect 511398 496170 511494 496226
rect 510874 496102 511494 496170
rect 510874 496046 510970 496102
rect 511026 496046 511094 496102
rect 511150 496046 511218 496102
rect 511274 496046 511342 496102
rect 511398 496046 511494 496102
rect 510874 495978 511494 496046
rect 510874 495922 510970 495978
rect 511026 495922 511094 495978
rect 511150 495922 511218 495978
rect 511274 495922 511342 495978
rect 511398 495922 511494 495978
rect 510874 478350 511494 495922
rect 510874 478294 510970 478350
rect 511026 478294 511094 478350
rect 511150 478294 511218 478350
rect 511274 478294 511342 478350
rect 511398 478294 511494 478350
rect 510874 478226 511494 478294
rect 510874 478170 510970 478226
rect 511026 478170 511094 478226
rect 511150 478170 511218 478226
rect 511274 478170 511342 478226
rect 511398 478170 511494 478226
rect 510874 478102 511494 478170
rect 510874 478046 510970 478102
rect 511026 478046 511094 478102
rect 511150 478046 511218 478102
rect 511274 478046 511342 478102
rect 511398 478046 511494 478102
rect 510874 477978 511494 478046
rect 510874 477922 510970 477978
rect 511026 477922 511094 477978
rect 511150 477922 511218 477978
rect 511274 477922 511342 477978
rect 511398 477922 511494 477978
rect 510874 460350 511494 477922
rect 510874 460294 510970 460350
rect 511026 460294 511094 460350
rect 511150 460294 511218 460350
rect 511274 460294 511342 460350
rect 511398 460294 511494 460350
rect 510874 460226 511494 460294
rect 510874 460170 510970 460226
rect 511026 460170 511094 460226
rect 511150 460170 511218 460226
rect 511274 460170 511342 460226
rect 511398 460170 511494 460226
rect 510874 460102 511494 460170
rect 510874 460046 510970 460102
rect 511026 460046 511094 460102
rect 511150 460046 511218 460102
rect 511274 460046 511342 460102
rect 511398 460046 511494 460102
rect 510874 459978 511494 460046
rect 510874 459922 510970 459978
rect 511026 459922 511094 459978
rect 511150 459922 511218 459978
rect 511274 459922 511342 459978
rect 511398 459922 511494 459978
rect 510874 458342 511494 459922
rect 525154 597212 525774 598268
rect 525154 597156 525250 597212
rect 525306 597156 525374 597212
rect 525430 597156 525498 597212
rect 525554 597156 525622 597212
rect 525678 597156 525774 597212
rect 525154 597088 525774 597156
rect 525154 597032 525250 597088
rect 525306 597032 525374 597088
rect 525430 597032 525498 597088
rect 525554 597032 525622 597088
rect 525678 597032 525774 597088
rect 525154 596964 525774 597032
rect 525154 596908 525250 596964
rect 525306 596908 525374 596964
rect 525430 596908 525498 596964
rect 525554 596908 525622 596964
rect 525678 596908 525774 596964
rect 525154 596840 525774 596908
rect 525154 596784 525250 596840
rect 525306 596784 525374 596840
rect 525430 596784 525498 596840
rect 525554 596784 525622 596840
rect 525678 596784 525774 596840
rect 525154 580350 525774 596784
rect 525154 580294 525250 580350
rect 525306 580294 525374 580350
rect 525430 580294 525498 580350
rect 525554 580294 525622 580350
rect 525678 580294 525774 580350
rect 525154 580226 525774 580294
rect 525154 580170 525250 580226
rect 525306 580170 525374 580226
rect 525430 580170 525498 580226
rect 525554 580170 525622 580226
rect 525678 580170 525774 580226
rect 525154 580102 525774 580170
rect 525154 580046 525250 580102
rect 525306 580046 525374 580102
rect 525430 580046 525498 580102
rect 525554 580046 525622 580102
rect 525678 580046 525774 580102
rect 525154 579978 525774 580046
rect 525154 579922 525250 579978
rect 525306 579922 525374 579978
rect 525430 579922 525498 579978
rect 525554 579922 525622 579978
rect 525678 579922 525774 579978
rect 525154 562350 525774 579922
rect 525154 562294 525250 562350
rect 525306 562294 525374 562350
rect 525430 562294 525498 562350
rect 525554 562294 525622 562350
rect 525678 562294 525774 562350
rect 525154 562226 525774 562294
rect 525154 562170 525250 562226
rect 525306 562170 525374 562226
rect 525430 562170 525498 562226
rect 525554 562170 525622 562226
rect 525678 562170 525774 562226
rect 525154 562102 525774 562170
rect 525154 562046 525250 562102
rect 525306 562046 525374 562102
rect 525430 562046 525498 562102
rect 525554 562046 525622 562102
rect 525678 562046 525774 562102
rect 525154 561978 525774 562046
rect 525154 561922 525250 561978
rect 525306 561922 525374 561978
rect 525430 561922 525498 561978
rect 525554 561922 525622 561978
rect 525678 561922 525774 561978
rect 525154 544350 525774 561922
rect 525154 544294 525250 544350
rect 525306 544294 525374 544350
rect 525430 544294 525498 544350
rect 525554 544294 525622 544350
rect 525678 544294 525774 544350
rect 525154 544226 525774 544294
rect 525154 544170 525250 544226
rect 525306 544170 525374 544226
rect 525430 544170 525498 544226
rect 525554 544170 525622 544226
rect 525678 544170 525774 544226
rect 525154 544102 525774 544170
rect 525154 544046 525250 544102
rect 525306 544046 525374 544102
rect 525430 544046 525498 544102
rect 525554 544046 525622 544102
rect 525678 544046 525774 544102
rect 525154 543978 525774 544046
rect 525154 543922 525250 543978
rect 525306 543922 525374 543978
rect 525430 543922 525498 543978
rect 525554 543922 525622 543978
rect 525678 543922 525774 543978
rect 525154 526350 525774 543922
rect 525154 526294 525250 526350
rect 525306 526294 525374 526350
rect 525430 526294 525498 526350
rect 525554 526294 525622 526350
rect 525678 526294 525774 526350
rect 525154 526226 525774 526294
rect 525154 526170 525250 526226
rect 525306 526170 525374 526226
rect 525430 526170 525498 526226
rect 525554 526170 525622 526226
rect 525678 526170 525774 526226
rect 525154 526102 525774 526170
rect 525154 526046 525250 526102
rect 525306 526046 525374 526102
rect 525430 526046 525498 526102
rect 525554 526046 525622 526102
rect 525678 526046 525774 526102
rect 525154 525978 525774 526046
rect 525154 525922 525250 525978
rect 525306 525922 525374 525978
rect 525430 525922 525498 525978
rect 525554 525922 525622 525978
rect 525678 525922 525774 525978
rect 525154 508350 525774 525922
rect 525154 508294 525250 508350
rect 525306 508294 525374 508350
rect 525430 508294 525498 508350
rect 525554 508294 525622 508350
rect 525678 508294 525774 508350
rect 525154 508226 525774 508294
rect 525154 508170 525250 508226
rect 525306 508170 525374 508226
rect 525430 508170 525498 508226
rect 525554 508170 525622 508226
rect 525678 508170 525774 508226
rect 525154 508102 525774 508170
rect 525154 508046 525250 508102
rect 525306 508046 525374 508102
rect 525430 508046 525498 508102
rect 525554 508046 525622 508102
rect 525678 508046 525774 508102
rect 525154 507978 525774 508046
rect 525154 507922 525250 507978
rect 525306 507922 525374 507978
rect 525430 507922 525498 507978
rect 525554 507922 525622 507978
rect 525678 507922 525774 507978
rect 525154 490350 525774 507922
rect 525154 490294 525250 490350
rect 525306 490294 525374 490350
rect 525430 490294 525498 490350
rect 525554 490294 525622 490350
rect 525678 490294 525774 490350
rect 525154 490226 525774 490294
rect 525154 490170 525250 490226
rect 525306 490170 525374 490226
rect 525430 490170 525498 490226
rect 525554 490170 525622 490226
rect 525678 490170 525774 490226
rect 525154 490102 525774 490170
rect 525154 490046 525250 490102
rect 525306 490046 525374 490102
rect 525430 490046 525498 490102
rect 525554 490046 525622 490102
rect 525678 490046 525774 490102
rect 525154 489978 525774 490046
rect 525154 489922 525250 489978
rect 525306 489922 525374 489978
rect 525430 489922 525498 489978
rect 525554 489922 525622 489978
rect 525678 489922 525774 489978
rect 525154 472350 525774 489922
rect 525154 472294 525250 472350
rect 525306 472294 525374 472350
rect 525430 472294 525498 472350
rect 525554 472294 525622 472350
rect 525678 472294 525774 472350
rect 525154 472226 525774 472294
rect 525154 472170 525250 472226
rect 525306 472170 525374 472226
rect 525430 472170 525498 472226
rect 525554 472170 525622 472226
rect 525678 472170 525774 472226
rect 525154 472102 525774 472170
rect 525154 472046 525250 472102
rect 525306 472046 525374 472102
rect 525430 472046 525498 472102
rect 525554 472046 525622 472102
rect 525678 472046 525774 472102
rect 525154 471978 525774 472046
rect 525154 471922 525250 471978
rect 525306 471922 525374 471978
rect 525430 471922 525498 471978
rect 525554 471922 525622 471978
rect 525678 471922 525774 471978
rect 525154 458342 525774 471922
rect 528874 598172 529494 598268
rect 528874 598116 528970 598172
rect 529026 598116 529094 598172
rect 529150 598116 529218 598172
rect 529274 598116 529342 598172
rect 529398 598116 529494 598172
rect 528874 598048 529494 598116
rect 528874 597992 528970 598048
rect 529026 597992 529094 598048
rect 529150 597992 529218 598048
rect 529274 597992 529342 598048
rect 529398 597992 529494 598048
rect 528874 597924 529494 597992
rect 528874 597868 528970 597924
rect 529026 597868 529094 597924
rect 529150 597868 529218 597924
rect 529274 597868 529342 597924
rect 529398 597868 529494 597924
rect 528874 597800 529494 597868
rect 528874 597744 528970 597800
rect 529026 597744 529094 597800
rect 529150 597744 529218 597800
rect 529274 597744 529342 597800
rect 529398 597744 529494 597800
rect 528874 586350 529494 597744
rect 528874 586294 528970 586350
rect 529026 586294 529094 586350
rect 529150 586294 529218 586350
rect 529274 586294 529342 586350
rect 529398 586294 529494 586350
rect 528874 586226 529494 586294
rect 528874 586170 528970 586226
rect 529026 586170 529094 586226
rect 529150 586170 529218 586226
rect 529274 586170 529342 586226
rect 529398 586170 529494 586226
rect 528874 586102 529494 586170
rect 528874 586046 528970 586102
rect 529026 586046 529094 586102
rect 529150 586046 529218 586102
rect 529274 586046 529342 586102
rect 529398 586046 529494 586102
rect 528874 585978 529494 586046
rect 528874 585922 528970 585978
rect 529026 585922 529094 585978
rect 529150 585922 529218 585978
rect 529274 585922 529342 585978
rect 529398 585922 529494 585978
rect 528874 568350 529494 585922
rect 528874 568294 528970 568350
rect 529026 568294 529094 568350
rect 529150 568294 529218 568350
rect 529274 568294 529342 568350
rect 529398 568294 529494 568350
rect 528874 568226 529494 568294
rect 528874 568170 528970 568226
rect 529026 568170 529094 568226
rect 529150 568170 529218 568226
rect 529274 568170 529342 568226
rect 529398 568170 529494 568226
rect 528874 568102 529494 568170
rect 528874 568046 528970 568102
rect 529026 568046 529094 568102
rect 529150 568046 529218 568102
rect 529274 568046 529342 568102
rect 529398 568046 529494 568102
rect 528874 567978 529494 568046
rect 528874 567922 528970 567978
rect 529026 567922 529094 567978
rect 529150 567922 529218 567978
rect 529274 567922 529342 567978
rect 529398 567922 529494 567978
rect 528874 550350 529494 567922
rect 528874 550294 528970 550350
rect 529026 550294 529094 550350
rect 529150 550294 529218 550350
rect 529274 550294 529342 550350
rect 529398 550294 529494 550350
rect 528874 550226 529494 550294
rect 528874 550170 528970 550226
rect 529026 550170 529094 550226
rect 529150 550170 529218 550226
rect 529274 550170 529342 550226
rect 529398 550170 529494 550226
rect 528874 550102 529494 550170
rect 528874 550046 528970 550102
rect 529026 550046 529094 550102
rect 529150 550046 529218 550102
rect 529274 550046 529342 550102
rect 529398 550046 529494 550102
rect 528874 549978 529494 550046
rect 528874 549922 528970 549978
rect 529026 549922 529094 549978
rect 529150 549922 529218 549978
rect 529274 549922 529342 549978
rect 529398 549922 529494 549978
rect 528874 532350 529494 549922
rect 528874 532294 528970 532350
rect 529026 532294 529094 532350
rect 529150 532294 529218 532350
rect 529274 532294 529342 532350
rect 529398 532294 529494 532350
rect 528874 532226 529494 532294
rect 528874 532170 528970 532226
rect 529026 532170 529094 532226
rect 529150 532170 529218 532226
rect 529274 532170 529342 532226
rect 529398 532170 529494 532226
rect 528874 532102 529494 532170
rect 528874 532046 528970 532102
rect 529026 532046 529094 532102
rect 529150 532046 529218 532102
rect 529274 532046 529342 532102
rect 529398 532046 529494 532102
rect 528874 531978 529494 532046
rect 528874 531922 528970 531978
rect 529026 531922 529094 531978
rect 529150 531922 529218 531978
rect 529274 531922 529342 531978
rect 529398 531922 529494 531978
rect 528874 514350 529494 531922
rect 528874 514294 528970 514350
rect 529026 514294 529094 514350
rect 529150 514294 529218 514350
rect 529274 514294 529342 514350
rect 529398 514294 529494 514350
rect 528874 514226 529494 514294
rect 528874 514170 528970 514226
rect 529026 514170 529094 514226
rect 529150 514170 529218 514226
rect 529274 514170 529342 514226
rect 529398 514170 529494 514226
rect 528874 514102 529494 514170
rect 528874 514046 528970 514102
rect 529026 514046 529094 514102
rect 529150 514046 529218 514102
rect 529274 514046 529342 514102
rect 529398 514046 529494 514102
rect 528874 513978 529494 514046
rect 528874 513922 528970 513978
rect 529026 513922 529094 513978
rect 529150 513922 529218 513978
rect 529274 513922 529342 513978
rect 529398 513922 529494 513978
rect 528874 496350 529494 513922
rect 528874 496294 528970 496350
rect 529026 496294 529094 496350
rect 529150 496294 529218 496350
rect 529274 496294 529342 496350
rect 529398 496294 529494 496350
rect 528874 496226 529494 496294
rect 528874 496170 528970 496226
rect 529026 496170 529094 496226
rect 529150 496170 529218 496226
rect 529274 496170 529342 496226
rect 529398 496170 529494 496226
rect 528874 496102 529494 496170
rect 528874 496046 528970 496102
rect 529026 496046 529094 496102
rect 529150 496046 529218 496102
rect 529274 496046 529342 496102
rect 529398 496046 529494 496102
rect 528874 495978 529494 496046
rect 528874 495922 528970 495978
rect 529026 495922 529094 495978
rect 529150 495922 529218 495978
rect 529274 495922 529342 495978
rect 529398 495922 529494 495978
rect 528874 478350 529494 495922
rect 528874 478294 528970 478350
rect 529026 478294 529094 478350
rect 529150 478294 529218 478350
rect 529274 478294 529342 478350
rect 529398 478294 529494 478350
rect 528874 478226 529494 478294
rect 528874 478170 528970 478226
rect 529026 478170 529094 478226
rect 529150 478170 529218 478226
rect 529274 478170 529342 478226
rect 529398 478170 529494 478226
rect 528874 478102 529494 478170
rect 528874 478046 528970 478102
rect 529026 478046 529094 478102
rect 529150 478046 529218 478102
rect 529274 478046 529342 478102
rect 529398 478046 529494 478102
rect 528874 477978 529494 478046
rect 528874 477922 528970 477978
rect 529026 477922 529094 477978
rect 529150 477922 529218 477978
rect 529274 477922 529342 477978
rect 529398 477922 529494 477978
rect 528874 460350 529494 477922
rect 528874 460294 528970 460350
rect 529026 460294 529094 460350
rect 529150 460294 529218 460350
rect 529274 460294 529342 460350
rect 529398 460294 529494 460350
rect 528874 460226 529494 460294
rect 528874 460170 528970 460226
rect 529026 460170 529094 460226
rect 529150 460170 529218 460226
rect 529274 460170 529342 460226
rect 529398 460170 529494 460226
rect 528874 460102 529494 460170
rect 528874 460046 528970 460102
rect 529026 460046 529094 460102
rect 529150 460046 529218 460102
rect 529274 460046 529342 460102
rect 529398 460046 529494 460102
rect 528874 459978 529494 460046
rect 528874 459922 528970 459978
rect 529026 459922 529094 459978
rect 529150 459922 529218 459978
rect 529274 459922 529342 459978
rect 529398 459922 529494 459978
rect 528874 458342 529494 459922
rect 543154 597212 543774 598268
rect 543154 597156 543250 597212
rect 543306 597156 543374 597212
rect 543430 597156 543498 597212
rect 543554 597156 543622 597212
rect 543678 597156 543774 597212
rect 543154 597088 543774 597156
rect 543154 597032 543250 597088
rect 543306 597032 543374 597088
rect 543430 597032 543498 597088
rect 543554 597032 543622 597088
rect 543678 597032 543774 597088
rect 543154 596964 543774 597032
rect 543154 596908 543250 596964
rect 543306 596908 543374 596964
rect 543430 596908 543498 596964
rect 543554 596908 543622 596964
rect 543678 596908 543774 596964
rect 543154 596840 543774 596908
rect 543154 596784 543250 596840
rect 543306 596784 543374 596840
rect 543430 596784 543498 596840
rect 543554 596784 543622 596840
rect 543678 596784 543774 596840
rect 543154 580350 543774 596784
rect 543154 580294 543250 580350
rect 543306 580294 543374 580350
rect 543430 580294 543498 580350
rect 543554 580294 543622 580350
rect 543678 580294 543774 580350
rect 543154 580226 543774 580294
rect 543154 580170 543250 580226
rect 543306 580170 543374 580226
rect 543430 580170 543498 580226
rect 543554 580170 543622 580226
rect 543678 580170 543774 580226
rect 543154 580102 543774 580170
rect 543154 580046 543250 580102
rect 543306 580046 543374 580102
rect 543430 580046 543498 580102
rect 543554 580046 543622 580102
rect 543678 580046 543774 580102
rect 543154 579978 543774 580046
rect 543154 579922 543250 579978
rect 543306 579922 543374 579978
rect 543430 579922 543498 579978
rect 543554 579922 543622 579978
rect 543678 579922 543774 579978
rect 543154 562350 543774 579922
rect 543154 562294 543250 562350
rect 543306 562294 543374 562350
rect 543430 562294 543498 562350
rect 543554 562294 543622 562350
rect 543678 562294 543774 562350
rect 543154 562226 543774 562294
rect 543154 562170 543250 562226
rect 543306 562170 543374 562226
rect 543430 562170 543498 562226
rect 543554 562170 543622 562226
rect 543678 562170 543774 562226
rect 543154 562102 543774 562170
rect 543154 562046 543250 562102
rect 543306 562046 543374 562102
rect 543430 562046 543498 562102
rect 543554 562046 543622 562102
rect 543678 562046 543774 562102
rect 543154 561978 543774 562046
rect 543154 561922 543250 561978
rect 543306 561922 543374 561978
rect 543430 561922 543498 561978
rect 543554 561922 543622 561978
rect 543678 561922 543774 561978
rect 543154 544350 543774 561922
rect 543154 544294 543250 544350
rect 543306 544294 543374 544350
rect 543430 544294 543498 544350
rect 543554 544294 543622 544350
rect 543678 544294 543774 544350
rect 543154 544226 543774 544294
rect 543154 544170 543250 544226
rect 543306 544170 543374 544226
rect 543430 544170 543498 544226
rect 543554 544170 543622 544226
rect 543678 544170 543774 544226
rect 543154 544102 543774 544170
rect 543154 544046 543250 544102
rect 543306 544046 543374 544102
rect 543430 544046 543498 544102
rect 543554 544046 543622 544102
rect 543678 544046 543774 544102
rect 543154 543978 543774 544046
rect 543154 543922 543250 543978
rect 543306 543922 543374 543978
rect 543430 543922 543498 543978
rect 543554 543922 543622 543978
rect 543678 543922 543774 543978
rect 543154 526350 543774 543922
rect 543154 526294 543250 526350
rect 543306 526294 543374 526350
rect 543430 526294 543498 526350
rect 543554 526294 543622 526350
rect 543678 526294 543774 526350
rect 543154 526226 543774 526294
rect 543154 526170 543250 526226
rect 543306 526170 543374 526226
rect 543430 526170 543498 526226
rect 543554 526170 543622 526226
rect 543678 526170 543774 526226
rect 543154 526102 543774 526170
rect 543154 526046 543250 526102
rect 543306 526046 543374 526102
rect 543430 526046 543498 526102
rect 543554 526046 543622 526102
rect 543678 526046 543774 526102
rect 543154 525978 543774 526046
rect 543154 525922 543250 525978
rect 543306 525922 543374 525978
rect 543430 525922 543498 525978
rect 543554 525922 543622 525978
rect 543678 525922 543774 525978
rect 543154 508350 543774 525922
rect 543154 508294 543250 508350
rect 543306 508294 543374 508350
rect 543430 508294 543498 508350
rect 543554 508294 543622 508350
rect 543678 508294 543774 508350
rect 543154 508226 543774 508294
rect 543154 508170 543250 508226
rect 543306 508170 543374 508226
rect 543430 508170 543498 508226
rect 543554 508170 543622 508226
rect 543678 508170 543774 508226
rect 543154 508102 543774 508170
rect 543154 508046 543250 508102
rect 543306 508046 543374 508102
rect 543430 508046 543498 508102
rect 543554 508046 543622 508102
rect 543678 508046 543774 508102
rect 543154 507978 543774 508046
rect 543154 507922 543250 507978
rect 543306 507922 543374 507978
rect 543430 507922 543498 507978
rect 543554 507922 543622 507978
rect 543678 507922 543774 507978
rect 543154 490350 543774 507922
rect 543154 490294 543250 490350
rect 543306 490294 543374 490350
rect 543430 490294 543498 490350
rect 543554 490294 543622 490350
rect 543678 490294 543774 490350
rect 543154 490226 543774 490294
rect 543154 490170 543250 490226
rect 543306 490170 543374 490226
rect 543430 490170 543498 490226
rect 543554 490170 543622 490226
rect 543678 490170 543774 490226
rect 543154 490102 543774 490170
rect 543154 490046 543250 490102
rect 543306 490046 543374 490102
rect 543430 490046 543498 490102
rect 543554 490046 543622 490102
rect 543678 490046 543774 490102
rect 543154 489978 543774 490046
rect 543154 489922 543250 489978
rect 543306 489922 543374 489978
rect 543430 489922 543498 489978
rect 543554 489922 543622 489978
rect 543678 489922 543774 489978
rect 543154 472350 543774 489922
rect 543154 472294 543250 472350
rect 543306 472294 543374 472350
rect 543430 472294 543498 472350
rect 543554 472294 543622 472350
rect 543678 472294 543774 472350
rect 543154 472226 543774 472294
rect 543154 472170 543250 472226
rect 543306 472170 543374 472226
rect 543430 472170 543498 472226
rect 543554 472170 543622 472226
rect 543678 472170 543774 472226
rect 543154 472102 543774 472170
rect 543154 472046 543250 472102
rect 543306 472046 543374 472102
rect 543430 472046 543498 472102
rect 543554 472046 543622 472102
rect 543678 472046 543774 472102
rect 543154 471978 543774 472046
rect 543154 471922 543250 471978
rect 543306 471922 543374 471978
rect 543430 471922 543498 471978
rect 543554 471922 543622 471978
rect 543678 471922 543774 471978
rect 543154 458342 543774 471922
rect 546874 598172 547494 598268
rect 546874 598116 546970 598172
rect 547026 598116 547094 598172
rect 547150 598116 547218 598172
rect 547274 598116 547342 598172
rect 547398 598116 547494 598172
rect 546874 598048 547494 598116
rect 546874 597992 546970 598048
rect 547026 597992 547094 598048
rect 547150 597992 547218 598048
rect 547274 597992 547342 598048
rect 547398 597992 547494 598048
rect 546874 597924 547494 597992
rect 546874 597868 546970 597924
rect 547026 597868 547094 597924
rect 547150 597868 547218 597924
rect 547274 597868 547342 597924
rect 547398 597868 547494 597924
rect 546874 597800 547494 597868
rect 546874 597744 546970 597800
rect 547026 597744 547094 597800
rect 547150 597744 547218 597800
rect 547274 597744 547342 597800
rect 547398 597744 547494 597800
rect 546874 586350 547494 597744
rect 546874 586294 546970 586350
rect 547026 586294 547094 586350
rect 547150 586294 547218 586350
rect 547274 586294 547342 586350
rect 547398 586294 547494 586350
rect 546874 586226 547494 586294
rect 546874 586170 546970 586226
rect 547026 586170 547094 586226
rect 547150 586170 547218 586226
rect 547274 586170 547342 586226
rect 547398 586170 547494 586226
rect 546874 586102 547494 586170
rect 546874 586046 546970 586102
rect 547026 586046 547094 586102
rect 547150 586046 547218 586102
rect 547274 586046 547342 586102
rect 547398 586046 547494 586102
rect 546874 585978 547494 586046
rect 546874 585922 546970 585978
rect 547026 585922 547094 585978
rect 547150 585922 547218 585978
rect 547274 585922 547342 585978
rect 547398 585922 547494 585978
rect 546874 568350 547494 585922
rect 546874 568294 546970 568350
rect 547026 568294 547094 568350
rect 547150 568294 547218 568350
rect 547274 568294 547342 568350
rect 547398 568294 547494 568350
rect 546874 568226 547494 568294
rect 546874 568170 546970 568226
rect 547026 568170 547094 568226
rect 547150 568170 547218 568226
rect 547274 568170 547342 568226
rect 547398 568170 547494 568226
rect 546874 568102 547494 568170
rect 546874 568046 546970 568102
rect 547026 568046 547094 568102
rect 547150 568046 547218 568102
rect 547274 568046 547342 568102
rect 547398 568046 547494 568102
rect 546874 567978 547494 568046
rect 546874 567922 546970 567978
rect 547026 567922 547094 567978
rect 547150 567922 547218 567978
rect 547274 567922 547342 567978
rect 547398 567922 547494 567978
rect 546874 550350 547494 567922
rect 546874 550294 546970 550350
rect 547026 550294 547094 550350
rect 547150 550294 547218 550350
rect 547274 550294 547342 550350
rect 547398 550294 547494 550350
rect 546874 550226 547494 550294
rect 546874 550170 546970 550226
rect 547026 550170 547094 550226
rect 547150 550170 547218 550226
rect 547274 550170 547342 550226
rect 547398 550170 547494 550226
rect 546874 550102 547494 550170
rect 546874 550046 546970 550102
rect 547026 550046 547094 550102
rect 547150 550046 547218 550102
rect 547274 550046 547342 550102
rect 547398 550046 547494 550102
rect 546874 549978 547494 550046
rect 546874 549922 546970 549978
rect 547026 549922 547094 549978
rect 547150 549922 547218 549978
rect 547274 549922 547342 549978
rect 547398 549922 547494 549978
rect 546874 532350 547494 549922
rect 546874 532294 546970 532350
rect 547026 532294 547094 532350
rect 547150 532294 547218 532350
rect 547274 532294 547342 532350
rect 547398 532294 547494 532350
rect 546874 532226 547494 532294
rect 546874 532170 546970 532226
rect 547026 532170 547094 532226
rect 547150 532170 547218 532226
rect 547274 532170 547342 532226
rect 547398 532170 547494 532226
rect 546874 532102 547494 532170
rect 546874 532046 546970 532102
rect 547026 532046 547094 532102
rect 547150 532046 547218 532102
rect 547274 532046 547342 532102
rect 547398 532046 547494 532102
rect 546874 531978 547494 532046
rect 546874 531922 546970 531978
rect 547026 531922 547094 531978
rect 547150 531922 547218 531978
rect 547274 531922 547342 531978
rect 547398 531922 547494 531978
rect 546874 514350 547494 531922
rect 546874 514294 546970 514350
rect 547026 514294 547094 514350
rect 547150 514294 547218 514350
rect 547274 514294 547342 514350
rect 547398 514294 547494 514350
rect 546874 514226 547494 514294
rect 546874 514170 546970 514226
rect 547026 514170 547094 514226
rect 547150 514170 547218 514226
rect 547274 514170 547342 514226
rect 547398 514170 547494 514226
rect 546874 514102 547494 514170
rect 546874 514046 546970 514102
rect 547026 514046 547094 514102
rect 547150 514046 547218 514102
rect 547274 514046 547342 514102
rect 547398 514046 547494 514102
rect 546874 513978 547494 514046
rect 546874 513922 546970 513978
rect 547026 513922 547094 513978
rect 547150 513922 547218 513978
rect 547274 513922 547342 513978
rect 547398 513922 547494 513978
rect 546874 496350 547494 513922
rect 546874 496294 546970 496350
rect 547026 496294 547094 496350
rect 547150 496294 547218 496350
rect 547274 496294 547342 496350
rect 547398 496294 547494 496350
rect 546874 496226 547494 496294
rect 546874 496170 546970 496226
rect 547026 496170 547094 496226
rect 547150 496170 547218 496226
rect 547274 496170 547342 496226
rect 547398 496170 547494 496226
rect 546874 496102 547494 496170
rect 546874 496046 546970 496102
rect 547026 496046 547094 496102
rect 547150 496046 547218 496102
rect 547274 496046 547342 496102
rect 547398 496046 547494 496102
rect 546874 495978 547494 496046
rect 546874 495922 546970 495978
rect 547026 495922 547094 495978
rect 547150 495922 547218 495978
rect 547274 495922 547342 495978
rect 547398 495922 547494 495978
rect 546874 478350 547494 495922
rect 546874 478294 546970 478350
rect 547026 478294 547094 478350
rect 547150 478294 547218 478350
rect 547274 478294 547342 478350
rect 547398 478294 547494 478350
rect 546874 478226 547494 478294
rect 546874 478170 546970 478226
rect 547026 478170 547094 478226
rect 547150 478170 547218 478226
rect 547274 478170 547342 478226
rect 547398 478170 547494 478226
rect 546874 478102 547494 478170
rect 546874 478046 546970 478102
rect 547026 478046 547094 478102
rect 547150 478046 547218 478102
rect 547274 478046 547342 478102
rect 547398 478046 547494 478102
rect 546874 477978 547494 478046
rect 546874 477922 546970 477978
rect 547026 477922 547094 477978
rect 547150 477922 547218 477978
rect 547274 477922 547342 477978
rect 547398 477922 547494 477978
rect 546874 460350 547494 477922
rect 546874 460294 546970 460350
rect 547026 460294 547094 460350
rect 547150 460294 547218 460350
rect 547274 460294 547342 460350
rect 547398 460294 547494 460350
rect 546874 460226 547494 460294
rect 546874 460170 546970 460226
rect 547026 460170 547094 460226
rect 547150 460170 547218 460226
rect 547274 460170 547342 460226
rect 547398 460170 547494 460226
rect 546874 460102 547494 460170
rect 546874 460046 546970 460102
rect 547026 460046 547094 460102
rect 547150 460046 547218 460102
rect 547274 460046 547342 460102
rect 547398 460046 547494 460102
rect 546874 459978 547494 460046
rect 546874 459922 546970 459978
rect 547026 459922 547094 459978
rect 547150 459922 547218 459978
rect 547274 459922 547342 459978
rect 547398 459922 547494 459978
rect 546874 458342 547494 459922
rect 561154 597212 561774 598268
rect 561154 597156 561250 597212
rect 561306 597156 561374 597212
rect 561430 597156 561498 597212
rect 561554 597156 561622 597212
rect 561678 597156 561774 597212
rect 561154 597088 561774 597156
rect 561154 597032 561250 597088
rect 561306 597032 561374 597088
rect 561430 597032 561498 597088
rect 561554 597032 561622 597088
rect 561678 597032 561774 597088
rect 561154 596964 561774 597032
rect 561154 596908 561250 596964
rect 561306 596908 561374 596964
rect 561430 596908 561498 596964
rect 561554 596908 561622 596964
rect 561678 596908 561774 596964
rect 561154 596840 561774 596908
rect 561154 596784 561250 596840
rect 561306 596784 561374 596840
rect 561430 596784 561498 596840
rect 561554 596784 561622 596840
rect 561678 596784 561774 596840
rect 561154 580350 561774 596784
rect 561154 580294 561250 580350
rect 561306 580294 561374 580350
rect 561430 580294 561498 580350
rect 561554 580294 561622 580350
rect 561678 580294 561774 580350
rect 561154 580226 561774 580294
rect 561154 580170 561250 580226
rect 561306 580170 561374 580226
rect 561430 580170 561498 580226
rect 561554 580170 561622 580226
rect 561678 580170 561774 580226
rect 561154 580102 561774 580170
rect 561154 580046 561250 580102
rect 561306 580046 561374 580102
rect 561430 580046 561498 580102
rect 561554 580046 561622 580102
rect 561678 580046 561774 580102
rect 561154 579978 561774 580046
rect 561154 579922 561250 579978
rect 561306 579922 561374 579978
rect 561430 579922 561498 579978
rect 561554 579922 561622 579978
rect 561678 579922 561774 579978
rect 561154 562350 561774 579922
rect 561154 562294 561250 562350
rect 561306 562294 561374 562350
rect 561430 562294 561498 562350
rect 561554 562294 561622 562350
rect 561678 562294 561774 562350
rect 561154 562226 561774 562294
rect 561154 562170 561250 562226
rect 561306 562170 561374 562226
rect 561430 562170 561498 562226
rect 561554 562170 561622 562226
rect 561678 562170 561774 562226
rect 561154 562102 561774 562170
rect 561154 562046 561250 562102
rect 561306 562046 561374 562102
rect 561430 562046 561498 562102
rect 561554 562046 561622 562102
rect 561678 562046 561774 562102
rect 561154 561978 561774 562046
rect 561154 561922 561250 561978
rect 561306 561922 561374 561978
rect 561430 561922 561498 561978
rect 561554 561922 561622 561978
rect 561678 561922 561774 561978
rect 561154 544350 561774 561922
rect 561154 544294 561250 544350
rect 561306 544294 561374 544350
rect 561430 544294 561498 544350
rect 561554 544294 561622 544350
rect 561678 544294 561774 544350
rect 561154 544226 561774 544294
rect 561154 544170 561250 544226
rect 561306 544170 561374 544226
rect 561430 544170 561498 544226
rect 561554 544170 561622 544226
rect 561678 544170 561774 544226
rect 561154 544102 561774 544170
rect 561154 544046 561250 544102
rect 561306 544046 561374 544102
rect 561430 544046 561498 544102
rect 561554 544046 561622 544102
rect 561678 544046 561774 544102
rect 561154 543978 561774 544046
rect 561154 543922 561250 543978
rect 561306 543922 561374 543978
rect 561430 543922 561498 543978
rect 561554 543922 561622 543978
rect 561678 543922 561774 543978
rect 561154 526350 561774 543922
rect 561154 526294 561250 526350
rect 561306 526294 561374 526350
rect 561430 526294 561498 526350
rect 561554 526294 561622 526350
rect 561678 526294 561774 526350
rect 561154 526226 561774 526294
rect 561154 526170 561250 526226
rect 561306 526170 561374 526226
rect 561430 526170 561498 526226
rect 561554 526170 561622 526226
rect 561678 526170 561774 526226
rect 561154 526102 561774 526170
rect 561154 526046 561250 526102
rect 561306 526046 561374 526102
rect 561430 526046 561498 526102
rect 561554 526046 561622 526102
rect 561678 526046 561774 526102
rect 561154 525978 561774 526046
rect 561154 525922 561250 525978
rect 561306 525922 561374 525978
rect 561430 525922 561498 525978
rect 561554 525922 561622 525978
rect 561678 525922 561774 525978
rect 561154 508350 561774 525922
rect 561154 508294 561250 508350
rect 561306 508294 561374 508350
rect 561430 508294 561498 508350
rect 561554 508294 561622 508350
rect 561678 508294 561774 508350
rect 561154 508226 561774 508294
rect 561154 508170 561250 508226
rect 561306 508170 561374 508226
rect 561430 508170 561498 508226
rect 561554 508170 561622 508226
rect 561678 508170 561774 508226
rect 561154 508102 561774 508170
rect 561154 508046 561250 508102
rect 561306 508046 561374 508102
rect 561430 508046 561498 508102
rect 561554 508046 561622 508102
rect 561678 508046 561774 508102
rect 561154 507978 561774 508046
rect 561154 507922 561250 507978
rect 561306 507922 561374 507978
rect 561430 507922 561498 507978
rect 561554 507922 561622 507978
rect 561678 507922 561774 507978
rect 561154 490350 561774 507922
rect 561154 490294 561250 490350
rect 561306 490294 561374 490350
rect 561430 490294 561498 490350
rect 561554 490294 561622 490350
rect 561678 490294 561774 490350
rect 561154 490226 561774 490294
rect 561154 490170 561250 490226
rect 561306 490170 561374 490226
rect 561430 490170 561498 490226
rect 561554 490170 561622 490226
rect 561678 490170 561774 490226
rect 561154 490102 561774 490170
rect 561154 490046 561250 490102
rect 561306 490046 561374 490102
rect 561430 490046 561498 490102
rect 561554 490046 561622 490102
rect 561678 490046 561774 490102
rect 561154 489978 561774 490046
rect 561154 489922 561250 489978
rect 561306 489922 561374 489978
rect 561430 489922 561498 489978
rect 561554 489922 561622 489978
rect 561678 489922 561774 489978
rect 561154 472350 561774 489922
rect 561154 472294 561250 472350
rect 561306 472294 561374 472350
rect 561430 472294 561498 472350
rect 561554 472294 561622 472350
rect 561678 472294 561774 472350
rect 561154 472226 561774 472294
rect 561154 472170 561250 472226
rect 561306 472170 561374 472226
rect 561430 472170 561498 472226
rect 561554 472170 561622 472226
rect 561678 472170 561774 472226
rect 561154 472102 561774 472170
rect 561154 472046 561250 472102
rect 561306 472046 561374 472102
rect 561430 472046 561498 472102
rect 561554 472046 561622 472102
rect 561678 472046 561774 472102
rect 561154 471978 561774 472046
rect 561154 471922 561250 471978
rect 561306 471922 561374 471978
rect 561430 471922 561498 471978
rect 561554 471922 561622 471978
rect 561678 471922 561774 471978
rect 561154 458342 561774 471922
rect 564874 598172 565494 598268
rect 564874 598116 564970 598172
rect 565026 598116 565094 598172
rect 565150 598116 565218 598172
rect 565274 598116 565342 598172
rect 565398 598116 565494 598172
rect 564874 598048 565494 598116
rect 564874 597992 564970 598048
rect 565026 597992 565094 598048
rect 565150 597992 565218 598048
rect 565274 597992 565342 598048
rect 565398 597992 565494 598048
rect 564874 597924 565494 597992
rect 564874 597868 564970 597924
rect 565026 597868 565094 597924
rect 565150 597868 565218 597924
rect 565274 597868 565342 597924
rect 565398 597868 565494 597924
rect 564874 597800 565494 597868
rect 564874 597744 564970 597800
rect 565026 597744 565094 597800
rect 565150 597744 565218 597800
rect 565274 597744 565342 597800
rect 565398 597744 565494 597800
rect 564874 586350 565494 597744
rect 564874 586294 564970 586350
rect 565026 586294 565094 586350
rect 565150 586294 565218 586350
rect 565274 586294 565342 586350
rect 565398 586294 565494 586350
rect 564874 586226 565494 586294
rect 564874 586170 564970 586226
rect 565026 586170 565094 586226
rect 565150 586170 565218 586226
rect 565274 586170 565342 586226
rect 565398 586170 565494 586226
rect 564874 586102 565494 586170
rect 564874 586046 564970 586102
rect 565026 586046 565094 586102
rect 565150 586046 565218 586102
rect 565274 586046 565342 586102
rect 565398 586046 565494 586102
rect 564874 585978 565494 586046
rect 564874 585922 564970 585978
rect 565026 585922 565094 585978
rect 565150 585922 565218 585978
rect 565274 585922 565342 585978
rect 565398 585922 565494 585978
rect 564874 568350 565494 585922
rect 564874 568294 564970 568350
rect 565026 568294 565094 568350
rect 565150 568294 565218 568350
rect 565274 568294 565342 568350
rect 565398 568294 565494 568350
rect 564874 568226 565494 568294
rect 564874 568170 564970 568226
rect 565026 568170 565094 568226
rect 565150 568170 565218 568226
rect 565274 568170 565342 568226
rect 565398 568170 565494 568226
rect 564874 568102 565494 568170
rect 564874 568046 564970 568102
rect 565026 568046 565094 568102
rect 565150 568046 565218 568102
rect 565274 568046 565342 568102
rect 565398 568046 565494 568102
rect 564874 567978 565494 568046
rect 564874 567922 564970 567978
rect 565026 567922 565094 567978
rect 565150 567922 565218 567978
rect 565274 567922 565342 567978
rect 565398 567922 565494 567978
rect 564874 550350 565494 567922
rect 564874 550294 564970 550350
rect 565026 550294 565094 550350
rect 565150 550294 565218 550350
rect 565274 550294 565342 550350
rect 565398 550294 565494 550350
rect 564874 550226 565494 550294
rect 564874 550170 564970 550226
rect 565026 550170 565094 550226
rect 565150 550170 565218 550226
rect 565274 550170 565342 550226
rect 565398 550170 565494 550226
rect 564874 550102 565494 550170
rect 564874 550046 564970 550102
rect 565026 550046 565094 550102
rect 565150 550046 565218 550102
rect 565274 550046 565342 550102
rect 565398 550046 565494 550102
rect 564874 549978 565494 550046
rect 564874 549922 564970 549978
rect 565026 549922 565094 549978
rect 565150 549922 565218 549978
rect 565274 549922 565342 549978
rect 565398 549922 565494 549978
rect 564874 532350 565494 549922
rect 564874 532294 564970 532350
rect 565026 532294 565094 532350
rect 565150 532294 565218 532350
rect 565274 532294 565342 532350
rect 565398 532294 565494 532350
rect 564874 532226 565494 532294
rect 564874 532170 564970 532226
rect 565026 532170 565094 532226
rect 565150 532170 565218 532226
rect 565274 532170 565342 532226
rect 565398 532170 565494 532226
rect 564874 532102 565494 532170
rect 564874 532046 564970 532102
rect 565026 532046 565094 532102
rect 565150 532046 565218 532102
rect 565274 532046 565342 532102
rect 565398 532046 565494 532102
rect 564874 531978 565494 532046
rect 564874 531922 564970 531978
rect 565026 531922 565094 531978
rect 565150 531922 565218 531978
rect 565274 531922 565342 531978
rect 565398 531922 565494 531978
rect 564874 514350 565494 531922
rect 564874 514294 564970 514350
rect 565026 514294 565094 514350
rect 565150 514294 565218 514350
rect 565274 514294 565342 514350
rect 565398 514294 565494 514350
rect 564874 514226 565494 514294
rect 564874 514170 564970 514226
rect 565026 514170 565094 514226
rect 565150 514170 565218 514226
rect 565274 514170 565342 514226
rect 565398 514170 565494 514226
rect 564874 514102 565494 514170
rect 564874 514046 564970 514102
rect 565026 514046 565094 514102
rect 565150 514046 565218 514102
rect 565274 514046 565342 514102
rect 565398 514046 565494 514102
rect 564874 513978 565494 514046
rect 564874 513922 564970 513978
rect 565026 513922 565094 513978
rect 565150 513922 565218 513978
rect 565274 513922 565342 513978
rect 565398 513922 565494 513978
rect 564874 496350 565494 513922
rect 564874 496294 564970 496350
rect 565026 496294 565094 496350
rect 565150 496294 565218 496350
rect 565274 496294 565342 496350
rect 565398 496294 565494 496350
rect 564874 496226 565494 496294
rect 564874 496170 564970 496226
rect 565026 496170 565094 496226
rect 565150 496170 565218 496226
rect 565274 496170 565342 496226
rect 565398 496170 565494 496226
rect 564874 496102 565494 496170
rect 564874 496046 564970 496102
rect 565026 496046 565094 496102
rect 565150 496046 565218 496102
rect 565274 496046 565342 496102
rect 565398 496046 565494 496102
rect 564874 495978 565494 496046
rect 564874 495922 564970 495978
rect 565026 495922 565094 495978
rect 565150 495922 565218 495978
rect 565274 495922 565342 495978
rect 565398 495922 565494 495978
rect 564874 478350 565494 495922
rect 564874 478294 564970 478350
rect 565026 478294 565094 478350
rect 565150 478294 565218 478350
rect 565274 478294 565342 478350
rect 565398 478294 565494 478350
rect 564874 478226 565494 478294
rect 564874 478170 564970 478226
rect 565026 478170 565094 478226
rect 565150 478170 565218 478226
rect 565274 478170 565342 478226
rect 565398 478170 565494 478226
rect 564874 478102 565494 478170
rect 564874 478046 564970 478102
rect 565026 478046 565094 478102
rect 565150 478046 565218 478102
rect 565274 478046 565342 478102
rect 565398 478046 565494 478102
rect 564874 477978 565494 478046
rect 564874 477922 564970 477978
rect 565026 477922 565094 477978
rect 565150 477922 565218 477978
rect 565274 477922 565342 477978
rect 565398 477922 565494 477978
rect 564874 460350 565494 477922
rect 564874 460294 564970 460350
rect 565026 460294 565094 460350
rect 565150 460294 565218 460350
rect 565274 460294 565342 460350
rect 565398 460294 565494 460350
rect 564874 460226 565494 460294
rect 564874 460170 564970 460226
rect 565026 460170 565094 460226
rect 565150 460170 565218 460226
rect 565274 460170 565342 460226
rect 565398 460170 565494 460226
rect 564874 460102 565494 460170
rect 564874 460046 564970 460102
rect 565026 460046 565094 460102
rect 565150 460046 565218 460102
rect 565274 460046 565342 460102
rect 565398 460046 565494 460102
rect 564874 459978 565494 460046
rect 564874 459922 564970 459978
rect 565026 459922 565094 459978
rect 565150 459922 565218 459978
rect 565274 459922 565342 459978
rect 565398 459922 565494 459978
rect 564874 458342 565494 459922
rect 579154 597212 579774 598268
rect 579154 597156 579250 597212
rect 579306 597156 579374 597212
rect 579430 597156 579498 597212
rect 579554 597156 579622 597212
rect 579678 597156 579774 597212
rect 579154 597088 579774 597156
rect 579154 597032 579250 597088
rect 579306 597032 579374 597088
rect 579430 597032 579498 597088
rect 579554 597032 579622 597088
rect 579678 597032 579774 597088
rect 579154 596964 579774 597032
rect 579154 596908 579250 596964
rect 579306 596908 579374 596964
rect 579430 596908 579498 596964
rect 579554 596908 579622 596964
rect 579678 596908 579774 596964
rect 579154 596840 579774 596908
rect 579154 596784 579250 596840
rect 579306 596784 579374 596840
rect 579430 596784 579498 596840
rect 579554 596784 579622 596840
rect 579678 596784 579774 596840
rect 579154 580350 579774 596784
rect 579154 580294 579250 580350
rect 579306 580294 579374 580350
rect 579430 580294 579498 580350
rect 579554 580294 579622 580350
rect 579678 580294 579774 580350
rect 579154 580226 579774 580294
rect 579154 580170 579250 580226
rect 579306 580170 579374 580226
rect 579430 580170 579498 580226
rect 579554 580170 579622 580226
rect 579678 580170 579774 580226
rect 579154 580102 579774 580170
rect 579154 580046 579250 580102
rect 579306 580046 579374 580102
rect 579430 580046 579498 580102
rect 579554 580046 579622 580102
rect 579678 580046 579774 580102
rect 579154 579978 579774 580046
rect 579154 579922 579250 579978
rect 579306 579922 579374 579978
rect 579430 579922 579498 579978
rect 579554 579922 579622 579978
rect 579678 579922 579774 579978
rect 579154 562350 579774 579922
rect 579154 562294 579250 562350
rect 579306 562294 579374 562350
rect 579430 562294 579498 562350
rect 579554 562294 579622 562350
rect 579678 562294 579774 562350
rect 579154 562226 579774 562294
rect 579154 562170 579250 562226
rect 579306 562170 579374 562226
rect 579430 562170 579498 562226
rect 579554 562170 579622 562226
rect 579678 562170 579774 562226
rect 579154 562102 579774 562170
rect 579154 562046 579250 562102
rect 579306 562046 579374 562102
rect 579430 562046 579498 562102
rect 579554 562046 579622 562102
rect 579678 562046 579774 562102
rect 579154 561978 579774 562046
rect 579154 561922 579250 561978
rect 579306 561922 579374 561978
rect 579430 561922 579498 561978
rect 579554 561922 579622 561978
rect 579678 561922 579774 561978
rect 579154 544350 579774 561922
rect 579154 544294 579250 544350
rect 579306 544294 579374 544350
rect 579430 544294 579498 544350
rect 579554 544294 579622 544350
rect 579678 544294 579774 544350
rect 579154 544226 579774 544294
rect 579154 544170 579250 544226
rect 579306 544170 579374 544226
rect 579430 544170 579498 544226
rect 579554 544170 579622 544226
rect 579678 544170 579774 544226
rect 579154 544102 579774 544170
rect 579154 544046 579250 544102
rect 579306 544046 579374 544102
rect 579430 544046 579498 544102
rect 579554 544046 579622 544102
rect 579678 544046 579774 544102
rect 579154 543978 579774 544046
rect 579154 543922 579250 543978
rect 579306 543922 579374 543978
rect 579430 543922 579498 543978
rect 579554 543922 579622 543978
rect 579678 543922 579774 543978
rect 579154 526350 579774 543922
rect 579154 526294 579250 526350
rect 579306 526294 579374 526350
rect 579430 526294 579498 526350
rect 579554 526294 579622 526350
rect 579678 526294 579774 526350
rect 579154 526226 579774 526294
rect 579154 526170 579250 526226
rect 579306 526170 579374 526226
rect 579430 526170 579498 526226
rect 579554 526170 579622 526226
rect 579678 526170 579774 526226
rect 579154 526102 579774 526170
rect 579154 526046 579250 526102
rect 579306 526046 579374 526102
rect 579430 526046 579498 526102
rect 579554 526046 579622 526102
rect 579678 526046 579774 526102
rect 579154 525978 579774 526046
rect 579154 525922 579250 525978
rect 579306 525922 579374 525978
rect 579430 525922 579498 525978
rect 579554 525922 579622 525978
rect 579678 525922 579774 525978
rect 579154 508350 579774 525922
rect 579154 508294 579250 508350
rect 579306 508294 579374 508350
rect 579430 508294 579498 508350
rect 579554 508294 579622 508350
rect 579678 508294 579774 508350
rect 579154 508226 579774 508294
rect 579154 508170 579250 508226
rect 579306 508170 579374 508226
rect 579430 508170 579498 508226
rect 579554 508170 579622 508226
rect 579678 508170 579774 508226
rect 579154 508102 579774 508170
rect 579154 508046 579250 508102
rect 579306 508046 579374 508102
rect 579430 508046 579498 508102
rect 579554 508046 579622 508102
rect 579678 508046 579774 508102
rect 579154 507978 579774 508046
rect 579154 507922 579250 507978
rect 579306 507922 579374 507978
rect 579430 507922 579498 507978
rect 579554 507922 579622 507978
rect 579678 507922 579774 507978
rect 579154 490350 579774 507922
rect 579154 490294 579250 490350
rect 579306 490294 579374 490350
rect 579430 490294 579498 490350
rect 579554 490294 579622 490350
rect 579678 490294 579774 490350
rect 579154 490226 579774 490294
rect 579154 490170 579250 490226
rect 579306 490170 579374 490226
rect 579430 490170 579498 490226
rect 579554 490170 579622 490226
rect 579678 490170 579774 490226
rect 579154 490102 579774 490170
rect 579154 490046 579250 490102
rect 579306 490046 579374 490102
rect 579430 490046 579498 490102
rect 579554 490046 579622 490102
rect 579678 490046 579774 490102
rect 579154 489978 579774 490046
rect 579154 489922 579250 489978
rect 579306 489922 579374 489978
rect 579430 489922 579498 489978
rect 579554 489922 579622 489978
rect 579678 489922 579774 489978
rect 579154 472350 579774 489922
rect 579154 472294 579250 472350
rect 579306 472294 579374 472350
rect 579430 472294 579498 472350
rect 579554 472294 579622 472350
rect 579678 472294 579774 472350
rect 579154 472226 579774 472294
rect 579154 472170 579250 472226
rect 579306 472170 579374 472226
rect 579430 472170 579498 472226
rect 579554 472170 579622 472226
rect 579678 472170 579774 472226
rect 579154 472102 579774 472170
rect 579154 472046 579250 472102
rect 579306 472046 579374 472102
rect 579430 472046 579498 472102
rect 579554 472046 579622 472102
rect 579678 472046 579774 472102
rect 579154 471978 579774 472046
rect 579154 471922 579250 471978
rect 579306 471922 579374 471978
rect 579430 471922 579498 471978
rect 579554 471922 579622 471978
rect 579678 471922 579774 471978
rect 402874 442294 402970 442350
rect 403026 442294 403094 442350
rect 403150 442294 403218 442350
rect 403274 442294 403342 442350
rect 403398 442294 403494 442350
rect 402874 442226 403494 442294
rect 402874 442170 402970 442226
rect 403026 442170 403094 442226
rect 403150 442170 403218 442226
rect 403274 442170 403342 442226
rect 403398 442170 403494 442226
rect 402874 442102 403494 442170
rect 402874 442046 402970 442102
rect 403026 442046 403094 442102
rect 403150 442046 403218 442102
rect 403274 442046 403342 442102
rect 403398 442046 403494 442102
rect 402874 441978 403494 442046
rect 402874 441922 402970 441978
rect 403026 441922 403094 441978
rect 403150 441922 403218 441978
rect 403274 441922 403342 441978
rect 403398 441922 403494 441978
rect 402874 424350 403494 441922
rect 402874 424294 402970 424350
rect 403026 424294 403094 424350
rect 403150 424294 403218 424350
rect 403274 424294 403342 424350
rect 403398 424294 403494 424350
rect 402874 424226 403494 424294
rect 402874 424170 402970 424226
rect 403026 424170 403094 424226
rect 403150 424170 403218 424226
rect 403274 424170 403342 424226
rect 403398 424170 403494 424226
rect 402874 424102 403494 424170
rect 402874 424046 402970 424102
rect 403026 424046 403094 424102
rect 403150 424046 403218 424102
rect 403274 424046 403342 424102
rect 403398 424046 403494 424102
rect 402874 423978 403494 424046
rect 402874 423922 402970 423978
rect 403026 423922 403094 423978
rect 403150 423922 403218 423978
rect 403274 423922 403342 423978
rect 403398 423922 403494 423978
rect 402874 406350 403494 423922
rect 402874 406294 402970 406350
rect 403026 406294 403094 406350
rect 403150 406294 403218 406350
rect 403274 406294 403342 406350
rect 403398 406294 403494 406350
rect 402874 406226 403494 406294
rect 402874 406170 402970 406226
rect 403026 406170 403094 406226
rect 403150 406170 403218 406226
rect 403274 406170 403342 406226
rect 403398 406170 403494 406226
rect 402874 406102 403494 406170
rect 402874 406046 402970 406102
rect 403026 406046 403094 406102
rect 403150 406046 403218 406102
rect 403274 406046 403342 406102
rect 403398 406046 403494 406102
rect 402874 405978 403494 406046
rect 402874 405922 402970 405978
rect 403026 405922 403094 405978
rect 403150 405922 403218 405978
rect 403274 405922 403342 405978
rect 403398 405922 403494 405978
rect 402874 388350 403494 405922
rect 402874 388294 402970 388350
rect 403026 388294 403094 388350
rect 403150 388294 403218 388350
rect 403274 388294 403342 388350
rect 403398 388294 403494 388350
rect 402874 388226 403494 388294
rect 402874 388170 402970 388226
rect 403026 388170 403094 388226
rect 403150 388170 403218 388226
rect 403274 388170 403342 388226
rect 403398 388170 403494 388226
rect 402874 388102 403494 388170
rect 402874 388046 402970 388102
rect 403026 388046 403094 388102
rect 403150 388046 403218 388102
rect 403274 388046 403342 388102
rect 403398 388046 403494 388102
rect 402874 387978 403494 388046
rect 402874 387922 402970 387978
rect 403026 387922 403094 387978
rect 403150 387922 403218 387978
rect 403274 387922 403342 387978
rect 403398 387922 403494 387978
rect 402874 370350 403494 387922
rect 402874 370294 402970 370350
rect 403026 370294 403094 370350
rect 403150 370294 403218 370350
rect 403274 370294 403342 370350
rect 403398 370294 403494 370350
rect 402874 370226 403494 370294
rect 402874 370170 402970 370226
rect 403026 370170 403094 370226
rect 403150 370170 403218 370226
rect 403274 370170 403342 370226
rect 403398 370170 403494 370226
rect 402874 370102 403494 370170
rect 402874 370046 402970 370102
rect 403026 370046 403094 370102
rect 403150 370046 403218 370102
rect 403274 370046 403342 370102
rect 403398 370046 403494 370102
rect 402874 369978 403494 370046
rect 402874 369922 402970 369978
rect 403026 369922 403094 369978
rect 403150 369922 403218 369978
rect 403274 369922 403342 369978
rect 403398 369922 403494 369978
rect 402874 352350 403494 369922
rect 402874 352294 402970 352350
rect 403026 352294 403094 352350
rect 403150 352294 403218 352350
rect 403274 352294 403342 352350
rect 403398 352294 403494 352350
rect 402874 352226 403494 352294
rect 402874 352170 402970 352226
rect 403026 352170 403094 352226
rect 403150 352170 403218 352226
rect 403274 352170 403342 352226
rect 403398 352170 403494 352226
rect 402874 352102 403494 352170
rect 402874 352046 402970 352102
rect 403026 352046 403094 352102
rect 403150 352046 403218 352102
rect 403274 352046 403342 352102
rect 403398 352046 403494 352102
rect 402874 351978 403494 352046
rect 402874 351922 402970 351978
rect 403026 351922 403094 351978
rect 403150 351922 403218 351978
rect 403274 351922 403342 351978
rect 403398 351922 403494 351978
rect 402874 334350 403494 351922
rect 402874 334294 402970 334350
rect 403026 334294 403094 334350
rect 403150 334294 403218 334350
rect 403274 334294 403342 334350
rect 403398 334294 403494 334350
rect 402874 334226 403494 334294
rect 402874 334170 402970 334226
rect 403026 334170 403094 334226
rect 403150 334170 403218 334226
rect 403274 334170 403342 334226
rect 403398 334170 403494 334226
rect 402874 334102 403494 334170
rect 402874 334046 402970 334102
rect 403026 334046 403094 334102
rect 403150 334046 403218 334102
rect 403274 334046 403342 334102
rect 403398 334046 403494 334102
rect 402874 333978 403494 334046
rect 402874 333922 402970 333978
rect 403026 333922 403094 333978
rect 403150 333922 403218 333978
rect 403274 333922 403342 333978
rect 403398 333922 403494 333978
rect 402874 316350 403494 333922
rect 579154 454350 579774 471922
rect 579154 454294 579250 454350
rect 579306 454294 579374 454350
rect 579430 454294 579498 454350
rect 579554 454294 579622 454350
rect 579678 454294 579774 454350
rect 579154 454226 579774 454294
rect 579154 454170 579250 454226
rect 579306 454170 579374 454226
rect 579430 454170 579498 454226
rect 579554 454170 579622 454226
rect 579678 454170 579774 454226
rect 579154 454102 579774 454170
rect 579154 454046 579250 454102
rect 579306 454046 579374 454102
rect 579430 454046 579498 454102
rect 579554 454046 579622 454102
rect 579678 454046 579774 454102
rect 579154 453978 579774 454046
rect 579154 453922 579250 453978
rect 579306 453922 579374 453978
rect 579430 453922 579498 453978
rect 579554 453922 579622 453978
rect 579678 453922 579774 453978
rect 579154 436350 579774 453922
rect 579154 436294 579250 436350
rect 579306 436294 579374 436350
rect 579430 436294 579498 436350
rect 579554 436294 579622 436350
rect 579678 436294 579774 436350
rect 579154 436226 579774 436294
rect 579154 436170 579250 436226
rect 579306 436170 579374 436226
rect 579430 436170 579498 436226
rect 579554 436170 579622 436226
rect 579678 436170 579774 436226
rect 579154 436102 579774 436170
rect 579154 436046 579250 436102
rect 579306 436046 579374 436102
rect 579430 436046 579498 436102
rect 579554 436046 579622 436102
rect 579678 436046 579774 436102
rect 579154 435978 579774 436046
rect 579154 435922 579250 435978
rect 579306 435922 579374 435978
rect 579430 435922 579498 435978
rect 579554 435922 579622 435978
rect 579678 435922 579774 435978
rect 579154 418350 579774 435922
rect 579154 418294 579250 418350
rect 579306 418294 579374 418350
rect 579430 418294 579498 418350
rect 579554 418294 579622 418350
rect 579678 418294 579774 418350
rect 579154 418226 579774 418294
rect 579154 418170 579250 418226
rect 579306 418170 579374 418226
rect 579430 418170 579498 418226
rect 579554 418170 579622 418226
rect 579678 418170 579774 418226
rect 579154 418102 579774 418170
rect 579154 418046 579250 418102
rect 579306 418046 579374 418102
rect 579430 418046 579498 418102
rect 579554 418046 579622 418102
rect 579678 418046 579774 418102
rect 579154 417978 579774 418046
rect 579154 417922 579250 417978
rect 579306 417922 579374 417978
rect 579430 417922 579498 417978
rect 579554 417922 579622 417978
rect 579678 417922 579774 417978
rect 579154 400350 579774 417922
rect 579154 400294 579250 400350
rect 579306 400294 579374 400350
rect 579430 400294 579498 400350
rect 579554 400294 579622 400350
rect 579678 400294 579774 400350
rect 579154 400226 579774 400294
rect 579154 400170 579250 400226
rect 579306 400170 579374 400226
rect 579430 400170 579498 400226
rect 579554 400170 579622 400226
rect 579678 400170 579774 400226
rect 579154 400102 579774 400170
rect 579154 400046 579250 400102
rect 579306 400046 579374 400102
rect 579430 400046 579498 400102
rect 579554 400046 579622 400102
rect 579678 400046 579774 400102
rect 579154 399978 579774 400046
rect 579154 399922 579250 399978
rect 579306 399922 579374 399978
rect 579430 399922 579498 399978
rect 579554 399922 579622 399978
rect 579678 399922 579774 399978
rect 579154 382350 579774 399922
rect 579154 382294 579250 382350
rect 579306 382294 579374 382350
rect 579430 382294 579498 382350
rect 579554 382294 579622 382350
rect 579678 382294 579774 382350
rect 579154 382226 579774 382294
rect 579154 382170 579250 382226
rect 579306 382170 579374 382226
rect 579430 382170 579498 382226
rect 579554 382170 579622 382226
rect 579678 382170 579774 382226
rect 579154 382102 579774 382170
rect 579154 382046 579250 382102
rect 579306 382046 579374 382102
rect 579430 382046 579498 382102
rect 579554 382046 579622 382102
rect 579678 382046 579774 382102
rect 579154 381978 579774 382046
rect 579154 381922 579250 381978
rect 579306 381922 579374 381978
rect 579430 381922 579498 381978
rect 579554 381922 579622 381978
rect 579678 381922 579774 381978
rect 579154 364350 579774 381922
rect 579154 364294 579250 364350
rect 579306 364294 579374 364350
rect 579430 364294 579498 364350
rect 579554 364294 579622 364350
rect 579678 364294 579774 364350
rect 579154 364226 579774 364294
rect 579154 364170 579250 364226
rect 579306 364170 579374 364226
rect 579430 364170 579498 364226
rect 579554 364170 579622 364226
rect 579678 364170 579774 364226
rect 579154 364102 579774 364170
rect 579154 364046 579250 364102
rect 579306 364046 579374 364102
rect 579430 364046 579498 364102
rect 579554 364046 579622 364102
rect 579678 364046 579774 364102
rect 579154 363978 579774 364046
rect 579154 363922 579250 363978
rect 579306 363922 579374 363978
rect 579430 363922 579498 363978
rect 579554 363922 579622 363978
rect 579678 363922 579774 363978
rect 579154 346350 579774 363922
rect 579154 346294 579250 346350
rect 579306 346294 579374 346350
rect 579430 346294 579498 346350
rect 579554 346294 579622 346350
rect 579678 346294 579774 346350
rect 579154 346226 579774 346294
rect 579154 346170 579250 346226
rect 579306 346170 579374 346226
rect 579430 346170 579498 346226
rect 579554 346170 579622 346226
rect 579678 346170 579774 346226
rect 579154 346102 579774 346170
rect 579154 346046 579250 346102
rect 579306 346046 579374 346102
rect 579430 346046 579498 346102
rect 579554 346046 579622 346102
rect 579678 346046 579774 346102
rect 579154 345978 579774 346046
rect 579154 345922 579250 345978
rect 579306 345922 579374 345978
rect 579430 345922 579498 345978
rect 579554 345922 579622 345978
rect 579678 345922 579774 345978
rect 579154 328350 579774 345922
rect 579154 328294 579250 328350
rect 579306 328294 579374 328350
rect 579430 328294 579498 328350
rect 579554 328294 579622 328350
rect 579678 328294 579774 328350
rect 579154 328226 579774 328294
rect 579154 328170 579250 328226
rect 579306 328170 579374 328226
rect 579430 328170 579498 328226
rect 579554 328170 579622 328226
rect 579678 328170 579774 328226
rect 579154 328102 579774 328170
rect 579154 328046 579250 328102
rect 579306 328046 579374 328102
rect 579430 328046 579498 328102
rect 579554 328046 579622 328102
rect 579678 328046 579774 328102
rect 579154 327978 579774 328046
rect 579154 327922 579250 327978
rect 579306 327922 579374 327978
rect 579430 327922 579498 327978
rect 579554 327922 579622 327978
rect 579678 327922 579774 327978
rect 402874 316294 402970 316350
rect 403026 316294 403094 316350
rect 403150 316294 403218 316350
rect 403274 316294 403342 316350
rect 403398 316294 403494 316350
rect 402874 316226 403494 316294
rect 402874 316170 402970 316226
rect 403026 316170 403094 316226
rect 403150 316170 403218 316226
rect 403274 316170 403342 316226
rect 403398 316170 403494 316226
rect 402874 316102 403494 316170
rect 402874 316046 402970 316102
rect 403026 316046 403094 316102
rect 403150 316046 403218 316102
rect 403274 316046 403342 316102
rect 403398 316046 403494 316102
rect 402874 315978 403494 316046
rect 402874 315922 402970 315978
rect 403026 315922 403094 315978
rect 403150 315922 403218 315978
rect 403274 315922 403342 315978
rect 403398 315922 403494 315978
rect 402874 298350 403494 315922
rect 402874 298294 402970 298350
rect 403026 298294 403094 298350
rect 403150 298294 403218 298350
rect 403274 298294 403342 298350
rect 403398 298294 403494 298350
rect 420874 316350 421494 318858
rect 420874 316294 420970 316350
rect 421026 316294 421094 316350
rect 421150 316294 421218 316350
rect 421274 316294 421342 316350
rect 421398 316294 421494 316350
rect 420874 316226 421494 316294
rect 420874 316170 420970 316226
rect 421026 316170 421094 316226
rect 421150 316170 421218 316226
rect 421274 316170 421342 316226
rect 421398 316170 421494 316226
rect 420874 316102 421494 316170
rect 420874 316046 420970 316102
rect 421026 316046 421094 316102
rect 421150 316046 421218 316102
rect 421274 316046 421342 316102
rect 421398 316046 421494 316102
rect 420874 315978 421494 316046
rect 420874 315922 420970 315978
rect 421026 315922 421094 315978
rect 421150 315922 421218 315978
rect 421274 315922 421342 315978
rect 421398 315922 421494 315978
rect 420874 298422 421494 315922
rect 420874 298366 420970 298422
rect 421026 298366 421094 298422
rect 421150 298366 421218 298422
rect 421274 298366 421342 298422
rect 421398 298366 421494 298422
rect 420874 298342 421494 298366
rect 438874 316350 439494 318858
rect 438874 316294 438970 316350
rect 439026 316294 439094 316350
rect 439150 316294 439218 316350
rect 439274 316294 439342 316350
rect 439398 316294 439494 316350
rect 438874 316226 439494 316294
rect 438874 316170 438970 316226
rect 439026 316170 439094 316226
rect 439150 316170 439218 316226
rect 439274 316170 439342 316226
rect 439398 316170 439494 316226
rect 438874 316102 439494 316170
rect 438874 316046 438970 316102
rect 439026 316046 439094 316102
rect 439150 316046 439218 316102
rect 439274 316046 439342 316102
rect 439398 316046 439494 316102
rect 438874 315978 439494 316046
rect 438874 315922 438970 315978
rect 439026 315922 439094 315978
rect 439150 315922 439218 315978
rect 439274 315922 439342 315978
rect 439398 315922 439494 315978
rect 438874 298422 439494 315922
rect 438874 298366 438970 298422
rect 439026 298366 439094 298422
rect 439150 298366 439218 298422
rect 439274 298366 439342 298422
rect 439398 298366 439494 298422
rect 438874 298342 439494 298366
rect 456874 316350 457494 318858
rect 456874 316294 456970 316350
rect 457026 316294 457094 316350
rect 457150 316294 457218 316350
rect 457274 316294 457342 316350
rect 457398 316294 457494 316350
rect 456874 316226 457494 316294
rect 456874 316170 456970 316226
rect 457026 316170 457094 316226
rect 457150 316170 457218 316226
rect 457274 316170 457342 316226
rect 457398 316170 457494 316226
rect 456874 316102 457494 316170
rect 456874 316046 456970 316102
rect 457026 316046 457094 316102
rect 457150 316046 457218 316102
rect 457274 316046 457342 316102
rect 457398 316046 457494 316102
rect 456874 315978 457494 316046
rect 456874 315922 456970 315978
rect 457026 315922 457094 315978
rect 457150 315922 457218 315978
rect 457274 315922 457342 315978
rect 457398 315922 457494 315978
rect 456874 298422 457494 315922
rect 456874 298366 456970 298422
rect 457026 298366 457094 298422
rect 457150 298366 457218 298422
rect 457274 298366 457342 298422
rect 457398 298366 457494 298422
rect 456874 298342 457494 298366
rect 474874 316350 475494 318858
rect 474874 316294 474970 316350
rect 475026 316294 475094 316350
rect 475150 316294 475218 316350
rect 475274 316294 475342 316350
rect 475398 316294 475494 316350
rect 474874 316226 475494 316294
rect 474874 316170 474970 316226
rect 475026 316170 475094 316226
rect 475150 316170 475218 316226
rect 475274 316170 475342 316226
rect 475398 316170 475494 316226
rect 474874 316102 475494 316170
rect 474874 316046 474970 316102
rect 475026 316046 475094 316102
rect 475150 316046 475218 316102
rect 475274 316046 475342 316102
rect 475398 316046 475494 316102
rect 474874 315978 475494 316046
rect 474874 315922 474970 315978
rect 475026 315922 475094 315978
rect 475150 315922 475218 315978
rect 475274 315922 475342 315978
rect 475398 315922 475494 315978
rect 474874 298422 475494 315922
rect 474874 298366 474970 298422
rect 475026 298366 475094 298422
rect 475150 298366 475218 298422
rect 475274 298366 475342 298422
rect 475398 298366 475494 298422
rect 474874 298342 475494 298366
rect 492874 316350 493494 318858
rect 492874 316294 492970 316350
rect 493026 316294 493094 316350
rect 493150 316294 493218 316350
rect 493274 316294 493342 316350
rect 493398 316294 493494 316350
rect 492874 316226 493494 316294
rect 492874 316170 492970 316226
rect 493026 316170 493094 316226
rect 493150 316170 493218 316226
rect 493274 316170 493342 316226
rect 493398 316170 493494 316226
rect 492874 316102 493494 316170
rect 492874 316046 492970 316102
rect 493026 316046 493094 316102
rect 493150 316046 493218 316102
rect 493274 316046 493342 316102
rect 493398 316046 493494 316102
rect 492874 315978 493494 316046
rect 492874 315922 492970 315978
rect 493026 315922 493094 315978
rect 493150 315922 493218 315978
rect 493274 315922 493342 315978
rect 493398 315922 493494 315978
rect 492874 298422 493494 315922
rect 492874 298366 492970 298422
rect 493026 298366 493094 298422
rect 493150 298366 493218 298422
rect 493274 298366 493342 298422
rect 493398 298366 493494 298422
rect 492874 298342 493494 298366
rect 510874 316350 511494 318858
rect 510874 316294 510970 316350
rect 511026 316294 511094 316350
rect 511150 316294 511218 316350
rect 511274 316294 511342 316350
rect 511398 316294 511494 316350
rect 510874 316226 511494 316294
rect 510874 316170 510970 316226
rect 511026 316170 511094 316226
rect 511150 316170 511218 316226
rect 511274 316170 511342 316226
rect 511398 316170 511494 316226
rect 510874 316102 511494 316170
rect 510874 316046 510970 316102
rect 511026 316046 511094 316102
rect 511150 316046 511218 316102
rect 511274 316046 511342 316102
rect 511398 316046 511494 316102
rect 510874 315978 511494 316046
rect 510874 315922 510970 315978
rect 511026 315922 511094 315978
rect 511150 315922 511218 315978
rect 511274 315922 511342 315978
rect 511398 315922 511494 315978
rect 510874 298422 511494 315922
rect 510874 298366 510970 298422
rect 511026 298366 511094 298422
rect 511150 298366 511218 298422
rect 511274 298366 511342 298422
rect 511398 298366 511494 298422
rect 510874 298342 511494 298366
rect 528874 316350 529494 318858
rect 528874 316294 528970 316350
rect 529026 316294 529094 316350
rect 529150 316294 529218 316350
rect 529274 316294 529342 316350
rect 529398 316294 529494 316350
rect 528874 316226 529494 316294
rect 528874 316170 528970 316226
rect 529026 316170 529094 316226
rect 529150 316170 529218 316226
rect 529274 316170 529342 316226
rect 529398 316170 529494 316226
rect 528874 316102 529494 316170
rect 528874 316046 528970 316102
rect 529026 316046 529094 316102
rect 529150 316046 529218 316102
rect 529274 316046 529342 316102
rect 529398 316046 529494 316102
rect 528874 315978 529494 316046
rect 528874 315922 528970 315978
rect 529026 315922 529094 315978
rect 529150 315922 529218 315978
rect 529274 315922 529342 315978
rect 529398 315922 529494 315978
rect 528874 298422 529494 315922
rect 528874 298366 528970 298422
rect 529026 298366 529094 298422
rect 529150 298366 529218 298422
rect 529274 298366 529342 298422
rect 529398 298366 529494 298422
rect 528874 298342 529494 298366
rect 546874 316350 547494 318858
rect 546874 316294 546970 316350
rect 547026 316294 547094 316350
rect 547150 316294 547218 316350
rect 547274 316294 547342 316350
rect 547398 316294 547494 316350
rect 546874 316226 547494 316294
rect 546874 316170 546970 316226
rect 547026 316170 547094 316226
rect 547150 316170 547218 316226
rect 547274 316170 547342 316226
rect 547398 316170 547494 316226
rect 546874 316102 547494 316170
rect 546874 316046 546970 316102
rect 547026 316046 547094 316102
rect 547150 316046 547218 316102
rect 547274 316046 547342 316102
rect 547398 316046 547494 316102
rect 546874 315978 547494 316046
rect 546874 315922 546970 315978
rect 547026 315922 547094 315978
rect 547150 315922 547218 315978
rect 547274 315922 547342 315978
rect 547398 315922 547494 315978
rect 546874 298422 547494 315922
rect 546874 298366 546970 298422
rect 547026 298366 547094 298422
rect 547150 298366 547218 298422
rect 547274 298366 547342 298422
rect 547398 298366 547494 298422
rect 546874 298342 547494 298366
rect 564874 316350 565494 318858
rect 564874 316294 564970 316350
rect 565026 316294 565094 316350
rect 565150 316294 565218 316350
rect 565274 316294 565342 316350
rect 565398 316294 565494 316350
rect 564874 316226 565494 316294
rect 564874 316170 564970 316226
rect 565026 316170 565094 316226
rect 565150 316170 565218 316226
rect 565274 316170 565342 316226
rect 565398 316170 565494 316226
rect 564874 316102 565494 316170
rect 564874 316046 564970 316102
rect 565026 316046 565094 316102
rect 565150 316046 565218 316102
rect 565274 316046 565342 316102
rect 565398 316046 565494 316102
rect 564874 315978 565494 316046
rect 564874 315922 564970 315978
rect 565026 315922 565094 315978
rect 565150 315922 565218 315978
rect 565274 315922 565342 315978
rect 565398 315922 565494 315978
rect 564874 298422 565494 315922
rect 564874 298366 564970 298422
rect 565026 298366 565094 298422
rect 565150 298366 565218 298422
rect 565274 298366 565342 298422
rect 565398 298366 565494 298422
rect 564874 298342 565494 298366
rect 579154 310350 579774 327922
rect 579154 310294 579250 310350
rect 579306 310294 579374 310350
rect 579430 310294 579498 310350
rect 579554 310294 579622 310350
rect 579678 310294 579774 310350
rect 579154 310226 579774 310294
rect 579154 310170 579250 310226
rect 579306 310170 579374 310226
rect 579430 310170 579498 310226
rect 579554 310170 579622 310226
rect 579678 310170 579774 310226
rect 579154 310102 579774 310170
rect 579154 310046 579250 310102
rect 579306 310046 579374 310102
rect 579430 310046 579498 310102
rect 579554 310046 579622 310102
rect 579678 310046 579774 310102
rect 579154 309978 579774 310046
rect 579154 309922 579250 309978
rect 579306 309922 579374 309978
rect 579430 309922 579498 309978
rect 579554 309922 579622 309978
rect 579678 309922 579774 309978
rect 402874 298226 403494 298294
rect 402874 298170 402970 298226
rect 403026 298170 403094 298226
rect 403150 298170 403218 298226
rect 403274 298170 403342 298226
rect 403398 298170 403494 298226
rect 402874 298102 403494 298170
rect 402874 298046 402970 298102
rect 403026 298046 403094 298102
rect 403150 298046 403218 298102
rect 403274 298046 403342 298102
rect 403398 298046 403494 298102
rect 402874 297978 403494 298046
rect 402874 297922 402970 297978
rect 403026 297922 403094 297978
rect 403150 297922 403218 297978
rect 403274 297922 403342 297978
rect 403398 297922 403494 297978
rect 402874 280350 403494 297922
rect 402874 280294 402970 280350
rect 403026 280294 403094 280350
rect 403150 280294 403218 280350
rect 403274 280294 403342 280350
rect 403398 280294 403494 280350
rect 402874 280226 403494 280294
rect 402874 280170 402970 280226
rect 403026 280170 403094 280226
rect 403150 280170 403218 280226
rect 403274 280170 403342 280226
rect 403398 280170 403494 280226
rect 402874 280102 403494 280170
rect 402874 280046 402970 280102
rect 403026 280046 403094 280102
rect 403150 280046 403218 280102
rect 403274 280046 403342 280102
rect 403398 280046 403494 280102
rect 402874 279978 403494 280046
rect 402874 279922 402970 279978
rect 403026 279922 403094 279978
rect 403150 279922 403218 279978
rect 403274 279922 403342 279978
rect 403398 279922 403494 279978
rect 402874 262350 403494 279922
rect 402874 262294 402970 262350
rect 403026 262294 403094 262350
rect 403150 262294 403218 262350
rect 403274 262294 403342 262350
rect 403398 262294 403494 262350
rect 402874 262226 403494 262294
rect 402874 262170 402970 262226
rect 403026 262170 403094 262226
rect 403150 262170 403218 262226
rect 403274 262170 403342 262226
rect 403398 262170 403494 262226
rect 402874 262102 403494 262170
rect 402874 262046 402970 262102
rect 403026 262046 403094 262102
rect 403150 262046 403218 262102
rect 403274 262046 403342 262102
rect 403398 262046 403494 262102
rect 402874 261978 403494 262046
rect 402874 261922 402970 261978
rect 403026 261922 403094 261978
rect 403150 261922 403218 261978
rect 403274 261922 403342 261978
rect 403398 261922 403494 261978
rect 402874 244350 403494 261922
rect 402874 244294 402970 244350
rect 403026 244294 403094 244350
rect 403150 244294 403218 244350
rect 403274 244294 403342 244350
rect 403398 244294 403494 244350
rect 402874 244226 403494 244294
rect 402874 244170 402970 244226
rect 403026 244170 403094 244226
rect 403150 244170 403218 244226
rect 403274 244170 403342 244226
rect 403398 244170 403494 244226
rect 402874 244102 403494 244170
rect 402874 244046 402970 244102
rect 403026 244046 403094 244102
rect 403150 244046 403218 244102
rect 403274 244046 403342 244102
rect 403398 244046 403494 244102
rect 402874 243978 403494 244046
rect 402874 243922 402970 243978
rect 403026 243922 403094 243978
rect 403150 243922 403218 243978
rect 403274 243922 403342 243978
rect 403398 243922 403494 243978
rect 402874 226350 403494 243922
rect 402874 226294 402970 226350
rect 403026 226294 403094 226350
rect 403150 226294 403218 226350
rect 403274 226294 403342 226350
rect 403398 226294 403494 226350
rect 402874 226226 403494 226294
rect 402874 226170 402970 226226
rect 403026 226170 403094 226226
rect 403150 226170 403218 226226
rect 403274 226170 403342 226226
rect 403398 226170 403494 226226
rect 402874 226102 403494 226170
rect 402874 226046 402970 226102
rect 403026 226046 403094 226102
rect 403150 226046 403218 226102
rect 403274 226046 403342 226102
rect 403398 226046 403494 226102
rect 402874 225978 403494 226046
rect 402874 225922 402970 225978
rect 403026 225922 403094 225978
rect 403150 225922 403218 225978
rect 403274 225922 403342 225978
rect 403398 225922 403494 225978
rect 402874 208350 403494 225922
rect 402874 208294 402970 208350
rect 403026 208294 403094 208350
rect 403150 208294 403218 208350
rect 403274 208294 403342 208350
rect 403398 208294 403494 208350
rect 402874 208226 403494 208294
rect 402874 208170 402970 208226
rect 403026 208170 403094 208226
rect 403150 208170 403218 208226
rect 403274 208170 403342 208226
rect 403398 208170 403494 208226
rect 402874 208102 403494 208170
rect 402874 208046 402970 208102
rect 403026 208046 403094 208102
rect 403150 208046 403218 208102
rect 403274 208046 403342 208102
rect 403398 208046 403494 208102
rect 402874 207978 403494 208046
rect 402874 207922 402970 207978
rect 403026 207922 403094 207978
rect 403150 207922 403218 207978
rect 403274 207922 403342 207978
rect 403398 207922 403494 207978
rect 402874 190350 403494 207922
rect 402874 190294 402970 190350
rect 403026 190294 403094 190350
rect 403150 190294 403218 190350
rect 403274 190294 403342 190350
rect 403398 190294 403494 190350
rect 402874 190226 403494 190294
rect 402874 190170 402970 190226
rect 403026 190170 403094 190226
rect 403150 190170 403218 190226
rect 403274 190170 403342 190226
rect 403398 190170 403494 190226
rect 402874 190102 403494 190170
rect 402874 190046 402970 190102
rect 403026 190046 403094 190102
rect 403150 190046 403218 190102
rect 403274 190046 403342 190102
rect 403398 190046 403494 190102
rect 402874 189978 403494 190046
rect 402874 189922 402970 189978
rect 403026 189922 403094 189978
rect 403150 189922 403218 189978
rect 403274 189922 403342 189978
rect 403398 189922 403494 189978
rect 402874 172350 403494 189922
rect 402874 172294 402970 172350
rect 403026 172294 403094 172350
rect 403150 172294 403218 172350
rect 403274 172294 403342 172350
rect 403398 172294 403494 172350
rect 402874 172226 403494 172294
rect 402874 172170 402970 172226
rect 403026 172170 403094 172226
rect 403150 172170 403218 172226
rect 403274 172170 403342 172226
rect 403398 172170 403494 172226
rect 402874 172102 403494 172170
rect 402874 172046 402970 172102
rect 403026 172046 403094 172102
rect 403150 172046 403218 172102
rect 403274 172046 403342 172102
rect 403398 172046 403494 172102
rect 402874 171978 403494 172046
rect 402874 171922 402970 171978
rect 403026 171922 403094 171978
rect 403150 171922 403218 171978
rect 403274 171922 403342 171978
rect 403398 171922 403494 171978
rect 402874 154350 403494 171922
rect 579154 292350 579774 309922
rect 579154 292294 579250 292350
rect 579306 292294 579374 292350
rect 579430 292294 579498 292350
rect 579554 292294 579622 292350
rect 579678 292294 579774 292350
rect 579154 292226 579774 292294
rect 579154 292170 579250 292226
rect 579306 292170 579374 292226
rect 579430 292170 579498 292226
rect 579554 292170 579622 292226
rect 579678 292170 579774 292226
rect 579154 292102 579774 292170
rect 579154 292046 579250 292102
rect 579306 292046 579374 292102
rect 579430 292046 579498 292102
rect 579554 292046 579622 292102
rect 579678 292046 579774 292102
rect 579154 291978 579774 292046
rect 579154 291922 579250 291978
rect 579306 291922 579374 291978
rect 579430 291922 579498 291978
rect 579554 291922 579622 291978
rect 579678 291922 579774 291978
rect 579154 274350 579774 291922
rect 579154 274294 579250 274350
rect 579306 274294 579374 274350
rect 579430 274294 579498 274350
rect 579554 274294 579622 274350
rect 579678 274294 579774 274350
rect 579154 274226 579774 274294
rect 579154 274170 579250 274226
rect 579306 274170 579374 274226
rect 579430 274170 579498 274226
rect 579554 274170 579622 274226
rect 579678 274170 579774 274226
rect 579154 274102 579774 274170
rect 579154 274046 579250 274102
rect 579306 274046 579374 274102
rect 579430 274046 579498 274102
rect 579554 274046 579622 274102
rect 579678 274046 579774 274102
rect 579154 273978 579774 274046
rect 579154 273922 579250 273978
rect 579306 273922 579374 273978
rect 579430 273922 579498 273978
rect 579554 273922 579622 273978
rect 579678 273922 579774 273978
rect 579154 256350 579774 273922
rect 579154 256294 579250 256350
rect 579306 256294 579374 256350
rect 579430 256294 579498 256350
rect 579554 256294 579622 256350
rect 579678 256294 579774 256350
rect 579154 256226 579774 256294
rect 579154 256170 579250 256226
rect 579306 256170 579374 256226
rect 579430 256170 579498 256226
rect 579554 256170 579622 256226
rect 579678 256170 579774 256226
rect 579154 256102 579774 256170
rect 579154 256046 579250 256102
rect 579306 256046 579374 256102
rect 579430 256046 579498 256102
rect 579554 256046 579622 256102
rect 579678 256046 579774 256102
rect 579154 255978 579774 256046
rect 579154 255922 579250 255978
rect 579306 255922 579374 255978
rect 579430 255922 579498 255978
rect 579554 255922 579622 255978
rect 579678 255922 579774 255978
rect 579154 238350 579774 255922
rect 579154 238294 579250 238350
rect 579306 238294 579374 238350
rect 579430 238294 579498 238350
rect 579554 238294 579622 238350
rect 579678 238294 579774 238350
rect 579154 238226 579774 238294
rect 579154 238170 579250 238226
rect 579306 238170 579374 238226
rect 579430 238170 579498 238226
rect 579554 238170 579622 238226
rect 579678 238170 579774 238226
rect 579154 238102 579774 238170
rect 579154 238046 579250 238102
rect 579306 238046 579374 238102
rect 579430 238046 579498 238102
rect 579554 238046 579622 238102
rect 579678 238046 579774 238102
rect 579154 237978 579774 238046
rect 579154 237922 579250 237978
rect 579306 237922 579374 237978
rect 579430 237922 579498 237978
rect 579554 237922 579622 237978
rect 579678 237922 579774 237978
rect 579154 220350 579774 237922
rect 579154 220294 579250 220350
rect 579306 220294 579374 220350
rect 579430 220294 579498 220350
rect 579554 220294 579622 220350
rect 579678 220294 579774 220350
rect 579154 220226 579774 220294
rect 579154 220170 579250 220226
rect 579306 220170 579374 220226
rect 579430 220170 579498 220226
rect 579554 220170 579622 220226
rect 579678 220170 579774 220226
rect 579154 220102 579774 220170
rect 579154 220046 579250 220102
rect 579306 220046 579374 220102
rect 579430 220046 579498 220102
rect 579554 220046 579622 220102
rect 579678 220046 579774 220102
rect 579154 219978 579774 220046
rect 579154 219922 579250 219978
rect 579306 219922 579374 219978
rect 579430 219922 579498 219978
rect 579554 219922 579622 219978
rect 579678 219922 579774 219978
rect 579154 202350 579774 219922
rect 579154 202294 579250 202350
rect 579306 202294 579374 202350
rect 579430 202294 579498 202350
rect 579554 202294 579622 202350
rect 579678 202294 579774 202350
rect 579154 202226 579774 202294
rect 579154 202170 579250 202226
rect 579306 202170 579374 202226
rect 579430 202170 579498 202226
rect 579554 202170 579622 202226
rect 579678 202170 579774 202226
rect 579154 202102 579774 202170
rect 579154 202046 579250 202102
rect 579306 202046 579374 202102
rect 579430 202046 579498 202102
rect 579554 202046 579622 202102
rect 579678 202046 579774 202102
rect 579154 201978 579774 202046
rect 579154 201922 579250 201978
rect 579306 201922 579374 201978
rect 579430 201922 579498 201978
rect 579554 201922 579622 201978
rect 579678 201922 579774 201978
rect 579154 184350 579774 201922
rect 579154 184294 579250 184350
rect 579306 184294 579374 184350
rect 579430 184294 579498 184350
rect 579554 184294 579622 184350
rect 579678 184294 579774 184350
rect 579154 184226 579774 184294
rect 579154 184170 579250 184226
rect 579306 184170 579374 184226
rect 579430 184170 579498 184226
rect 579554 184170 579622 184226
rect 579678 184170 579774 184226
rect 579154 184102 579774 184170
rect 579154 184046 579250 184102
rect 579306 184046 579374 184102
rect 579430 184046 579498 184102
rect 579554 184046 579622 184102
rect 579678 184046 579774 184102
rect 579154 183978 579774 184046
rect 579154 183922 579250 183978
rect 579306 183922 579374 183978
rect 579430 183922 579498 183978
rect 579554 183922 579622 183978
rect 579678 183922 579774 183978
rect 579154 166350 579774 183922
rect 579154 166294 579250 166350
rect 579306 166294 579374 166350
rect 579430 166294 579498 166350
rect 579554 166294 579622 166350
rect 579678 166294 579774 166350
rect 579154 166226 579774 166294
rect 579154 166170 579250 166226
rect 579306 166170 579374 166226
rect 579430 166170 579498 166226
rect 579554 166170 579622 166226
rect 579678 166170 579774 166226
rect 579154 166102 579774 166170
rect 579154 166046 579250 166102
rect 579306 166046 579374 166102
rect 579430 166046 579498 166102
rect 579554 166046 579622 166102
rect 579678 166046 579774 166102
rect 579154 165978 579774 166046
rect 579154 165922 579250 165978
rect 579306 165922 579374 165978
rect 579430 165922 579498 165978
rect 579554 165922 579622 165978
rect 579678 165922 579774 165978
rect 402874 154294 402970 154350
rect 403026 154294 403094 154350
rect 403150 154294 403218 154350
rect 403274 154294 403342 154350
rect 403398 154294 403494 154350
rect 402874 154226 403494 154294
rect 402874 154170 402970 154226
rect 403026 154170 403094 154226
rect 403150 154170 403218 154226
rect 403274 154170 403342 154226
rect 403398 154170 403494 154226
rect 402874 154102 403494 154170
rect 402874 154046 402970 154102
rect 403026 154046 403094 154102
rect 403150 154046 403218 154102
rect 403274 154046 403342 154102
rect 403398 154046 403494 154102
rect 402874 153978 403494 154046
rect 402874 153922 402970 153978
rect 403026 153922 403094 153978
rect 403150 153922 403218 153978
rect 403274 153922 403342 153978
rect 403398 153922 403494 153978
rect 402874 136350 403494 153922
rect 402874 136294 402970 136350
rect 403026 136294 403094 136350
rect 403150 136294 403218 136350
rect 403274 136294 403342 136350
rect 403398 136294 403494 136350
rect 402874 136226 403494 136294
rect 402874 136170 402970 136226
rect 403026 136170 403094 136226
rect 403150 136170 403218 136226
rect 403274 136170 403342 136226
rect 403398 136170 403494 136226
rect 402874 136102 403494 136170
rect 402874 136046 402970 136102
rect 403026 136046 403094 136102
rect 403150 136046 403218 136102
rect 403274 136046 403342 136102
rect 403398 136046 403494 136102
rect 402874 135978 403494 136046
rect 402874 135922 402970 135978
rect 403026 135922 403094 135978
rect 403150 135922 403218 135978
rect 403274 135922 403342 135978
rect 403398 135922 403494 135978
rect 402874 118350 403494 135922
rect 402874 118294 402970 118350
rect 403026 118294 403094 118350
rect 403150 118294 403218 118350
rect 403274 118294 403342 118350
rect 403398 118294 403494 118350
rect 402874 118226 403494 118294
rect 402874 118170 402970 118226
rect 403026 118170 403094 118226
rect 403150 118170 403218 118226
rect 403274 118170 403342 118226
rect 403398 118170 403494 118226
rect 402874 118102 403494 118170
rect 402874 118046 402970 118102
rect 403026 118046 403094 118102
rect 403150 118046 403218 118102
rect 403274 118046 403342 118102
rect 403398 118046 403494 118102
rect 402874 117978 403494 118046
rect 402874 117922 402970 117978
rect 403026 117922 403094 117978
rect 403150 117922 403218 117978
rect 403274 117922 403342 117978
rect 403398 117922 403494 117978
rect 402874 100350 403494 117922
rect 402874 100294 402970 100350
rect 403026 100294 403094 100350
rect 403150 100294 403218 100350
rect 403274 100294 403342 100350
rect 403398 100294 403494 100350
rect 402874 100226 403494 100294
rect 402874 100170 402970 100226
rect 403026 100170 403094 100226
rect 403150 100170 403218 100226
rect 403274 100170 403342 100226
rect 403398 100170 403494 100226
rect 402874 100102 403494 100170
rect 402874 100046 402970 100102
rect 403026 100046 403094 100102
rect 403150 100046 403218 100102
rect 403274 100046 403342 100102
rect 403398 100046 403494 100102
rect 402874 99978 403494 100046
rect 402874 99922 402970 99978
rect 403026 99922 403094 99978
rect 403150 99922 403218 99978
rect 403274 99922 403342 99978
rect 403398 99922 403494 99978
rect 402874 82350 403494 99922
rect 402874 82294 402970 82350
rect 403026 82294 403094 82350
rect 403150 82294 403218 82350
rect 403274 82294 403342 82350
rect 403398 82294 403494 82350
rect 402874 82226 403494 82294
rect 402874 82170 402970 82226
rect 403026 82170 403094 82226
rect 403150 82170 403218 82226
rect 403274 82170 403342 82226
rect 403398 82170 403494 82226
rect 402874 82102 403494 82170
rect 402874 82046 402970 82102
rect 403026 82046 403094 82102
rect 403150 82046 403218 82102
rect 403274 82046 403342 82102
rect 403398 82046 403494 82102
rect 402874 81978 403494 82046
rect 402874 81922 402970 81978
rect 403026 81922 403094 81978
rect 403150 81922 403218 81978
rect 403274 81922 403342 81978
rect 403398 81922 403494 81978
rect 402874 64350 403494 81922
rect 402874 64294 402970 64350
rect 403026 64294 403094 64350
rect 403150 64294 403218 64350
rect 403274 64294 403342 64350
rect 403398 64294 403494 64350
rect 402874 64226 403494 64294
rect 402874 64170 402970 64226
rect 403026 64170 403094 64226
rect 403150 64170 403218 64226
rect 403274 64170 403342 64226
rect 403398 64170 403494 64226
rect 402874 64102 403494 64170
rect 402874 64046 402970 64102
rect 403026 64046 403094 64102
rect 403150 64046 403218 64102
rect 403274 64046 403342 64102
rect 403398 64046 403494 64102
rect 402874 63978 403494 64046
rect 402874 63922 402970 63978
rect 403026 63922 403094 63978
rect 403150 63922 403218 63978
rect 403274 63922 403342 63978
rect 403398 63922 403494 63978
rect 402874 46350 403494 63922
rect 402874 46294 402970 46350
rect 403026 46294 403094 46350
rect 403150 46294 403218 46350
rect 403274 46294 403342 46350
rect 403398 46294 403494 46350
rect 402874 46226 403494 46294
rect 402874 46170 402970 46226
rect 403026 46170 403094 46226
rect 403150 46170 403218 46226
rect 403274 46170 403342 46226
rect 403398 46170 403494 46226
rect 402874 46102 403494 46170
rect 402874 46046 402970 46102
rect 403026 46046 403094 46102
rect 403150 46046 403218 46102
rect 403274 46046 403342 46102
rect 403398 46046 403494 46102
rect 402874 45978 403494 46046
rect 402874 45922 402970 45978
rect 403026 45922 403094 45978
rect 403150 45922 403218 45978
rect 403274 45922 403342 45978
rect 403398 45922 403494 45978
rect 402874 28350 403494 45922
rect 402874 28294 402970 28350
rect 403026 28294 403094 28350
rect 403150 28294 403218 28350
rect 403274 28294 403342 28350
rect 403398 28294 403494 28350
rect 402874 28226 403494 28294
rect 402874 28170 402970 28226
rect 403026 28170 403094 28226
rect 403150 28170 403218 28226
rect 403274 28170 403342 28226
rect 403398 28170 403494 28226
rect 402874 28102 403494 28170
rect 402874 28046 402970 28102
rect 403026 28046 403094 28102
rect 403150 28046 403218 28102
rect 403274 28046 403342 28102
rect 403398 28046 403494 28102
rect 402874 27978 403494 28046
rect 402874 27922 402970 27978
rect 403026 27922 403094 27978
rect 403150 27922 403218 27978
rect 403274 27922 403342 27978
rect 403398 27922 403494 27978
rect 402874 10350 403494 27922
rect 402874 10294 402970 10350
rect 403026 10294 403094 10350
rect 403150 10294 403218 10350
rect 403274 10294 403342 10350
rect 403398 10294 403494 10350
rect 402874 10226 403494 10294
rect 402874 10170 402970 10226
rect 403026 10170 403094 10226
rect 403150 10170 403218 10226
rect 403274 10170 403342 10226
rect 403398 10170 403494 10226
rect 402874 10102 403494 10170
rect 402874 10046 402970 10102
rect 403026 10046 403094 10102
rect 403150 10046 403218 10102
rect 403274 10046 403342 10102
rect 403398 10046 403494 10102
rect 402874 9978 403494 10046
rect 402874 9922 402970 9978
rect 403026 9922 403094 9978
rect 403150 9922 403218 9978
rect 403274 9922 403342 9978
rect 403398 9922 403494 9978
rect 402874 -1120 403494 9922
rect 402874 -1176 402970 -1120
rect 403026 -1176 403094 -1120
rect 403150 -1176 403218 -1120
rect 403274 -1176 403342 -1120
rect 403398 -1176 403494 -1120
rect 402874 -1244 403494 -1176
rect 402874 -1300 402970 -1244
rect 403026 -1300 403094 -1244
rect 403150 -1300 403218 -1244
rect 403274 -1300 403342 -1244
rect 403398 -1300 403494 -1244
rect 402874 -1368 403494 -1300
rect 402874 -1424 402970 -1368
rect 403026 -1424 403094 -1368
rect 403150 -1424 403218 -1368
rect 403274 -1424 403342 -1368
rect 403398 -1424 403494 -1368
rect 402874 -1492 403494 -1424
rect 402874 -1548 402970 -1492
rect 403026 -1548 403094 -1492
rect 403150 -1548 403218 -1492
rect 403274 -1548 403342 -1492
rect 403398 -1548 403494 -1492
rect 402874 -1644 403494 -1548
rect 417154 148350 417774 158858
rect 417154 148294 417250 148350
rect 417306 148294 417374 148350
rect 417430 148294 417498 148350
rect 417554 148294 417622 148350
rect 417678 148294 417774 148350
rect 417154 148226 417774 148294
rect 417154 148170 417250 148226
rect 417306 148170 417374 148226
rect 417430 148170 417498 148226
rect 417554 148170 417622 148226
rect 417678 148170 417774 148226
rect 417154 148102 417774 148170
rect 417154 148046 417250 148102
rect 417306 148046 417374 148102
rect 417430 148046 417498 148102
rect 417554 148046 417622 148102
rect 417678 148046 417774 148102
rect 417154 147978 417774 148046
rect 417154 147922 417250 147978
rect 417306 147922 417374 147978
rect 417430 147922 417498 147978
rect 417554 147922 417622 147978
rect 417678 147922 417774 147978
rect 417154 130350 417774 147922
rect 417154 130294 417250 130350
rect 417306 130294 417374 130350
rect 417430 130294 417498 130350
rect 417554 130294 417622 130350
rect 417678 130294 417774 130350
rect 417154 130226 417774 130294
rect 417154 130170 417250 130226
rect 417306 130170 417374 130226
rect 417430 130170 417498 130226
rect 417554 130170 417622 130226
rect 417678 130170 417774 130226
rect 417154 130102 417774 130170
rect 417154 130046 417250 130102
rect 417306 130046 417374 130102
rect 417430 130046 417498 130102
rect 417554 130046 417622 130102
rect 417678 130046 417774 130102
rect 417154 129978 417774 130046
rect 417154 129922 417250 129978
rect 417306 129922 417374 129978
rect 417430 129922 417498 129978
rect 417554 129922 417622 129978
rect 417678 129922 417774 129978
rect 417154 112350 417774 129922
rect 417154 112294 417250 112350
rect 417306 112294 417374 112350
rect 417430 112294 417498 112350
rect 417554 112294 417622 112350
rect 417678 112294 417774 112350
rect 417154 112226 417774 112294
rect 417154 112170 417250 112226
rect 417306 112170 417374 112226
rect 417430 112170 417498 112226
rect 417554 112170 417622 112226
rect 417678 112170 417774 112226
rect 417154 112102 417774 112170
rect 417154 112046 417250 112102
rect 417306 112046 417374 112102
rect 417430 112046 417498 112102
rect 417554 112046 417622 112102
rect 417678 112046 417774 112102
rect 417154 111978 417774 112046
rect 417154 111922 417250 111978
rect 417306 111922 417374 111978
rect 417430 111922 417498 111978
rect 417554 111922 417622 111978
rect 417678 111922 417774 111978
rect 417154 94350 417774 111922
rect 417154 94294 417250 94350
rect 417306 94294 417374 94350
rect 417430 94294 417498 94350
rect 417554 94294 417622 94350
rect 417678 94294 417774 94350
rect 417154 94226 417774 94294
rect 417154 94170 417250 94226
rect 417306 94170 417374 94226
rect 417430 94170 417498 94226
rect 417554 94170 417622 94226
rect 417678 94170 417774 94226
rect 417154 94102 417774 94170
rect 417154 94046 417250 94102
rect 417306 94046 417374 94102
rect 417430 94046 417498 94102
rect 417554 94046 417622 94102
rect 417678 94046 417774 94102
rect 417154 93978 417774 94046
rect 417154 93922 417250 93978
rect 417306 93922 417374 93978
rect 417430 93922 417498 93978
rect 417554 93922 417622 93978
rect 417678 93922 417774 93978
rect 417154 76350 417774 93922
rect 417154 76294 417250 76350
rect 417306 76294 417374 76350
rect 417430 76294 417498 76350
rect 417554 76294 417622 76350
rect 417678 76294 417774 76350
rect 417154 76226 417774 76294
rect 417154 76170 417250 76226
rect 417306 76170 417374 76226
rect 417430 76170 417498 76226
rect 417554 76170 417622 76226
rect 417678 76170 417774 76226
rect 417154 76102 417774 76170
rect 417154 76046 417250 76102
rect 417306 76046 417374 76102
rect 417430 76046 417498 76102
rect 417554 76046 417622 76102
rect 417678 76046 417774 76102
rect 417154 75978 417774 76046
rect 417154 75922 417250 75978
rect 417306 75922 417374 75978
rect 417430 75922 417498 75978
rect 417554 75922 417622 75978
rect 417678 75922 417774 75978
rect 417154 58350 417774 75922
rect 417154 58294 417250 58350
rect 417306 58294 417374 58350
rect 417430 58294 417498 58350
rect 417554 58294 417622 58350
rect 417678 58294 417774 58350
rect 417154 58226 417774 58294
rect 417154 58170 417250 58226
rect 417306 58170 417374 58226
rect 417430 58170 417498 58226
rect 417554 58170 417622 58226
rect 417678 58170 417774 58226
rect 417154 58102 417774 58170
rect 417154 58046 417250 58102
rect 417306 58046 417374 58102
rect 417430 58046 417498 58102
rect 417554 58046 417622 58102
rect 417678 58046 417774 58102
rect 417154 57978 417774 58046
rect 417154 57922 417250 57978
rect 417306 57922 417374 57978
rect 417430 57922 417498 57978
rect 417554 57922 417622 57978
rect 417678 57922 417774 57978
rect 417154 40350 417774 57922
rect 417154 40294 417250 40350
rect 417306 40294 417374 40350
rect 417430 40294 417498 40350
rect 417554 40294 417622 40350
rect 417678 40294 417774 40350
rect 417154 40226 417774 40294
rect 417154 40170 417250 40226
rect 417306 40170 417374 40226
rect 417430 40170 417498 40226
rect 417554 40170 417622 40226
rect 417678 40170 417774 40226
rect 417154 40102 417774 40170
rect 417154 40046 417250 40102
rect 417306 40046 417374 40102
rect 417430 40046 417498 40102
rect 417554 40046 417622 40102
rect 417678 40046 417774 40102
rect 417154 39978 417774 40046
rect 417154 39922 417250 39978
rect 417306 39922 417374 39978
rect 417430 39922 417498 39978
rect 417554 39922 417622 39978
rect 417678 39922 417774 39978
rect 417154 22350 417774 39922
rect 417154 22294 417250 22350
rect 417306 22294 417374 22350
rect 417430 22294 417498 22350
rect 417554 22294 417622 22350
rect 417678 22294 417774 22350
rect 417154 22226 417774 22294
rect 417154 22170 417250 22226
rect 417306 22170 417374 22226
rect 417430 22170 417498 22226
rect 417554 22170 417622 22226
rect 417678 22170 417774 22226
rect 417154 22102 417774 22170
rect 417154 22046 417250 22102
rect 417306 22046 417374 22102
rect 417430 22046 417498 22102
rect 417554 22046 417622 22102
rect 417678 22046 417774 22102
rect 417154 21978 417774 22046
rect 417154 21922 417250 21978
rect 417306 21922 417374 21978
rect 417430 21922 417498 21978
rect 417554 21922 417622 21978
rect 417678 21922 417774 21978
rect 417154 4350 417774 21922
rect 417154 4294 417250 4350
rect 417306 4294 417374 4350
rect 417430 4294 417498 4350
rect 417554 4294 417622 4350
rect 417678 4294 417774 4350
rect 417154 4226 417774 4294
rect 417154 4170 417250 4226
rect 417306 4170 417374 4226
rect 417430 4170 417498 4226
rect 417554 4170 417622 4226
rect 417678 4170 417774 4226
rect 417154 4102 417774 4170
rect 417154 4046 417250 4102
rect 417306 4046 417374 4102
rect 417430 4046 417498 4102
rect 417554 4046 417622 4102
rect 417678 4046 417774 4102
rect 417154 3978 417774 4046
rect 417154 3922 417250 3978
rect 417306 3922 417374 3978
rect 417430 3922 417498 3978
rect 417554 3922 417622 3978
rect 417678 3922 417774 3978
rect 417154 -160 417774 3922
rect 417154 -216 417250 -160
rect 417306 -216 417374 -160
rect 417430 -216 417498 -160
rect 417554 -216 417622 -160
rect 417678 -216 417774 -160
rect 417154 -284 417774 -216
rect 417154 -340 417250 -284
rect 417306 -340 417374 -284
rect 417430 -340 417498 -284
rect 417554 -340 417622 -284
rect 417678 -340 417774 -284
rect 417154 -408 417774 -340
rect 417154 -464 417250 -408
rect 417306 -464 417374 -408
rect 417430 -464 417498 -408
rect 417554 -464 417622 -408
rect 417678 -464 417774 -408
rect 417154 -532 417774 -464
rect 417154 -588 417250 -532
rect 417306 -588 417374 -532
rect 417430 -588 417498 -532
rect 417554 -588 417622 -532
rect 417678 -588 417774 -532
rect 417154 -1644 417774 -588
rect 420874 154350 421494 158858
rect 420874 154294 420970 154350
rect 421026 154294 421094 154350
rect 421150 154294 421218 154350
rect 421274 154294 421342 154350
rect 421398 154294 421494 154350
rect 420874 154226 421494 154294
rect 420874 154170 420970 154226
rect 421026 154170 421094 154226
rect 421150 154170 421218 154226
rect 421274 154170 421342 154226
rect 421398 154170 421494 154226
rect 420874 154102 421494 154170
rect 420874 154046 420970 154102
rect 421026 154046 421094 154102
rect 421150 154046 421218 154102
rect 421274 154046 421342 154102
rect 421398 154046 421494 154102
rect 420874 153978 421494 154046
rect 420874 153922 420970 153978
rect 421026 153922 421094 153978
rect 421150 153922 421218 153978
rect 421274 153922 421342 153978
rect 421398 153922 421494 153978
rect 420874 136350 421494 153922
rect 420874 136294 420970 136350
rect 421026 136294 421094 136350
rect 421150 136294 421218 136350
rect 421274 136294 421342 136350
rect 421398 136294 421494 136350
rect 420874 136226 421494 136294
rect 420874 136170 420970 136226
rect 421026 136170 421094 136226
rect 421150 136170 421218 136226
rect 421274 136170 421342 136226
rect 421398 136170 421494 136226
rect 420874 136102 421494 136170
rect 420874 136046 420970 136102
rect 421026 136046 421094 136102
rect 421150 136046 421218 136102
rect 421274 136046 421342 136102
rect 421398 136046 421494 136102
rect 420874 135978 421494 136046
rect 420874 135922 420970 135978
rect 421026 135922 421094 135978
rect 421150 135922 421218 135978
rect 421274 135922 421342 135978
rect 421398 135922 421494 135978
rect 420874 118350 421494 135922
rect 420874 118294 420970 118350
rect 421026 118294 421094 118350
rect 421150 118294 421218 118350
rect 421274 118294 421342 118350
rect 421398 118294 421494 118350
rect 420874 118226 421494 118294
rect 420874 118170 420970 118226
rect 421026 118170 421094 118226
rect 421150 118170 421218 118226
rect 421274 118170 421342 118226
rect 421398 118170 421494 118226
rect 420874 118102 421494 118170
rect 420874 118046 420970 118102
rect 421026 118046 421094 118102
rect 421150 118046 421218 118102
rect 421274 118046 421342 118102
rect 421398 118046 421494 118102
rect 420874 117978 421494 118046
rect 420874 117922 420970 117978
rect 421026 117922 421094 117978
rect 421150 117922 421218 117978
rect 421274 117922 421342 117978
rect 421398 117922 421494 117978
rect 420874 100350 421494 117922
rect 420874 100294 420970 100350
rect 421026 100294 421094 100350
rect 421150 100294 421218 100350
rect 421274 100294 421342 100350
rect 421398 100294 421494 100350
rect 420874 100226 421494 100294
rect 420874 100170 420970 100226
rect 421026 100170 421094 100226
rect 421150 100170 421218 100226
rect 421274 100170 421342 100226
rect 421398 100170 421494 100226
rect 420874 100102 421494 100170
rect 420874 100046 420970 100102
rect 421026 100046 421094 100102
rect 421150 100046 421218 100102
rect 421274 100046 421342 100102
rect 421398 100046 421494 100102
rect 420874 99978 421494 100046
rect 420874 99922 420970 99978
rect 421026 99922 421094 99978
rect 421150 99922 421218 99978
rect 421274 99922 421342 99978
rect 421398 99922 421494 99978
rect 420874 82350 421494 99922
rect 420874 82294 420970 82350
rect 421026 82294 421094 82350
rect 421150 82294 421218 82350
rect 421274 82294 421342 82350
rect 421398 82294 421494 82350
rect 420874 82226 421494 82294
rect 420874 82170 420970 82226
rect 421026 82170 421094 82226
rect 421150 82170 421218 82226
rect 421274 82170 421342 82226
rect 421398 82170 421494 82226
rect 420874 82102 421494 82170
rect 420874 82046 420970 82102
rect 421026 82046 421094 82102
rect 421150 82046 421218 82102
rect 421274 82046 421342 82102
rect 421398 82046 421494 82102
rect 420874 81978 421494 82046
rect 420874 81922 420970 81978
rect 421026 81922 421094 81978
rect 421150 81922 421218 81978
rect 421274 81922 421342 81978
rect 421398 81922 421494 81978
rect 420874 64350 421494 81922
rect 420874 64294 420970 64350
rect 421026 64294 421094 64350
rect 421150 64294 421218 64350
rect 421274 64294 421342 64350
rect 421398 64294 421494 64350
rect 420874 64226 421494 64294
rect 420874 64170 420970 64226
rect 421026 64170 421094 64226
rect 421150 64170 421218 64226
rect 421274 64170 421342 64226
rect 421398 64170 421494 64226
rect 420874 64102 421494 64170
rect 420874 64046 420970 64102
rect 421026 64046 421094 64102
rect 421150 64046 421218 64102
rect 421274 64046 421342 64102
rect 421398 64046 421494 64102
rect 420874 63978 421494 64046
rect 420874 63922 420970 63978
rect 421026 63922 421094 63978
rect 421150 63922 421218 63978
rect 421274 63922 421342 63978
rect 421398 63922 421494 63978
rect 420874 46350 421494 63922
rect 420874 46294 420970 46350
rect 421026 46294 421094 46350
rect 421150 46294 421218 46350
rect 421274 46294 421342 46350
rect 421398 46294 421494 46350
rect 420874 46226 421494 46294
rect 420874 46170 420970 46226
rect 421026 46170 421094 46226
rect 421150 46170 421218 46226
rect 421274 46170 421342 46226
rect 421398 46170 421494 46226
rect 420874 46102 421494 46170
rect 420874 46046 420970 46102
rect 421026 46046 421094 46102
rect 421150 46046 421218 46102
rect 421274 46046 421342 46102
rect 421398 46046 421494 46102
rect 420874 45978 421494 46046
rect 420874 45922 420970 45978
rect 421026 45922 421094 45978
rect 421150 45922 421218 45978
rect 421274 45922 421342 45978
rect 421398 45922 421494 45978
rect 420874 28350 421494 45922
rect 420874 28294 420970 28350
rect 421026 28294 421094 28350
rect 421150 28294 421218 28350
rect 421274 28294 421342 28350
rect 421398 28294 421494 28350
rect 420874 28226 421494 28294
rect 420874 28170 420970 28226
rect 421026 28170 421094 28226
rect 421150 28170 421218 28226
rect 421274 28170 421342 28226
rect 421398 28170 421494 28226
rect 420874 28102 421494 28170
rect 420874 28046 420970 28102
rect 421026 28046 421094 28102
rect 421150 28046 421218 28102
rect 421274 28046 421342 28102
rect 421398 28046 421494 28102
rect 420874 27978 421494 28046
rect 420874 27922 420970 27978
rect 421026 27922 421094 27978
rect 421150 27922 421218 27978
rect 421274 27922 421342 27978
rect 421398 27922 421494 27978
rect 420874 10350 421494 27922
rect 420874 10294 420970 10350
rect 421026 10294 421094 10350
rect 421150 10294 421218 10350
rect 421274 10294 421342 10350
rect 421398 10294 421494 10350
rect 420874 10226 421494 10294
rect 420874 10170 420970 10226
rect 421026 10170 421094 10226
rect 421150 10170 421218 10226
rect 421274 10170 421342 10226
rect 421398 10170 421494 10226
rect 420874 10102 421494 10170
rect 420874 10046 420970 10102
rect 421026 10046 421094 10102
rect 421150 10046 421218 10102
rect 421274 10046 421342 10102
rect 421398 10046 421494 10102
rect 420874 9978 421494 10046
rect 420874 9922 420970 9978
rect 421026 9922 421094 9978
rect 421150 9922 421218 9978
rect 421274 9922 421342 9978
rect 421398 9922 421494 9978
rect 420874 -1120 421494 9922
rect 420874 -1176 420970 -1120
rect 421026 -1176 421094 -1120
rect 421150 -1176 421218 -1120
rect 421274 -1176 421342 -1120
rect 421398 -1176 421494 -1120
rect 420874 -1244 421494 -1176
rect 420874 -1300 420970 -1244
rect 421026 -1300 421094 -1244
rect 421150 -1300 421218 -1244
rect 421274 -1300 421342 -1244
rect 421398 -1300 421494 -1244
rect 420874 -1368 421494 -1300
rect 420874 -1424 420970 -1368
rect 421026 -1424 421094 -1368
rect 421150 -1424 421218 -1368
rect 421274 -1424 421342 -1368
rect 421398 -1424 421494 -1368
rect 420874 -1492 421494 -1424
rect 420874 -1548 420970 -1492
rect 421026 -1548 421094 -1492
rect 421150 -1548 421218 -1492
rect 421274 -1548 421342 -1492
rect 421398 -1548 421494 -1492
rect 420874 -1644 421494 -1548
rect 435154 148350 435774 158858
rect 435154 148294 435250 148350
rect 435306 148294 435374 148350
rect 435430 148294 435498 148350
rect 435554 148294 435622 148350
rect 435678 148294 435774 148350
rect 435154 148226 435774 148294
rect 435154 148170 435250 148226
rect 435306 148170 435374 148226
rect 435430 148170 435498 148226
rect 435554 148170 435622 148226
rect 435678 148170 435774 148226
rect 435154 148102 435774 148170
rect 435154 148046 435250 148102
rect 435306 148046 435374 148102
rect 435430 148046 435498 148102
rect 435554 148046 435622 148102
rect 435678 148046 435774 148102
rect 435154 147978 435774 148046
rect 435154 147922 435250 147978
rect 435306 147922 435374 147978
rect 435430 147922 435498 147978
rect 435554 147922 435622 147978
rect 435678 147922 435774 147978
rect 435154 130350 435774 147922
rect 435154 130294 435250 130350
rect 435306 130294 435374 130350
rect 435430 130294 435498 130350
rect 435554 130294 435622 130350
rect 435678 130294 435774 130350
rect 435154 130226 435774 130294
rect 435154 130170 435250 130226
rect 435306 130170 435374 130226
rect 435430 130170 435498 130226
rect 435554 130170 435622 130226
rect 435678 130170 435774 130226
rect 435154 130102 435774 130170
rect 435154 130046 435250 130102
rect 435306 130046 435374 130102
rect 435430 130046 435498 130102
rect 435554 130046 435622 130102
rect 435678 130046 435774 130102
rect 435154 129978 435774 130046
rect 435154 129922 435250 129978
rect 435306 129922 435374 129978
rect 435430 129922 435498 129978
rect 435554 129922 435622 129978
rect 435678 129922 435774 129978
rect 435154 112350 435774 129922
rect 435154 112294 435250 112350
rect 435306 112294 435374 112350
rect 435430 112294 435498 112350
rect 435554 112294 435622 112350
rect 435678 112294 435774 112350
rect 435154 112226 435774 112294
rect 435154 112170 435250 112226
rect 435306 112170 435374 112226
rect 435430 112170 435498 112226
rect 435554 112170 435622 112226
rect 435678 112170 435774 112226
rect 435154 112102 435774 112170
rect 435154 112046 435250 112102
rect 435306 112046 435374 112102
rect 435430 112046 435498 112102
rect 435554 112046 435622 112102
rect 435678 112046 435774 112102
rect 435154 111978 435774 112046
rect 435154 111922 435250 111978
rect 435306 111922 435374 111978
rect 435430 111922 435498 111978
rect 435554 111922 435622 111978
rect 435678 111922 435774 111978
rect 435154 94350 435774 111922
rect 435154 94294 435250 94350
rect 435306 94294 435374 94350
rect 435430 94294 435498 94350
rect 435554 94294 435622 94350
rect 435678 94294 435774 94350
rect 435154 94226 435774 94294
rect 435154 94170 435250 94226
rect 435306 94170 435374 94226
rect 435430 94170 435498 94226
rect 435554 94170 435622 94226
rect 435678 94170 435774 94226
rect 435154 94102 435774 94170
rect 435154 94046 435250 94102
rect 435306 94046 435374 94102
rect 435430 94046 435498 94102
rect 435554 94046 435622 94102
rect 435678 94046 435774 94102
rect 435154 93978 435774 94046
rect 435154 93922 435250 93978
rect 435306 93922 435374 93978
rect 435430 93922 435498 93978
rect 435554 93922 435622 93978
rect 435678 93922 435774 93978
rect 435154 76350 435774 93922
rect 435154 76294 435250 76350
rect 435306 76294 435374 76350
rect 435430 76294 435498 76350
rect 435554 76294 435622 76350
rect 435678 76294 435774 76350
rect 435154 76226 435774 76294
rect 435154 76170 435250 76226
rect 435306 76170 435374 76226
rect 435430 76170 435498 76226
rect 435554 76170 435622 76226
rect 435678 76170 435774 76226
rect 435154 76102 435774 76170
rect 435154 76046 435250 76102
rect 435306 76046 435374 76102
rect 435430 76046 435498 76102
rect 435554 76046 435622 76102
rect 435678 76046 435774 76102
rect 435154 75978 435774 76046
rect 435154 75922 435250 75978
rect 435306 75922 435374 75978
rect 435430 75922 435498 75978
rect 435554 75922 435622 75978
rect 435678 75922 435774 75978
rect 435154 58350 435774 75922
rect 435154 58294 435250 58350
rect 435306 58294 435374 58350
rect 435430 58294 435498 58350
rect 435554 58294 435622 58350
rect 435678 58294 435774 58350
rect 435154 58226 435774 58294
rect 435154 58170 435250 58226
rect 435306 58170 435374 58226
rect 435430 58170 435498 58226
rect 435554 58170 435622 58226
rect 435678 58170 435774 58226
rect 435154 58102 435774 58170
rect 435154 58046 435250 58102
rect 435306 58046 435374 58102
rect 435430 58046 435498 58102
rect 435554 58046 435622 58102
rect 435678 58046 435774 58102
rect 435154 57978 435774 58046
rect 435154 57922 435250 57978
rect 435306 57922 435374 57978
rect 435430 57922 435498 57978
rect 435554 57922 435622 57978
rect 435678 57922 435774 57978
rect 435154 40350 435774 57922
rect 435154 40294 435250 40350
rect 435306 40294 435374 40350
rect 435430 40294 435498 40350
rect 435554 40294 435622 40350
rect 435678 40294 435774 40350
rect 435154 40226 435774 40294
rect 435154 40170 435250 40226
rect 435306 40170 435374 40226
rect 435430 40170 435498 40226
rect 435554 40170 435622 40226
rect 435678 40170 435774 40226
rect 435154 40102 435774 40170
rect 435154 40046 435250 40102
rect 435306 40046 435374 40102
rect 435430 40046 435498 40102
rect 435554 40046 435622 40102
rect 435678 40046 435774 40102
rect 435154 39978 435774 40046
rect 435154 39922 435250 39978
rect 435306 39922 435374 39978
rect 435430 39922 435498 39978
rect 435554 39922 435622 39978
rect 435678 39922 435774 39978
rect 435154 22350 435774 39922
rect 435154 22294 435250 22350
rect 435306 22294 435374 22350
rect 435430 22294 435498 22350
rect 435554 22294 435622 22350
rect 435678 22294 435774 22350
rect 435154 22226 435774 22294
rect 435154 22170 435250 22226
rect 435306 22170 435374 22226
rect 435430 22170 435498 22226
rect 435554 22170 435622 22226
rect 435678 22170 435774 22226
rect 435154 22102 435774 22170
rect 435154 22046 435250 22102
rect 435306 22046 435374 22102
rect 435430 22046 435498 22102
rect 435554 22046 435622 22102
rect 435678 22046 435774 22102
rect 435154 21978 435774 22046
rect 435154 21922 435250 21978
rect 435306 21922 435374 21978
rect 435430 21922 435498 21978
rect 435554 21922 435622 21978
rect 435678 21922 435774 21978
rect 435154 4350 435774 21922
rect 435154 4294 435250 4350
rect 435306 4294 435374 4350
rect 435430 4294 435498 4350
rect 435554 4294 435622 4350
rect 435678 4294 435774 4350
rect 435154 4226 435774 4294
rect 435154 4170 435250 4226
rect 435306 4170 435374 4226
rect 435430 4170 435498 4226
rect 435554 4170 435622 4226
rect 435678 4170 435774 4226
rect 435154 4102 435774 4170
rect 435154 4046 435250 4102
rect 435306 4046 435374 4102
rect 435430 4046 435498 4102
rect 435554 4046 435622 4102
rect 435678 4046 435774 4102
rect 435154 3978 435774 4046
rect 435154 3922 435250 3978
rect 435306 3922 435374 3978
rect 435430 3922 435498 3978
rect 435554 3922 435622 3978
rect 435678 3922 435774 3978
rect 435154 -160 435774 3922
rect 435154 -216 435250 -160
rect 435306 -216 435374 -160
rect 435430 -216 435498 -160
rect 435554 -216 435622 -160
rect 435678 -216 435774 -160
rect 435154 -284 435774 -216
rect 435154 -340 435250 -284
rect 435306 -340 435374 -284
rect 435430 -340 435498 -284
rect 435554 -340 435622 -284
rect 435678 -340 435774 -284
rect 435154 -408 435774 -340
rect 435154 -464 435250 -408
rect 435306 -464 435374 -408
rect 435430 -464 435498 -408
rect 435554 -464 435622 -408
rect 435678 -464 435774 -408
rect 435154 -532 435774 -464
rect 435154 -588 435250 -532
rect 435306 -588 435374 -532
rect 435430 -588 435498 -532
rect 435554 -588 435622 -532
rect 435678 -588 435774 -532
rect 435154 -1644 435774 -588
rect 438874 154350 439494 158858
rect 438874 154294 438970 154350
rect 439026 154294 439094 154350
rect 439150 154294 439218 154350
rect 439274 154294 439342 154350
rect 439398 154294 439494 154350
rect 438874 154226 439494 154294
rect 438874 154170 438970 154226
rect 439026 154170 439094 154226
rect 439150 154170 439218 154226
rect 439274 154170 439342 154226
rect 439398 154170 439494 154226
rect 438874 154102 439494 154170
rect 438874 154046 438970 154102
rect 439026 154046 439094 154102
rect 439150 154046 439218 154102
rect 439274 154046 439342 154102
rect 439398 154046 439494 154102
rect 438874 153978 439494 154046
rect 438874 153922 438970 153978
rect 439026 153922 439094 153978
rect 439150 153922 439218 153978
rect 439274 153922 439342 153978
rect 439398 153922 439494 153978
rect 438874 136350 439494 153922
rect 438874 136294 438970 136350
rect 439026 136294 439094 136350
rect 439150 136294 439218 136350
rect 439274 136294 439342 136350
rect 439398 136294 439494 136350
rect 438874 136226 439494 136294
rect 438874 136170 438970 136226
rect 439026 136170 439094 136226
rect 439150 136170 439218 136226
rect 439274 136170 439342 136226
rect 439398 136170 439494 136226
rect 438874 136102 439494 136170
rect 438874 136046 438970 136102
rect 439026 136046 439094 136102
rect 439150 136046 439218 136102
rect 439274 136046 439342 136102
rect 439398 136046 439494 136102
rect 438874 135978 439494 136046
rect 438874 135922 438970 135978
rect 439026 135922 439094 135978
rect 439150 135922 439218 135978
rect 439274 135922 439342 135978
rect 439398 135922 439494 135978
rect 438874 118350 439494 135922
rect 438874 118294 438970 118350
rect 439026 118294 439094 118350
rect 439150 118294 439218 118350
rect 439274 118294 439342 118350
rect 439398 118294 439494 118350
rect 438874 118226 439494 118294
rect 438874 118170 438970 118226
rect 439026 118170 439094 118226
rect 439150 118170 439218 118226
rect 439274 118170 439342 118226
rect 439398 118170 439494 118226
rect 438874 118102 439494 118170
rect 438874 118046 438970 118102
rect 439026 118046 439094 118102
rect 439150 118046 439218 118102
rect 439274 118046 439342 118102
rect 439398 118046 439494 118102
rect 438874 117978 439494 118046
rect 438874 117922 438970 117978
rect 439026 117922 439094 117978
rect 439150 117922 439218 117978
rect 439274 117922 439342 117978
rect 439398 117922 439494 117978
rect 438874 100350 439494 117922
rect 438874 100294 438970 100350
rect 439026 100294 439094 100350
rect 439150 100294 439218 100350
rect 439274 100294 439342 100350
rect 439398 100294 439494 100350
rect 438874 100226 439494 100294
rect 438874 100170 438970 100226
rect 439026 100170 439094 100226
rect 439150 100170 439218 100226
rect 439274 100170 439342 100226
rect 439398 100170 439494 100226
rect 438874 100102 439494 100170
rect 438874 100046 438970 100102
rect 439026 100046 439094 100102
rect 439150 100046 439218 100102
rect 439274 100046 439342 100102
rect 439398 100046 439494 100102
rect 438874 99978 439494 100046
rect 438874 99922 438970 99978
rect 439026 99922 439094 99978
rect 439150 99922 439218 99978
rect 439274 99922 439342 99978
rect 439398 99922 439494 99978
rect 438874 82350 439494 99922
rect 438874 82294 438970 82350
rect 439026 82294 439094 82350
rect 439150 82294 439218 82350
rect 439274 82294 439342 82350
rect 439398 82294 439494 82350
rect 438874 82226 439494 82294
rect 438874 82170 438970 82226
rect 439026 82170 439094 82226
rect 439150 82170 439218 82226
rect 439274 82170 439342 82226
rect 439398 82170 439494 82226
rect 438874 82102 439494 82170
rect 438874 82046 438970 82102
rect 439026 82046 439094 82102
rect 439150 82046 439218 82102
rect 439274 82046 439342 82102
rect 439398 82046 439494 82102
rect 438874 81978 439494 82046
rect 438874 81922 438970 81978
rect 439026 81922 439094 81978
rect 439150 81922 439218 81978
rect 439274 81922 439342 81978
rect 439398 81922 439494 81978
rect 438874 64350 439494 81922
rect 438874 64294 438970 64350
rect 439026 64294 439094 64350
rect 439150 64294 439218 64350
rect 439274 64294 439342 64350
rect 439398 64294 439494 64350
rect 438874 64226 439494 64294
rect 438874 64170 438970 64226
rect 439026 64170 439094 64226
rect 439150 64170 439218 64226
rect 439274 64170 439342 64226
rect 439398 64170 439494 64226
rect 438874 64102 439494 64170
rect 438874 64046 438970 64102
rect 439026 64046 439094 64102
rect 439150 64046 439218 64102
rect 439274 64046 439342 64102
rect 439398 64046 439494 64102
rect 438874 63978 439494 64046
rect 438874 63922 438970 63978
rect 439026 63922 439094 63978
rect 439150 63922 439218 63978
rect 439274 63922 439342 63978
rect 439398 63922 439494 63978
rect 438874 46350 439494 63922
rect 438874 46294 438970 46350
rect 439026 46294 439094 46350
rect 439150 46294 439218 46350
rect 439274 46294 439342 46350
rect 439398 46294 439494 46350
rect 438874 46226 439494 46294
rect 438874 46170 438970 46226
rect 439026 46170 439094 46226
rect 439150 46170 439218 46226
rect 439274 46170 439342 46226
rect 439398 46170 439494 46226
rect 438874 46102 439494 46170
rect 438874 46046 438970 46102
rect 439026 46046 439094 46102
rect 439150 46046 439218 46102
rect 439274 46046 439342 46102
rect 439398 46046 439494 46102
rect 438874 45978 439494 46046
rect 438874 45922 438970 45978
rect 439026 45922 439094 45978
rect 439150 45922 439218 45978
rect 439274 45922 439342 45978
rect 439398 45922 439494 45978
rect 438874 28350 439494 45922
rect 438874 28294 438970 28350
rect 439026 28294 439094 28350
rect 439150 28294 439218 28350
rect 439274 28294 439342 28350
rect 439398 28294 439494 28350
rect 438874 28226 439494 28294
rect 438874 28170 438970 28226
rect 439026 28170 439094 28226
rect 439150 28170 439218 28226
rect 439274 28170 439342 28226
rect 439398 28170 439494 28226
rect 438874 28102 439494 28170
rect 438874 28046 438970 28102
rect 439026 28046 439094 28102
rect 439150 28046 439218 28102
rect 439274 28046 439342 28102
rect 439398 28046 439494 28102
rect 438874 27978 439494 28046
rect 438874 27922 438970 27978
rect 439026 27922 439094 27978
rect 439150 27922 439218 27978
rect 439274 27922 439342 27978
rect 439398 27922 439494 27978
rect 438874 10350 439494 27922
rect 438874 10294 438970 10350
rect 439026 10294 439094 10350
rect 439150 10294 439218 10350
rect 439274 10294 439342 10350
rect 439398 10294 439494 10350
rect 438874 10226 439494 10294
rect 438874 10170 438970 10226
rect 439026 10170 439094 10226
rect 439150 10170 439218 10226
rect 439274 10170 439342 10226
rect 439398 10170 439494 10226
rect 438874 10102 439494 10170
rect 438874 10046 438970 10102
rect 439026 10046 439094 10102
rect 439150 10046 439218 10102
rect 439274 10046 439342 10102
rect 439398 10046 439494 10102
rect 438874 9978 439494 10046
rect 438874 9922 438970 9978
rect 439026 9922 439094 9978
rect 439150 9922 439218 9978
rect 439274 9922 439342 9978
rect 439398 9922 439494 9978
rect 438874 -1120 439494 9922
rect 438874 -1176 438970 -1120
rect 439026 -1176 439094 -1120
rect 439150 -1176 439218 -1120
rect 439274 -1176 439342 -1120
rect 439398 -1176 439494 -1120
rect 438874 -1244 439494 -1176
rect 438874 -1300 438970 -1244
rect 439026 -1300 439094 -1244
rect 439150 -1300 439218 -1244
rect 439274 -1300 439342 -1244
rect 439398 -1300 439494 -1244
rect 438874 -1368 439494 -1300
rect 438874 -1424 438970 -1368
rect 439026 -1424 439094 -1368
rect 439150 -1424 439218 -1368
rect 439274 -1424 439342 -1368
rect 439398 -1424 439494 -1368
rect 438874 -1492 439494 -1424
rect 438874 -1548 438970 -1492
rect 439026 -1548 439094 -1492
rect 439150 -1548 439218 -1492
rect 439274 -1548 439342 -1492
rect 439398 -1548 439494 -1492
rect 438874 -1644 439494 -1548
rect 453154 148350 453774 158858
rect 453154 148294 453250 148350
rect 453306 148294 453374 148350
rect 453430 148294 453498 148350
rect 453554 148294 453622 148350
rect 453678 148294 453774 148350
rect 453154 148226 453774 148294
rect 453154 148170 453250 148226
rect 453306 148170 453374 148226
rect 453430 148170 453498 148226
rect 453554 148170 453622 148226
rect 453678 148170 453774 148226
rect 453154 148102 453774 148170
rect 453154 148046 453250 148102
rect 453306 148046 453374 148102
rect 453430 148046 453498 148102
rect 453554 148046 453622 148102
rect 453678 148046 453774 148102
rect 453154 147978 453774 148046
rect 453154 147922 453250 147978
rect 453306 147922 453374 147978
rect 453430 147922 453498 147978
rect 453554 147922 453622 147978
rect 453678 147922 453774 147978
rect 453154 130350 453774 147922
rect 453154 130294 453250 130350
rect 453306 130294 453374 130350
rect 453430 130294 453498 130350
rect 453554 130294 453622 130350
rect 453678 130294 453774 130350
rect 453154 130226 453774 130294
rect 453154 130170 453250 130226
rect 453306 130170 453374 130226
rect 453430 130170 453498 130226
rect 453554 130170 453622 130226
rect 453678 130170 453774 130226
rect 453154 130102 453774 130170
rect 453154 130046 453250 130102
rect 453306 130046 453374 130102
rect 453430 130046 453498 130102
rect 453554 130046 453622 130102
rect 453678 130046 453774 130102
rect 453154 129978 453774 130046
rect 453154 129922 453250 129978
rect 453306 129922 453374 129978
rect 453430 129922 453498 129978
rect 453554 129922 453622 129978
rect 453678 129922 453774 129978
rect 453154 112350 453774 129922
rect 453154 112294 453250 112350
rect 453306 112294 453374 112350
rect 453430 112294 453498 112350
rect 453554 112294 453622 112350
rect 453678 112294 453774 112350
rect 453154 112226 453774 112294
rect 453154 112170 453250 112226
rect 453306 112170 453374 112226
rect 453430 112170 453498 112226
rect 453554 112170 453622 112226
rect 453678 112170 453774 112226
rect 453154 112102 453774 112170
rect 453154 112046 453250 112102
rect 453306 112046 453374 112102
rect 453430 112046 453498 112102
rect 453554 112046 453622 112102
rect 453678 112046 453774 112102
rect 453154 111978 453774 112046
rect 453154 111922 453250 111978
rect 453306 111922 453374 111978
rect 453430 111922 453498 111978
rect 453554 111922 453622 111978
rect 453678 111922 453774 111978
rect 453154 94350 453774 111922
rect 453154 94294 453250 94350
rect 453306 94294 453374 94350
rect 453430 94294 453498 94350
rect 453554 94294 453622 94350
rect 453678 94294 453774 94350
rect 453154 94226 453774 94294
rect 453154 94170 453250 94226
rect 453306 94170 453374 94226
rect 453430 94170 453498 94226
rect 453554 94170 453622 94226
rect 453678 94170 453774 94226
rect 453154 94102 453774 94170
rect 453154 94046 453250 94102
rect 453306 94046 453374 94102
rect 453430 94046 453498 94102
rect 453554 94046 453622 94102
rect 453678 94046 453774 94102
rect 453154 93978 453774 94046
rect 453154 93922 453250 93978
rect 453306 93922 453374 93978
rect 453430 93922 453498 93978
rect 453554 93922 453622 93978
rect 453678 93922 453774 93978
rect 453154 76350 453774 93922
rect 453154 76294 453250 76350
rect 453306 76294 453374 76350
rect 453430 76294 453498 76350
rect 453554 76294 453622 76350
rect 453678 76294 453774 76350
rect 453154 76226 453774 76294
rect 453154 76170 453250 76226
rect 453306 76170 453374 76226
rect 453430 76170 453498 76226
rect 453554 76170 453622 76226
rect 453678 76170 453774 76226
rect 453154 76102 453774 76170
rect 453154 76046 453250 76102
rect 453306 76046 453374 76102
rect 453430 76046 453498 76102
rect 453554 76046 453622 76102
rect 453678 76046 453774 76102
rect 453154 75978 453774 76046
rect 453154 75922 453250 75978
rect 453306 75922 453374 75978
rect 453430 75922 453498 75978
rect 453554 75922 453622 75978
rect 453678 75922 453774 75978
rect 453154 58350 453774 75922
rect 453154 58294 453250 58350
rect 453306 58294 453374 58350
rect 453430 58294 453498 58350
rect 453554 58294 453622 58350
rect 453678 58294 453774 58350
rect 453154 58226 453774 58294
rect 453154 58170 453250 58226
rect 453306 58170 453374 58226
rect 453430 58170 453498 58226
rect 453554 58170 453622 58226
rect 453678 58170 453774 58226
rect 453154 58102 453774 58170
rect 453154 58046 453250 58102
rect 453306 58046 453374 58102
rect 453430 58046 453498 58102
rect 453554 58046 453622 58102
rect 453678 58046 453774 58102
rect 453154 57978 453774 58046
rect 453154 57922 453250 57978
rect 453306 57922 453374 57978
rect 453430 57922 453498 57978
rect 453554 57922 453622 57978
rect 453678 57922 453774 57978
rect 453154 40350 453774 57922
rect 453154 40294 453250 40350
rect 453306 40294 453374 40350
rect 453430 40294 453498 40350
rect 453554 40294 453622 40350
rect 453678 40294 453774 40350
rect 453154 40226 453774 40294
rect 453154 40170 453250 40226
rect 453306 40170 453374 40226
rect 453430 40170 453498 40226
rect 453554 40170 453622 40226
rect 453678 40170 453774 40226
rect 453154 40102 453774 40170
rect 453154 40046 453250 40102
rect 453306 40046 453374 40102
rect 453430 40046 453498 40102
rect 453554 40046 453622 40102
rect 453678 40046 453774 40102
rect 453154 39978 453774 40046
rect 453154 39922 453250 39978
rect 453306 39922 453374 39978
rect 453430 39922 453498 39978
rect 453554 39922 453622 39978
rect 453678 39922 453774 39978
rect 453154 22350 453774 39922
rect 453154 22294 453250 22350
rect 453306 22294 453374 22350
rect 453430 22294 453498 22350
rect 453554 22294 453622 22350
rect 453678 22294 453774 22350
rect 453154 22226 453774 22294
rect 453154 22170 453250 22226
rect 453306 22170 453374 22226
rect 453430 22170 453498 22226
rect 453554 22170 453622 22226
rect 453678 22170 453774 22226
rect 453154 22102 453774 22170
rect 453154 22046 453250 22102
rect 453306 22046 453374 22102
rect 453430 22046 453498 22102
rect 453554 22046 453622 22102
rect 453678 22046 453774 22102
rect 453154 21978 453774 22046
rect 453154 21922 453250 21978
rect 453306 21922 453374 21978
rect 453430 21922 453498 21978
rect 453554 21922 453622 21978
rect 453678 21922 453774 21978
rect 453154 4350 453774 21922
rect 453154 4294 453250 4350
rect 453306 4294 453374 4350
rect 453430 4294 453498 4350
rect 453554 4294 453622 4350
rect 453678 4294 453774 4350
rect 453154 4226 453774 4294
rect 453154 4170 453250 4226
rect 453306 4170 453374 4226
rect 453430 4170 453498 4226
rect 453554 4170 453622 4226
rect 453678 4170 453774 4226
rect 453154 4102 453774 4170
rect 453154 4046 453250 4102
rect 453306 4046 453374 4102
rect 453430 4046 453498 4102
rect 453554 4046 453622 4102
rect 453678 4046 453774 4102
rect 453154 3978 453774 4046
rect 453154 3922 453250 3978
rect 453306 3922 453374 3978
rect 453430 3922 453498 3978
rect 453554 3922 453622 3978
rect 453678 3922 453774 3978
rect 453154 -160 453774 3922
rect 453154 -216 453250 -160
rect 453306 -216 453374 -160
rect 453430 -216 453498 -160
rect 453554 -216 453622 -160
rect 453678 -216 453774 -160
rect 453154 -284 453774 -216
rect 453154 -340 453250 -284
rect 453306 -340 453374 -284
rect 453430 -340 453498 -284
rect 453554 -340 453622 -284
rect 453678 -340 453774 -284
rect 453154 -408 453774 -340
rect 453154 -464 453250 -408
rect 453306 -464 453374 -408
rect 453430 -464 453498 -408
rect 453554 -464 453622 -408
rect 453678 -464 453774 -408
rect 453154 -532 453774 -464
rect 453154 -588 453250 -532
rect 453306 -588 453374 -532
rect 453430 -588 453498 -532
rect 453554 -588 453622 -532
rect 453678 -588 453774 -532
rect 453154 -1644 453774 -588
rect 456874 154350 457494 158858
rect 456874 154294 456970 154350
rect 457026 154294 457094 154350
rect 457150 154294 457218 154350
rect 457274 154294 457342 154350
rect 457398 154294 457494 154350
rect 456874 154226 457494 154294
rect 456874 154170 456970 154226
rect 457026 154170 457094 154226
rect 457150 154170 457218 154226
rect 457274 154170 457342 154226
rect 457398 154170 457494 154226
rect 456874 154102 457494 154170
rect 456874 154046 456970 154102
rect 457026 154046 457094 154102
rect 457150 154046 457218 154102
rect 457274 154046 457342 154102
rect 457398 154046 457494 154102
rect 456874 153978 457494 154046
rect 456874 153922 456970 153978
rect 457026 153922 457094 153978
rect 457150 153922 457218 153978
rect 457274 153922 457342 153978
rect 457398 153922 457494 153978
rect 456874 136350 457494 153922
rect 456874 136294 456970 136350
rect 457026 136294 457094 136350
rect 457150 136294 457218 136350
rect 457274 136294 457342 136350
rect 457398 136294 457494 136350
rect 456874 136226 457494 136294
rect 456874 136170 456970 136226
rect 457026 136170 457094 136226
rect 457150 136170 457218 136226
rect 457274 136170 457342 136226
rect 457398 136170 457494 136226
rect 456874 136102 457494 136170
rect 456874 136046 456970 136102
rect 457026 136046 457094 136102
rect 457150 136046 457218 136102
rect 457274 136046 457342 136102
rect 457398 136046 457494 136102
rect 456874 135978 457494 136046
rect 456874 135922 456970 135978
rect 457026 135922 457094 135978
rect 457150 135922 457218 135978
rect 457274 135922 457342 135978
rect 457398 135922 457494 135978
rect 456874 118350 457494 135922
rect 456874 118294 456970 118350
rect 457026 118294 457094 118350
rect 457150 118294 457218 118350
rect 457274 118294 457342 118350
rect 457398 118294 457494 118350
rect 456874 118226 457494 118294
rect 456874 118170 456970 118226
rect 457026 118170 457094 118226
rect 457150 118170 457218 118226
rect 457274 118170 457342 118226
rect 457398 118170 457494 118226
rect 456874 118102 457494 118170
rect 456874 118046 456970 118102
rect 457026 118046 457094 118102
rect 457150 118046 457218 118102
rect 457274 118046 457342 118102
rect 457398 118046 457494 118102
rect 456874 117978 457494 118046
rect 456874 117922 456970 117978
rect 457026 117922 457094 117978
rect 457150 117922 457218 117978
rect 457274 117922 457342 117978
rect 457398 117922 457494 117978
rect 456874 100350 457494 117922
rect 456874 100294 456970 100350
rect 457026 100294 457094 100350
rect 457150 100294 457218 100350
rect 457274 100294 457342 100350
rect 457398 100294 457494 100350
rect 456874 100226 457494 100294
rect 456874 100170 456970 100226
rect 457026 100170 457094 100226
rect 457150 100170 457218 100226
rect 457274 100170 457342 100226
rect 457398 100170 457494 100226
rect 456874 100102 457494 100170
rect 456874 100046 456970 100102
rect 457026 100046 457094 100102
rect 457150 100046 457218 100102
rect 457274 100046 457342 100102
rect 457398 100046 457494 100102
rect 456874 99978 457494 100046
rect 456874 99922 456970 99978
rect 457026 99922 457094 99978
rect 457150 99922 457218 99978
rect 457274 99922 457342 99978
rect 457398 99922 457494 99978
rect 456874 82350 457494 99922
rect 456874 82294 456970 82350
rect 457026 82294 457094 82350
rect 457150 82294 457218 82350
rect 457274 82294 457342 82350
rect 457398 82294 457494 82350
rect 456874 82226 457494 82294
rect 456874 82170 456970 82226
rect 457026 82170 457094 82226
rect 457150 82170 457218 82226
rect 457274 82170 457342 82226
rect 457398 82170 457494 82226
rect 456874 82102 457494 82170
rect 456874 82046 456970 82102
rect 457026 82046 457094 82102
rect 457150 82046 457218 82102
rect 457274 82046 457342 82102
rect 457398 82046 457494 82102
rect 456874 81978 457494 82046
rect 456874 81922 456970 81978
rect 457026 81922 457094 81978
rect 457150 81922 457218 81978
rect 457274 81922 457342 81978
rect 457398 81922 457494 81978
rect 456874 64350 457494 81922
rect 456874 64294 456970 64350
rect 457026 64294 457094 64350
rect 457150 64294 457218 64350
rect 457274 64294 457342 64350
rect 457398 64294 457494 64350
rect 456874 64226 457494 64294
rect 456874 64170 456970 64226
rect 457026 64170 457094 64226
rect 457150 64170 457218 64226
rect 457274 64170 457342 64226
rect 457398 64170 457494 64226
rect 456874 64102 457494 64170
rect 456874 64046 456970 64102
rect 457026 64046 457094 64102
rect 457150 64046 457218 64102
rect 457274 64046 457342 64102
rect 457398 64046 457494 64102
rect 456874 63978 457494 64046
rect 456874 63922 456970 63978
rect 457026 63922 457094 63978
rect 457150 63922 457218 63978
rect 457274 63922 457342 63978
rect 457398 63922 457494 63978
rect 456874 46350 457494 63922
rect 456874 46294 456970 46350
rect 457026 46294 457094 46350
rect 457150 46294 457218 46350
rect 457274 46294 457342 46350
rect 457398 46294 457494 46350
rect 456874 46226 457494 46294
rect 456874 46170 456970 46226
rect 457026 46170 457094 46226
rect 457150 46170 457218 46226
rect 457274 46170 457342 46226
rect 457398 46170 457494 46226
rect 456874 46102 457494 46170
rect 456874 46046 456970 46102
rect 457026 46046 457094 46102
rect 457150 46046 457218 46102
rect 457274 46046 457342 46102
rect 457398 46046 457494 46102
rect 456874 45978 457494 46046
rect 456874 45922 456970 45978
rect 457026 45922 457094 45978
rect 457150 45922 457218 45978
rect 457274 45922 457342 45978
rect 457398 45922 457494 45978
rect 456874 28350 457494 45922
rect 456874 28294 456970 28350
rect 457026 28294 457094 28350
rect 457150 28294 457218 28350
rect 457274 28294 457342 28350
rect 457398 28294 457494 28350
rect 456874 28226 457494 28294
rect 456874 28170 456970 28226
rect 457026 28170 457094 28226
rect 457150 28170 457218 28226
rect 457274 28170 457342 28226
rect 457398 28170 457494 28226
rect 456874 28102 457494 28170
rect 456874 28046 456970 28102
rect 457026 28046 457094 28102
rect 457150 28046 457218 28102
rect 457274 28046 457342 28102
rect 457398 28046 457494 28102
rect 456874 27978 457494 28046
rect 456874 27922 456970 27978
rect 457026 27922 457094 27978
rect 457150 27922 457218 27978
rect 457274 27922 457342 27978
rect 457398 27922 457494 27978
rect 456874 10350 457494 27922
rect 456874 10294 456970 10350
rect 457026 10294 457094 10350
rect 457150 10294 457218 10350
rect 457274 10294 457342 10350
rect 457398 10294 457494 10350
rect 456874 10226 457494 10294
rect 456874 10170 456970 10226
rect 457026 10170 457094 10226
rect 457150 10170 457218 10226
rect 457274 10170 457342 10226
rect 457398 10170 457494 10226
rect 456874 10102 457494 10170
rect 456874 10046 456970 10102
rect 457026 10046 457094 10102
rect 457150 10046 457218 10102
rect 457274 10046 457342 10102
rect 457398 10046 457494 10102
rect 456874 9978 457494 10046
rect 456874 9922 456970 9978
rect 457026 9922 457094 9978
rect 457150 9922 457218 9978
rect 457274 9922 457342 9978
rect 457398 9922 457494 9978
rect 456874 -1120 457494 9922
rect 456874 -1176 456970 -1120
rect 457026 -1176 457094 -1120
rect 457150 -1176 457218 -1120
rect 457274 -1176 457342 -1120
rect 457398 -1176 457494 -1120
rect 456874 -1244 457494 -1176
rect 456874 -1300 456970 -1244
rect 457026 -1300 457094 -1244
rect 457150 -1300 457218 -1244
rect 457274 -1300 457342 -1244
rect 457398 -1300 457494 -1244
rect 456874 -1368 457494 -1300
rect 456874 -1424 456970 -1368
rect 457026 -1424 457094 -1368
rect 457150 -1424 457218 -1368
rect 457274 -1424 457342 -1368
rect 457398 -1424 457494 -1368
rect 456874 -1492 457494 -1424
rect 456874 -1548 456970 -1492
rect 457026 -1548 457094 -1492
rect 457150 -1548 457218 -1492
rect 457274 -1548 457342 -1492
rect 457398 -1548 457494 -1492
rect 456874 -1644 457494 -1548
rect 471154 148350 471774 158858
rect 471154 148294 471250 148350
rect 471306 148294 471374 148350
rect 471430 148294 471498 148350
rect 471554 148294 471622 148350
rect 471678 148294 471774 148350
rect 471154 148226 471774 148294
rect 471154 148170 471250 148226
rect 471306 148170 471374 148226
rect 471430 148170 471498 148226
rect 471554 148170 471622 148226
rect 471678 148170 471774 148226
rect 471154 148102 471774 148170
rect 471154 148046 471250 148102
rect 471306 148046 471374 148102
rect 471430 148046 471498 148102
rect 471554 148046 471622 148102
rect 471678 148046 471774 148102
rect 471154 147978 471774 148046
rect 471154 147922 471250 147978
rect 471306 147922 471374 147978
rect 471430 147922 471498 147978
rect 471554 147922 471622 147978
rect 471678 147922 471774 147978
rect 471154 130350 471774 147922
rect 471154 130294 471250 130350
rect 471306 130294 471374 130350
rect 471430 130294 471498 130350
rect 471554 130294 471622 130350
rect 471678 130294 471774 130350
rect 471154 130226 471774 130294
rect 471154 130170 471250 130226
rect 471306 130170 471374 130226
rect 471430 130170 471498 130226
rect 471554 130170 471622 130226
rect 471678 130170 471774 130226
rect 471154 130102 471774 130170
rect 471154 130046 471250 130102
rect 471306 130046 471374 130102
rect 471430 130046 471498 130102
rect 471554 130046 471622 130102
rect 471678 130046 471774 130102
rect 471154 129978 471774 130046
rect 471154 129922 471250 129978
rect 471306 129922 471374 129978
rect 471430 129922 471498 129978
rect 471554 129922 471622 129978
rect 471678 129922 471774 129978
rect 471154 112350 471774 129922
rect 471154 112294 471250 112350
rect 471306 112294 471374 112350
rect 471430 112294 471498 112350
rect 471554 112294 471622 112350
rect 471678 112294 471774 112350
rect 471154 112226 471774 112294
rect 471154 112170 471250 112226
rect 471306 112170 471374 112226
rect 471430 112170 471498 112226
rect 471554 112170 471622 112226
rect 471678 112170 471774 112226
rect 471154 112102 471774 112170
rect 471154 112046 471250 112102
rect 471306 112046 471374 112102
rect 471430 112046 471498 112102
rect 471554 112046 471622 112102
rect 471678 112046 471774 112102
rect 471154 111978 471774 112046
rect 471154 111922 471250 111978
rect 471306 111922 471374 111978
rect 471430 111922 471498 111978
rect 471554 111922 471622 111978
rect 471678 111922 471774 111978
rect 471154 94350 471774 111922
rect 471154 94294 471250 94350
rect 471306 94294 471374 94350
rect 471430 94294 471498 94350
rect 471554 94294 471622 94350
rect 471678 94294 471774 94350
rect 471154 94226 471774 94294
rect 471154 94170 471250 94226
rect 471306 94170 471374 94226
rect 471430 94170 471498 94226
rect 471554 94170 471622 94226
rect 471678 94170 471774 94226
rect 471154 94102 471774 94170
rect 471154 94046 471250 94102
rect 471306 94046 471374 94102
rect 471430 94046 471498 94102
rect 471554 94046 471622 94102
rect 471678 94046 471774 94102
rect 471154 93978 471774 94046
rect 471154 93922 471250 93978
rect 471306 93922 471374 93978
rect 471430 93922 471498 93978
rect 471554 93922 471622 93978
rect 471678 93922 471774 93978
rect 471154 76350 471774 93922
rect 471154 76294 471250 76350
rect 471306 76294 471374 76350
rect 471430 76294 471498 76350
rect 471554 76294 471622 76350
rect 471678 76294 471774 76350
rect 471154 76226 471774 76294
rect 471154 76170 471250 76226
rect 471306 76170 471374 76226
rect 471430 76170 471498 76226
rect 471554 76170 471622 76226
rect 471678 76170 471774 76226
rect 471154 76102 471774 76170
rect 471154 76046 471250 76102
rect 471306 76046 471374 76102
rect 471430 76046 471498 76102
rect 471554 76046 471622 76102
rect 471678 76046 471774 76102
rect 471154 75978 471774 76046
rect 471154 75922 471250 75978
rect 471306 75922 471374 75978
rect 471430 75922 471498 75978
rect 471554 75922 471622 75978
rect 471678 75922 471774 75978
rect 471154 58350 471774 75922
rect 471154 58294 471250 58350
rect 471306 58294 471374 58350
rect 471430 58294 471498 58350
rect 471554 58294 471622 58350
rect 471678 58294 471774 58350
rect 471154 58226 471774 58294
rect 471154 58170 471250 58226
rect 471306 58170 471374 58226
rect 471430 58170 471498 58226
rect 471554 58170 471622 58226
rect 471678 58170 471774 58226
rect 471154 58102 471774 58170
rect 471154 58046 471250 58102
rect 471306 58046 471374 58102
rect 471430 58046 471498 58102
rect 471554 58046 471622 58102
rect 471678 58046 471774 58102
rect 471154 57978 471774 58046
rect 471154 57922 471250 57978
rect 471306 57922 471374 57978
rect 471430 57922 471498 57978
rect 471554 57922 471622 57978
rect 471678 57922 471774 57978
rect 471154 40350 471774 57922
rect 471154 40294 471250 40350
rect 471306 40294 471374 40350
rect 471430 40294 471498 40350
rect 471554 40294 471622 40350
rect 471678 40294 471774 40350
rect 471154 40226 471774 40294
rect 471154 40170 471250 40226
rect 471306 40170 471374 40226
rect 471430 40170 471498 40226
rect 471554 40170 471622 40226
rect 471678 40170 471774 40226
rect 471154 40102 471774 40170
rect 471154 40046 471250 40102
rect 471306 40046 471374 40102
rect 471430 40046 471498 40102
rect 471554 40046 471622 40102
rect 471678 40046 471774 40102
rect 471154 39978 471774 40046
rect 471154 39922 471250 39978
rect 471306 39922 471374 39978
rect 471430 39922 471498 39978
rect 471554 39922 471622 39978
rect 471678 39922 471774 39978
rect 471154 22350 471774 39922
rect 471154 22294 471250 22350
rect 471306 22294 471374 22350
rect 471430 22294 471498 22350
rect 471554 22294 471622 22350
rect 471678 22294 471774 22350
rect 471154 22226 471774 22294
rect 471154 22170 471250 22226
rect 471306 22170 471374 22226
rect 471430 22170 471498 22226
rect 471554 22170 471622 22226
rect 471678 22170 471774 22226
rect 471154 22102 471774 22170
rect 471154 22046 471250 22102
rect 471306 22046 471374 22102
rect 471430 22046 471498 22102
rect 471554 22046 471622 22102
rect 471678 22046 471774 22102
rect 471154 21978 471774 22046
rect 471154 21922 471250 21978
rect 471306 21922 471374 21978
rect 471430 21922 471498 21978
rect 471554 21922 471622 21978
rect 471678 21922 471774 21978
rect 471154 4350 471774 21922
rect 471154 4294 471250 4350
rect 471306 4294 471374 4350
rect 471430 4294 471498 4350
rect 471554 4294 471622 4350
rect 471678 4294 471774 4350
rect 471154 4226 471774 4294
rect 471154 4170 471250 4226
rect 471306 4170 471374 4226
rect 471430 4170 471498 4226
rect 471554 4170 471622 4226
rect 471678 4170 471774 4226
rect 471154 4102 471774 4170
rect 471154 4046 471250 4102
rect 471306 4046 471374 4102
rect 471430 4046 471498 4102
rect 471554 4046 471622 4102
rect 471678 4046 471774 4102
rect 471154 3978 471774 4046
rect 471154 3922 471250 3978
rect 471306 3922 471374 3978
rect 471430 3922 471498 3978
rect 471554 3922 471622 3978
rect 471678 3922 471774 3978
rect 471154 -160 471774 3922
rect 471154 -216 471250 -160
rect 471306 -216 471374 -160
rect 471430 -216 471498 -160
rect 471554 -216 471622 -160
rect 471678 -216 471774 -160
rect 471154 -284 471774 -216
rect 471154 -340 471250 -284
rect 471306 -340 471374 -284
rect 471430 -340 471498 -284
rect 471554 -340 471622 -284
rect 471678 -340 471774 -284
rect 471154 -408 471774 -340
rect 471154 -464 471250 -408
rect 471306 -464 471374 -408
rect 471430 -464 471498 -408
rect 471554 -464 471622 -408
rect 471678 -464 471774 -408
rect 471154 -532 471774 -464
rect 471154 -588 471250 -532
rect 471306 -588 471374 -532
rect 471430 -588 471498 -532
rect 471554 -588 471622 -532
rect 471678 -588 471774 -532
rect 471154 -1644 471774 -588
rect 474874 154350 475494 158858
rect 474874 154294 474970 154350
rect 475026 154294 475094 154350
rect 475150 154294 475218 154350
rect 475274 154294 475342 154350
rect 475398 154294 475494 154350
rect 474874 154226 475494 154294
rect 474874 154170 474970 154226
rect 475026 154170 475094 154226
rect 475150 154170 475218 154226
rect 475274 154170 475342 154226
rect 475398 154170 475494 154226
rect 474874 154102 475494 154170
rect 474874 154046 474970 154102
rect 475026 154046 475094 154102
rect 475150 154046 475218 154102
rect 475274 154046 475342 154102
rect 475398 154046 475494 154102
rect 474874 153978 475494 154046
rect 474874 153922 474970 153978
rect 475026 153922 475094 153978
rect 475150 153922 475218 153978
rect 475274 153922 475342 153978
rect 475398 153922 475494 153978
rect 474874 136350 475494 153922
rect 474874 136294 474970 136350
rect 475026 136294 475094 136350
rect 475150 136294 475218 136350
rect 475274 136294 475342 136350
rect 475398 136294 475494 136350
rect 474874 136226 475494 136294
rect 474874 136170 474970 136226
rect 475026 136170 475094 136226
rect 475150 136170 475218 136226
rect 475274 136170 475342 136226
rect 475398 136170 475494 136226
rect 474874 136102 475494 136170
rect 474874 136046 474970 136102
rect 475026 136046 475094 136102
rect 475150 136046 475218 136102
rect 475274 136046 475342 136102
rect 475398 136046 475494 136102
rect 474874 135978 475494 136046
rect 474874 135922 474970 135978
rect 475026 135922 475094 135978
rect 475150 135922 475218 135978
rect 475274 135922 475342 135978
rect 475398 135922 475494 135978
rect 474874 118350 475494 135922
rect 474874 118294 474970 118350
rect 475026 118294 475094 118350
rect 475150 118294 475218 118350
rect 475274 118294 475342 118350
rect 475398 118294 475494 118350
rect 474874 118226 475494 118294
rect 474874 118170 474970 118226
rect 475026 118170 475094 118226
rect 475150 118170 475218 118226
rect 475274 118170 475342 118226
rect 475398 118170 475494 118226
rect 474874 118102 475494 118170
rect 474874 118046 474970 118102
rect 475026 118046 475094 118102
rect 475150 118046 475218 118102
rect 475274 118046 475342 118102
rect 475398 118046 475494 118102
rect 474874 117978 475494 118046
rect 474874 117922 474970 117978
rect 475026 117922 475094 117978
rect 475150 117922 475218 117978
rect 475274 117922 475342 117978
rect 475398 117922 475494 117978
rect 474874 100350 475494 117922
rect 474874 100294 474970 100350
rect 475026 100294 475094 100350
rect 475150 100294 475218 100350
rect 475274 100294 475342 100350
rect 475398 100294 475494 100350
rect 474874 100226 475494 100294
rect 474874 100170 474970 100226
rect 475026 100170 475094 100226
rect 475150 100170 475218 100226
rect 475274 100170 475342 100226
rect 475398 100170 475494 100226
rect 474874 100102 475494 100170
rect 474874 100046 474970 100102
rect 475026 100046 475094 100102
rect 475150 100046 475218 100102
rect 475274 100046 475342 100102
rect 475398 100046 475494 100102
rect 474874 99978 475494 100046
rect 474874 99922 474970 99978
rect 475026 99922 475094 99978
rect 475150 99922 475218 99978
rect 475274 99922 475342 99978
rect 475398 99922 475494 99978
rect 474874 82350 475494 99922
rect 474874 82294 474970 82350
rect 475026 82294 475094 82350
rect 475150 82294 475218 82350
rect 475274 82294 475342 82350
rect 475398 82294 475494 82350
rect 474874 82226 475494 82294
rect 474874 82170 474970 82226
rect 475026 82170 475094 82226
rect 475150 82170 475218 82226
rect 475274 82170 475342 82226
rect 475398 82170 475494 82226
rect 474874 82102 475494 82170
rect 474874 82046 474970 82102
rect 475026 82046 475094 82102
rect 475150 82046 475218 82102
rect 475274 82046 475342 82102
rect 475398 82046 475494 82102
rect 474874 81978 475494 82046
rect 474874 81922 474970 81978
rect 475026 81922 475094 81978
rect 475150 81922 475218 81978
rect 475274 81922 475342 81978
rect 475398 81922 475494 81978
rect 474874 64350 475494 81922
rect 474874 64294 474970 64350
rect 475026 64294 475094 64350
rect 475150 64294 475218 64350
rect 475274 64294 475342 64350
rect 475398 64294 475494 64350
rect 474874 64226 475494 64294
rect 474874 64170 474970 64226
rect 475026 64170 475094 64226
rect 475150 64170 475218 64226
rect 475274 64170 475342 64226
rect 475398 64170 475494 64226
rect 474874 64102 475494 64170
rect 474874 64046 474970 64102
rect 475026 64046 475094 64102
rect 475150 64046 475218 64102
rect 475274 64046 475342 64102
rect 475398 64046 475494 64102
rect 474874 63978 475494 64046
rect 474874 63922 474970 63978
rect 475026 63922 475094 63978
rect 475150 63922 475218 63978
rect 475274 63922 475342 63978
rect 475398 63922 475494 63978
rect 474874 46350 475494 63922
rect 474874 46294 474970 46350
rect 475026 46294 475094 46350
rect 475150 46294 475218 46350
rect 475274 46294 475342 46350
rect 475398 46294 475494 46350
rect 474874 46226 475494 46294
rect 474874 46170 474970 46226
rect 475026 46170 475094 46226
rect 475150 46170 475218 46226
rect 475274 46170 475342 46226
rect 475398 46170 475494 46226
rect 474874 46102 475494 46170
rect 474874 46046 474970 46102
rect 475026 46046 475094 46102
rect 475150 46046 475218 46102
rect 475274 46046 475342 46102
rect 475398 46046 475494 46102
rect 474874 45978 475494 46046
rect 474874 45922 474970 45978
rect 475026 45922 475094 45978
rect 475150 45922 475218 45978
rect 475274 45922 475342 45978
rect 475398 45922 475494 45978
rect 474874 28350 475494 45922
rect 474874 28294 474970 28350
rect 475026 28294 475094 28350
rect 475150 28294 475218 28350
rect 475274 28294 475342 28350
rect 475398 28294 475494 28350
rect 474874 28226 475494 28294
rect 474874 28170 474970 28226
rect 475026 28170 475094 28226
rect 475150 28170 475218 28226
rect 475274 28170 475342 28226
rect 475398 28170 475494 28226
rect 474874 28102 475494 28170
rect 474874 28046 474970 28102
rect 475026 28046 475094 28102
rect 475150 28046 475218 28102
rect 475274 28046 475342 28102
rect 475398 28046 475494 28102
rect 474874 27978 475494 28046
rect 474874 27922 474970 27978
rect 475026 27922 475094 27978
rect 475150 27922 475218 27978
rect 475274 27922 475342 27978
rect 475398 27922 475494 27978
rect 474874 10350 475494 27922
rect 474874 10294 474970 10350
rect 475026 10294 475094 10350
rect 475150 10294 475218 10350
rect 475274 10294 475342 10350
rect 475398 10294 475494 10350
rect 474874 10226 475494 10294
rect 474874 10170 474970 10226
rect 475026 10170 475094 10226
rect 475150 10170 475218 10226
rect 475274 10170 475342 10226
rect 475398 10170 475494 10226
rect 474874 10102 475494 10170
rect 474874 10046 474970 10102
rect 475026 10046 475094 10102
rect 475150 10046 475218 10102
rect 475274 10046 475342 10102
rect 475398 10046 475494 10102
rect 474874 9978 475494 10046
rect 474874 9922 474970 9978
rect 475026 9922 475094 9978
rect 475150 9922 475218 9978
rect 475274 9922 475342 9978
rect 475398 9922 475494 9978
rect 474874 -1120 475494 9922
rect 474874 -1176 474970 -1120
rect 475026 -1176 475094 -1120
rect 475150 -1176 475218 -1120
rect 475274 -1176 475342 -1120
rect 475398 -1176 475494 -1120
rect 474874 -1244 475494 -1176
rect 474874 -1300 474970 -1244
rect 475026 -1300 475094 -1244
rect 475150 -1300 475218 -1244
rect 475274 -1300 475342 -1244
rect 475398 -1300 475494 -1244
rect 474874 -1368 475494 -1300
rect 474874 -1424 474970 -1368
rect 475026 -1424 475094 -1368
rect 475150 -1424 475218 -1368
rect 475274 -1424 475342 -1368
rect 475398 -1424 475494 -1368
rect 474874 -1492 475494 -1424
rect 474874 -1548 474970 -1492
rect 475026 -1548 475094 -1492
rect 475150 -1548 475218 -1492
rect 475274 -1548 475342 -1492
rect 475398 -1548 475494 -1492
rect 474874 -1644 475494 -1548
rect 489154 148350 489774 158858
rect 489154 148294 489250 148350
rect 489306 148294 489374 148350
rect 489430 148294 489498 148350
rect 489554 148294 489622 148350
rect 489678 148294 489774 148350
rect 489154 148226 489774 148294
rect 489154 148170 489250 148226
rect 489306 148170 489374 148226
rect 489430 148170 489498 148226
rect 489554 148170 489622 148226
rect 489678 148170 489774 148226
rect 489154 148102 489774 148170
rect 489154 148046 489250 148102
rect 489306 148046 489374 148102
rect 489430 148046 489498 148102
rect 489554 148046 489622 148102
rect 489678 148046 489774 148102
rect 489154 147978 489774 148046
rect 489154 147922 489250 147978
rect 489306 147922 489374 147978
rect 489430 147922 489498 147978
rect 489554 147922 489622 147978
rect 489678 147922 489774 147978
rect 489154 130350 489774 147922
rect 489154 130294 489250 130350
rect 489306 130294 489374 130350
rect 489430 130294 489498 130350
rect 489554 130294 489622 130350
rect 489678 130294 489774 130350
rect 489154 130226 489774 130294
rect 489154 130170 489250 130226
rect 489306 130170 489374 130226
rect 489430 130170 489498 130226
rect 489554 130170 489622 130226
rect 489678 130170 489774 130226
rect 489154 130102 489774 130170
rect 489154 130046 489250 130102
rect 489306 130046 489374 130102
rect 489430 130046 489498 130102
rect 489554 130046 489622 130102
rect 489678 130046 489774 130102
rect 489154 129978 489774 130046
rect 489154 129922 489250 129978
rect 489306 129922 489374 129978
rect 489430 129922 489498 129978
rect 489554 129922 489622 129978
rect 489678 129922 489774 129978
rect 489154 112350 489774 129922
rect 489154 112294 489250 112350
rect 489306 112294 489374 112350
rect 489430 112294 489498 112350
rect 489554 112294 489622 112350
rect 489678 112294 489774 112350
rect 489154 112226 489774 112294
rect 489154 112170 489250 112226
rect 489306 112170 489374 112226
rect 489430 112170 489498 112226
rect 489554 112170 489622 112226
rect 489678 112170 489774 112226
rect 489154 112102 489774 112170
rect 489154 112046 489250 112102
rect 489306 112046 489374 112102
rect 489430 112046 489498 112102
rect 489554 112046 489622 112102
rect 489678 112046 489774 112102
rect 489154 111978 489774 112046
rect 489154 111922 489250 111978
rect 489306 111922 489374 111978
rect 489430 111922 489498 111978
rect 489554 111922 489622 111978
rect 489678 111922 489774 111978
rect 489154 94350 489774 111922
rect 489154 94294 489250 94350
rect 489306 94294 489374 94350
rect 489430 94294 489498 94350
rect 489554 94294 489622 94350
rect 489678 94294 489774 94350
rect 489154 94226 489774 94294
rect 489154 94170 489250 94226
rect 489306 94170 489374 94226
rect 489430 94170 489498 94226
rect 489554 94170 489622 94226
rect 489678 94170 489774 94226
rect 489154 94102 489774 94170
rect 489154 94046 489250 94102
rect 489306 94046 489374 94102
rect 489430 94046 489498 94102
rect 489554 94046 489622 94102
rect 489678 94046 489774 94102
rect 489154 93978 489774 94046
rect 489154 93922 489250 93978
rect 489306 93922 489374 93978
rect 489430 93922 489498 93978
rect 489554 93922 489622 93978
rect 489678 93922 489774 93978
rect 489154 76350 489774 93922
rect 489154 76294 489250 76350
rect 489306 76294 489374 76350
rect 489430 76294 489498 76350
rect 489554 76294 489622 76350
rect 489678 76294 489774 76350
rect 489154 76226 489774 76294
rect 489154 76170 489250 76226
rect 489306 76170 489374 76226
rect 489430 76170 489498 76226
rect 489554 76170 489622 76226
rect 489678 76170 489774 76226
rect 489154 76102 489774 76170
rect 489154 76046 489250 76102
rect 489306 76046 489374 76102
rect 489430 76046 489498 76102
rect 489554 76046 489622 76102
rect 489678 76046 489774 76102
rect 489154 75978 489774 76046
rect 489154 75922 489250 75978
rect 489306 75922 489374 75978
rect 489430 75922 489498 75978
rect 489554 75922 489622 75978
rect 489678 75922 489774 75978
rect 489154 58350 489774 75922
rect 489154 58294 489250 58350
rect 489306 58294 489374 58350
rect 489430 58294 489498 58350
rect 489554 58294 489622 58350
rect 489678 58294 489774 58350
rect 489154 58226 489774 58294
rect 489154 58170 489250 58226
rect 489306 58170 489374 58226
rect 489430 58170 489498 58226
rect 489554 58170 489622 58226
rect 489678 58170 489774 58226
rect 489154 58102 489774 58170
rect 489154 58046 489250 58102
rect 489306 58046 489374 58102
rect 489430 58046 489498 58102
rect 489554 58046 489622 58102
rect 489678 58046 489774 58102
rect 489154 57978 489774 58046
rect 489154 57922 489250 57978
rect 489306 57922 489374 57978
rect 489430 57922 489498 57978
rect 489554 57922 489622 57978
rect 489678 57922 489774 57978
rect 489154 40350 489774 57922
rect 489154 40294 489250 40350
rect 489306 40294 489374 40350
rect 489430 40294 489498 40350
rect 489554 40294 489622 40350
rect 489678 40294 489774 40350
rect 489154 40226 489774 40294
rect 489154 40170 489250 40226
rect 489306 40170 489374 40226
rect 489430 40170 489498 40226
rect 489554 40170 489622 40226
rect 489678 40170 489774 40226
rect 489154 40102 489774 40170
rect 489154 40046 489250 40102
rect 489306 40046 489374 40102
rect 489430 40046 489498 40102
rect 489554 40046 489622 40102
rect 489678 40046 489774 40102
rect 489154 39978 489774 40046
rect 489154 39922 489250 39978
rect 489306 39922 489374 39978
rect 489430 39922 489498 39978
rect 489554 39922 489622 39978
rect 489678 39922 489774 39978
rect 489154 22350 489774 39922
rect 489154 22294 489250 22350
rect 489306 22294 489374 22350
rect 489430 22294 489498 22350
rect 489554 22294 489622 22350
rect 489678 22294 489774 22350
rect 489154 22226 489774 22294
rect 489154 22170 489250 22226
rect 489306 22170 489374 22226
rect 489430 22170 489498 22226
rect 489554 22170 489622 22226
rect 489678 22170 489774 22226
rect 489154 22102 489774 22170
rect 489154 22046 489250 22102
rect 489306 22046 489374 22102
rect 489430 22046 489498 22102
rect 489554 22046 489622 22102
rect 489678 22046 489774 22102
rect 489154 21978 489774 22046
rect 489154 21922 489250 21978
rect 489306 21922 489374 21978
rect 489430 21922 489498 21978
rect 489554 21922 489622 21978
rect 489678 21922 489774 21978
rect 489154 4350 489774 21922
rect 489154 4294 489250 4350
rect 489306 4294 489374 4350
rect 489430 4294 489498 4350
rect 489554 4294 489622 4350
rect 489678 4294 489774 4350
rect 489154 4226 489774 4294
rect 489154 4170 489250 4226
rect 489306 4170 489374 4226
rect 489430 4170 489498 4226
rect 489554 4170 489622 4226
rect 489678 4170 489774 4226
rect 489154 4102 489774 4170
rect 489154 4046 489250 4102
rect 489306 4046 489374 4102
rect 489430 4046 489498 4102
rect 489554 4046 489622 4102
rect 489678 4046 489774 4102
rect 489154 3978 489774 4046
rect 489154 3922 489250 3978
rect 489306 3922 489374 3978
rect 489430 3922 489498 3978
rect 489554 3922 489622 3978
rect 489678 3922 489774 3978
rect 489154 -160 489774 3922
rect 489154 -216 489250 -160
rect 489306 -216 489374 -160
rect 489430 -216 489498 -160
rect 489554 -216 489622 -160
rect 489678 -216 489774 -160
rect 489154 -284 489774 -216
rect 489154 -340 489250 -284
rect 489306 -340 489374 -284
rect 489430 -340 489498 -284
rect 489554 -340 489622 -284
rect 489678 -340 489774 -284
rect 489154 -408 489774 -340
rect 489154 -464 489250 -408
rect 489306 -464 489374 -408
rect 489430 -464 489498 -408
rect 489554 -464 489622 -408
rect 489678 -464 489774 -408
rect 489154 -532 489774 -464
rect 489154 -588 489250 -532
rect 489306 -588 489374 -532
rect 489430 -588 489498 -532
rect 489554 -588 489622 -532
rect 489678 -588 489774 -532
rect 489154 -1644 489774 -588
rect 492874 154350 493494 158858
rect 492874 154294 492970 154350
rect 493026 154294 493094 154350
rect 493150 154294 493218 154350
rect 493274 154294 493342 154350
rect 493398 154294 493494 154350
rect 492874 154226 493494 154294
rect 492874 154170 492970 154226
rect 493026 154170 493094 154226
rect 493150 154170 493218 154226
rect 493274 154170 493342 154226
rect 493398 154170 493494 154226
rect 492874 154102 493494 154170
rect 492874 154046 492970 154102
rect 493026 154046 493094 154102
rect 493150 154046 493218 154102
rect 493274 154046 493342 154102
rect 493398 154046 493494 154102
rect 492874 153978 493494 154046
rect 492874 153922 492970 153978
rect 493026 153922 493094 153978
rect 493150 153922 493218 153978
rect 493274 153922 493342 153978
rect 493398 153922 493494 153978
rect 492874 136350 493494 153922
rect 492874 136294 492970 136350
rect 493026 136294 493094 136350
rect 493150 136294 493218 136350
rect 493274 136294 493342 136350
rect 493398 136294 493494 136350
rect 492874 136226 493494 136294
rect 492874 136170 492970 136226
rect 493026 136170 493094 136226
rect 493150 136170 493218 136226
rect 493274 136170 493342 136226
rect 493398 136170 493494 136226
rect 492874 136102 493494 136170
rect 492874 136046 492970 136102
rect 493026 136046 493094 136102
rect 493150 136046 493218 136102
rect 493274 136046 493342 136102
rect 493398 136046 493494 136102
rect 492874 135978 493494 136046
rect 492874 135922 492970 135978
rect 493026 135922 493094 135978
rect 493150 135922 493218 135978
rect 493274 135922 493342 135978
rect 493398 135922 493494 135978
rect 492874 118350 493494 135922
rect 492874 118294 492970 118350
rect 493026 118294 493094 118350
rect 493150 118294 493218 118350
rect 493274 118294 493342 118350
rect 493398 118294 493494 118350
rect 492874 118226 493494 118294
rect 492874 118170 492970 118226
rect 493026 118170 493094 118226
rect 493150 118170 493218 118226
rect 493274 118170 493342 118226
rect 493398 118170 493494 118226
rect 492874 118102 493494 118170
rect 492874 118046 492970 118102
rect 493026 118046 493094 118102
rect 493150 118046 493218 118102
rect 493274 118046 493342 118102
rect 493398 118046 493494 118102
rect 492874 117978 493494 118046
rect 492874 117922 492970 117978
rect 493026 117922 493094 117978
rect 493150 117922 493218 117978
rect 493274 117922 493342 117978
rect 493398 117922 493494 117978
rect 492874 100350 493494 117922
rect 492874 100294 492970 100350
rect 493026 100294 493094 100350
rect 493150 100294 493218 100350
rect 493274 100294 493342 100350
rect 493398 100294 493494 100350
rect 492874 100226 493494 100294
rect 492874 100170 492970 100226
rect 493026 100170 493094 100226
rect 493150 100170 493218 100226
rect 493274 100170 493342 100226
rect 493398 100170 493494 100226
rect 492874 100102 493494 100170
rect 492874 100046 492970 100102
rect 493026 100046 493094 100102
rect 493150 100046 493218 100102
rect 493274 100046 493342 100102
rect 493398 100046 493494 100102
rect 492874 99978 493494 100046
rect 492874 99922 492970 99978
rect 493026 99922 493094 99978
rect 493150 99922 493218 99978
rect 493274 99922 493342 99978
rect 493398 99922 493494 99978
rect 492874 82350 493494 99922
rect 492874 82294 492970 82350
rect 493026 82294 493094 82350
rect 493150 82294 493218 82350
rect 493274 82294 493342 82350
rect 493398 82294 493494 82350
rect 492874 82226 493494 82294
rect 492874 82170 492970 82226
rect 493026 82170 493094 82226
rect 493150 82170 493218 82226
rect 493274 82170 493342 82226
rect 493398 82170 493494 82226
rect 492874 82102 493494 82170
rect 492874 82046 492970 82102
rect 493026 82046 493094 82102
rect 493150 82046 493218 82102
rect 493274 82046 493342 82102
rect 493398 82046 493494 82102
rect 492874 81978 493494 82046
rect 492874 81922 492970 81978
rect 493026 81922 493094 81978
rect 493150 81922 493218 81978
rect 493274 81922 493342 81978
rect 493398 81922 493494 81978
rect 492874 64350 493494 81922
rect 492874 64294 492970 64350
rect 493026 64294 493094 64350
rect 493150 64294 493218 64350
rect 493274 64294 493342 64350
rect 493398 64294 493494 64350
rect 492874 64226 493494 64294
rect 492874 64170 492970 64226
rect 493026 64170 493094 64226
rect 493150 64170 493218 64226
rect 493274 64170 493342 64226
rect 493398 64170 493494 64226
rect 492874 64102 493494 64170
rect 492874 64046 492970 64102
rect 493026 64046 493094 64102
rect 493150 64046 493218 64102
rect 493274 64046 493342 64102
rect 493398 64046 493494 64102
rect 492874 63978 493494 64046
rect 492874 63922 492970 63978
rect 493026 63922 493094 63978
rect 493150 63922 493218 63978
rect 493274 63922 493342 63978
rect 493398 63922 493494 63978
rect 492874 46350 493494 63922
rect 492874 46294 492970 46350
rect 493026 46294 493094 46350
rect 493150 46294 493218 46350
rect 493274 46294 493342 46350
rect 493398 46294 493494 46350
rect 492874 46226 493494 46294
rect 492874 46170 492970 46226
rect 493026 46170 493094 46226
rect 493150 46170 493218 46226
rect 493274 46170 493342 46226
rect 493398 46170 493494 46226
rect 492874 46102 493494 46170
rect 492874 46046 492970 46102
rect 493026 46046 493094 46102
rect 493150 46046 493218 46102
rect 493274 46046 493342 46102
rect 493398 46046 493494 46102
rect 492874 45978 493494 46046
rect 492874 45922 492970 45978
rect 493026 45922 493094 45978
rect 493150 45922 493218 45978
rect 493274 45922 493342 45978
rect 493398 45922 493494 45978
rect 492874 28350 493494 45922
rect 492874 28294 492970 28350
rect 493026 28294 493094 28350
rect 493150 28294 493218 28350
rect 493274 28294 493342 28350
rect 493398 28294 493494 28350
rect 492874 28226 493494 28294
rect 492874 28170 492970 28226
rect 493026 28170 493094 28226
rect 493150 28170 493218 28226
rect 493274 28170 493342 28226
rect 493398 28170 493494 28226
rect 492874 28102 493494 28170
rect 492874 28046 492970 28102
rect 493026 28046 493094 28102
rect 493150 28046 493218 28102
rect 493274 28046 493342 28102
rect 493398 28046 493494 28102
rect 492874 27978 493494 28046
rect 492874 27922 492970 27978
rect 493026 27922 493094 27978
rect 493150 27922 493218 27978
rect 493274 27922 493342 27978
rect 493398 27922 493494 27978
rect 492874 10350 493494 27922
rect 492874 10294 492970 10350
rect 493026 10294 493094 10350
rect 493150 10294 493218 10350
rect 493274 10294 493342 10350
rect 493398 10294 493494 10350
rect 492874 10226 493494 10294
rect 492874 10170 492970 10226
rect 493026 10170 493094 10226
rect 493150 10170 493218 10226
rect 493274 10170 493342 10226
rect 493398 10170 493494 10226
rect 492874 10102 493494 10170
rect 492874 10046 492970 10102
rect 493026 10046 493094 10102
rect 493150 10046 493218 10102
rect 493274 10046 493342 10102
rect 493398 10046 493494 10102
rect 492874 9978 493494 10046
rect 492874 9922 492970 9978
rect 493026 9922 493094 9978
rect 493150 9922 493218 9978
rect 493274 9922 493342 9978
rect 493398 9922 493494 9978
rect 492874 -1120 493494 9922
rect 492874 -1176 492970 -1120
rect 493026 -1176 493094 -1120
rect 493150 -1176 493218 -1120
rect 493274 -1176 493342 -1120
rect 493398 -1176 493494 -1120
rect 492874 -1244 493494 -1176
rect 492874 -1300 492970 -1244
rect 493026 -1300 493094 -1244
rect 493150 -1300 493218 -1244
rect 493274 -1300 493342 -1244
rect 493398 -1300 493494 -1244
rect 492874 -1368 493494 -1300
rect 492874 -1424 492970 -1368
rect 493026 -1424 493094 -1368
rect 493150 -1424 493218 -1368
rect 493274 -1424 493342 -1368
rect 493398 -1424 493494 -1368
rect 492874 -1492 493494 -1424
rect 492874 -1548 492970 -1492
rect 493026 -1548 493094 -1492
rect 493150 -1548 493218 -1492
rect 493274 -1548 493342 -1492
rect 493398 -1548 493494 -1492
rect 492874 -1644 493494 -1548
rect 507154 148350 507774 158858
rect 507154 148294 507250 148350
rect 507306 148294 507374 148350
rect 507430 148294 507498 148350
rect 507554 148294 507622 148350
rect 507678 148294 507774 148350
rect 507154 148226 507774 148294
rect 507154 148170 507250 148226
rect 507306 148170 507374 148226
rect 507430 148170 507498 148226
rect 507554 148170 507622 148226
rect 507678 148170 507774 148226
rect 507154 148102 507774 148170
rect 507154 148046 507250 148102
rect 507306 148046 507374 148102
rect 507430 148046 507498 148102
rect 507554 148046 507622 148102
rect 507678 148046 507774 148102
rect 507154 147978 507774 148046
rect 507154 147922 507250 147978
rect 507306 147922 507374 147978
rect 507430 147922 507498 147978
rect 507554 147922 507622 147978
rect 507678 147922 507774 147978
rect 507154 130350 507774 147922
rect 507154 130294 507250 130350
rect 507306 130294 507374 130350
rect 507430 130294 507498 130350
rect 507554 130294 507622 130350
rect 507678 130294 507774 130350
rect 507154 130226 507774 130294
rect 507154 130170 507250 130226
rect 507306 130170 507374 130226
rect 507430 130170 507498 130226
rect 507554 130170 507622 130226
rect 507678 130170 507774 130226
rect 507154 130102 507774 130170
rect 507154 130046 507250 130102
rect 507306 130046 507374 130102
rect 507430 130046 507498 130102
rect 507554 130046 507622 130102
rect 507678 130046 507774 130102
rect 507154 129978 507774 130046
rect 507154 129922 507250 129978
rect 507306 129922 507374 129978
rect 507430 129922 507498 129978
rect 507554 129922 507622 129978
rect 507678 129922 507774 129978
rect 507154 112350 507774 129922
rect 507154 112294 507250 112350
rect 507306 112294 507374 112350
rect 507430 112294 507498 112350
rect 507554 112294 507622 112350
rect 507678 112294 507774 112350
rect 507154 112226 507774 112294
rect 507154 112170 507250 112226
rect 507306 112170 507374 112226
rect 507430 112170 507498 112226
rect 507554 112170 507622 112226
rect 507678 112170 507774 112226
rect 507154 112102 507774 112170
rect 507154 112046 507250 112102
rect 507306 112046 507374 112102
rect 507430 112046 507498 112102
rect 507554 112046 507622 112102
rect 507678 112046 507774 112102
rect 507154 111978 507774 112046
rect 507154 111922 507250 111978
rect 507306 111922 507374 111978
rect 507430 111922 507498 111978
rect 507554 111922 507622 111978
rect 507678 111922 507774 111978
rect 507154 94350 507774 111922
rect 507154 94294 507250 94350
rect 507306 94294 507374 94350
rect 507430 94294 507498 94350
rect 507554 94294 507622 94350
rect 507678 94294 507774 94350
rect 507154 94226 507774 94294
rect 507154 94170 507250 94226
rect 507306 94170 507374 94226
rect 507430 94170 507498 94226
rect 507554 94170 507622 94226
rect 507678 94170 507774 94226
rect 507154 94102 507774 94170
rect 507154 94046 507250 94102
rect 507306 94046 507374 94102
rect 507430 94046 507498 94102
rect 507554 94046 507622 94102
rect 507678 94046 507774 94102
rect 507154 93978 507774 94046
rect 507154 93922 507250 93978
rect 507306 93922 507374 93978
rect 507430 93922 507498 93978
rect 507554 93922 507622 93978
rect 507678 93922 507774 93978
rect 507154 76350 507774 93922
rect 507154 76294 507250 76350
rect 507306 76294 507374 76350
rect 507430 76294 507498 76350
rect 507554 76294 507622 76350
rect 507678 76294 507774 76350
rect 507154 76226 507774 76294
rect 507154 76170 507250 76226
rect 507306 76170 507374 76226
rect 507430 76170 507498 76226
rect 507554 76170 507622 76226
rect 507678 76170 507774 76226
rect 507154 76102 507774 76170
rect 507154 76046 507250 76102
rect 507306 76046 507374 76102
rect 507430 76046 507498 76102
rect 507554 76046 507622 76102
rect 507678 76046 507774 76102
rect 507154 75978 507774 76046
rect 507154 75922 507250 75978
rect 507306 75922 507374 75978
rect 507430 75922 507498 75978
rect 507554 75922 507622 75978
rect 507678 75922 507774 75978
rect 507154 58350 507774 75922
rect 507154 58294 507250 58350
rect 507306 58294 507374 58350
rect 507430 58294 507498 58350
rect 507554 58294 507622 58350
rect 507678 58294 507774 58350
rect 507154 58226 507774 58294
rect 507154 58170 507250 58226
rect 507306 58170 507374 58226
rect 507430 58170 507498 58226
rect 507554 58170 507622 58226
rect 507678 58170 507774 58226
rect 507154 58102 507774 58170
rect 507154 58046 507250 58102
rect 507306 58046 507374 58102
rect 507430 58046 507498 58102
rect 507554 58046 507622 58102
rect 507678 58046 507774 58102
rect 507154 57978 507774 58046
rect 507154 57922 507250 57978
rect 507306 57922 507374 57978
rect 507430 57922 507498 57978
rect 507554 57922 507622 57978
rect 507678 57922 507774 57978
rect 507154 40350 507774 57922
rect 507154 40294 507250 40350
rect 507306 40294 507374 40350
rect 507430 40294 507498 40350
rect 507554 40294 507622 40350
rect 507678 40294 507774 40350
rect 507154 40226 507774 40294
rect 507154 40170 507250 40226
rect 507306 40170 507374 40226
rect 507430 40170 507498 40226
rect 507554 40170 507622 40226
rect 507678 40170 507774 40226
rect 507154 40102 507774 40170
rect 507154 40046 507250 40102
rect 507306 40046 507374 40102
rect 507430 40046 507498 40102
rect 507554 40046 507622 40102
rect 507678 40046 507774 40102
rect 507154 39978 507774 40046
rect 507154 39922 507250 39978
rect 507306 39922 507374 39978
rect 507430 39922 507498 39978
rect 507554 39922 507622 39978
rect 507678 39922 507774 39978
rect 507154 22350 507774 39922
rect 507154 22294 507250 22350
rect 507306 22294 507374 22350
rect 507430 22294 507498 22350
rect 507554 22294 507622 22350
rect 507678 22294 507774 22350
rect 507154 22226 507774 22294
rect 507154 22170 507250 22226
rect 507306 22170 507374 22226
rect 507430 22170 507498 22226
rect 507554 22170 507622 22226
rect 507678 22170 507774 22226
rect 507154 22102 507774 22170
rect 507154 22046 507250 22102
rect 507306 22046 507374 22102
rect 507430 22046 507498 22102
rect 507554 22046 507622 22102
rect 507678 22046 507774 22102
rect 507154 21978 507774 22046
rect 507154 21922 507250 21978
rect 507306 21922 507374 21978
rect 507430 21922 507498 21978
rect 507554 21922 507622 21978
rect 507678 21922 507774 21978
rect 507154 4350 507774 21922
rect 507154 4294 507250 4350
rect 507306 4294 507374 4350
rect 507430 4294 507498 4350
rect 507554 4294 507622 4350
rect 507678 4294 507774 4350
rect 507154 4226 507774 4294
rect 507154 4170 507250 4226
rect 507306 4170 507374 4226
rect 507430 4170 507498 4226
rect 507554 4170 507622 4226
rect 507678 4170 507774 4226
rect 507154 4102 507774 4170
rect 507154 4046 507250 4102
rect 507306 4046 507374 4102
rect 507430 4046 507498 4102
rect 507554 4046 507622 4102
rect 507678 4046 507774 4102
rect 507154 3978 507774 4046
rect 507154 3922 507250 3978
rect 507306 3922 507374 3978
rect 507430 3922 507498 3978
rect 507554 3922 507622 3978
rect 507678 3922 507774 3978
rect 507154 -160 507774 3922
rect 507154 -216 507250 -160
rect 507306 -216 507374 -160
rect 507430 -216 507498 -160
rect 507554 -216 507622 -160
rect 507678 -216 507774 -160
rect 507154 -284 507774 -216
rect 507154 -340 507250 -284
rect 507306 -340 507374 -284
rect 507430 -340 507498 -284
rect 507554 -340 507622 -284
rect 507678 -340 507774 -284
rect 507154 -408 507774 -340
rect 507154 -464 507250 -408
rect 507306 -464 507374 -408
rect 507430 -464 507498 -408
rect 507554 -464 507622 -408
rect 507678 -464 507774 -408
rect 507154 -532 507774 -464
rect 507154 -588 507250 -532
rect 507306 -588 507374 -532
rect 507430 -588 507498 -532
rect 507554 -588 507622 -532
rect 507678 -588 507774 -532
rect 507154 -1644 507774 -588
rect 510874 154350 511494 158858
rect 510874 154294 510970 154350
rect 511026 154294 511094 154350
rect 511150 154294 511218 154350
rect 511274 154294 511342 154350
rect 511398 154294 511494 154350
rect 510874 154226 511494 154294
rect 510874 154170 510970 154226
rect 511026 154170 511094 154226
rect 511150 154170 511218 154226
rect 511274 154170 511342 154226
rect 511398 154170 511494 154226
rect 510874 154102 511494 154170
rect 510874 154046 510970 154102
rect 511026 154046 511094 154102
rect 511150 154046 511218 154102
rect 511274 154046 511342 154102
rect 511398 154046 511494 154102
rect 510874 153978 511494 154046
rect 510874 153922 510970 153978
rect 511026 153922 511094 153978
rect 511150 153922 511218 153978
rect 511274 153922 511342 153978
rect 511398 153922 511494 153978
rect 510874 136350 511494 153922
rect 510874 136294 510970 136350
rect 511026 136294 511094 136350
rect 511150 136294 511218 136350
rect 511274 136294 511342 136350
rect 511398 136294 511494 136350
rect 510874 136226 511494 136294
rect 510874 136170 510970 136226
rect 511026 136170 511094 136226
rect 511150 136170 511218 136226
rect 511274 136170 511342 136226
rect 511398 136170 511494 136226
rect 510874 136102 511494 136170
rect 510874 136046 510970 136102
rect 511026 136046 511094 136102
rect 511150 136046 511218 136102
rect 511274 136046 511342 136102
rect 511398 136046 511494 136102
rect 510874 135978 511494 136046
rect 510874 135922 510970 135978
rect 511026 135922 511094 135978
rect 511150 135922 511218 135978
rect 511274 135922 511342 135978
rect 511398 135922 511494 135978
rect 510874 118350 511494 135922
rect 510874 118294 510970 118350
rect 511026 118294 511094 118350
rect 511150 118294 511218 118350
rect 511274 118294 511342 118350
rect 511398 118294 511494 118350
rect 510874 118226 511494 118294
rect 510874 118170 510970 118226
rect 511026 118170 511094 118226
rect 511150 118170 511218 118226
rect 511274 118170 511342 118226
rect 511398 118170 511494 118226
rect 510874 118102 511494 118170
rect 510874 118046 510970 118102
rect 511026 118046 511094 118102
rect 511150 118046 511218 118102
rect 511274 118046 511342 118102
rect 511398 118046 511494 118102
rect 510874 117978 511494 118046
rect 510874 117922 510970 117978
rect 511026 117922 511094 117978
rect 511150 117922 511218 117978
rect 511274 117922 511342 117978
rect 511398 117922 511494 117978
rect 510874 100350 511494 117922
rect 510874 100294 510970 100350
rect 511026 100294 511094 100350
rect 511150 100294 511218 100350
rect 511274 100294 511342 100350
rect 511398 100294 511494 100350
rect 510874 100226 511494 100294
rect 510874 100170 510970 100226
rect 511026 100170 511094 100226
rect 511150 100170 511218 100226
rect 511274 100170 511342 100226
rect 511398 100170 511494 100226
rect 510874 100102 511494 100170
rect 510874 100046 510970 100102
rect 511026 100046 511094 100102
rect 511150 100046 511218 100102
rect 511274 100046 511342 100102
rect 511398 100046 511494 100102
rect 510874 99978 511494 100046
rect 510874 99922 510970 99978
rect 511026 99922 511094 99978
rect 511150 99922 511218 99978
rect 511274 99922 511342 99978
rect 511398 99922 511494 99978
rect 510874 82350 511494 99922
rect 525154 148350 525774 158858
rect 525154 148294 525250 148350
rect 525306 148294 525374 148350
rect 525430 148294 525498 148350
rect 525554 148294 525622 148350
rect 525678 148294 525774 148350
rect 525154 148226 525774 148294
rect 525154 148170 525250 148226
rect 525306 148170 525374 148226
rect 525430 148170 525498 148226
rect 525554 148170 525622 148226
rect 525678 148170 525774 148226
rect 525154 148102 525774 148170
rect 525154 148046 525250 148102
rect 525306 148046 525374 148102
rect 525430 148046 525498 148102
rect 525554 148046 525622 148102
rect 525678 148046 525774 148102
rect 525154 147978 525774 148046
rect 525154 147922 525250 147978
rect 525306 147922 525374 147978
rect 525430 147922 525498 147978
rect 525554 147922 525622 147978
rect 525678 147922 525774 147978
rect 525154 130350 525774 147922
rect 525154 130294 525250 130350
rect 525306 130294 525374 130350
rect 525430 130294 525498 130350
rect 525554 130294 525622 130350
rect 525678 130294 525774 130350
rect 525154 130226 525774 130294
rect 525154 130170 525250 130226
rect 525306 130170 525374 130226
rect 525430 130170 525498 130226
rect 525554 130170 525622 130226
rect 525678 130170 525774 130226
rect 525154 130102 525774 130170
rect 525154 130046 525250 130102
rect 525306 130046 525374 130102
rect 525430 130046 525498 130102
rect 525554 130046 525622 130102
rect 525678 130046 525774 130102
rect 525154 129978 525774 130046
rect 525154 129922 525250 129978
rect 525306 129922 525374 129978
rect 525430 129922 525498 129978
rect 525554 129922 525622 129978
rect 525678 129922 525774 129978
rect 525154 112350 525774 129922
rect 525154 112294 525250 112350
rect 525306 112294 525374 112350
rect 525430 112294 525498 112350
rect 525554 112294 525622 112350
rect 525678 112294 525774 112350
rect 525154 112226 525774 112294
rect 525154 112170 525250 112226
rect 525306 112170 525374 112226
rect 525430 112170 525498 112226
rect 525554 112170 525622 112226
rect 525678 112170 525774 112226
rect 525154 112102 525774 112170
rect 525154 112046 525250 112102
rect 525306 112046 525374 112102
rect 525430 112046 525498 112102
rect 525554 112046 525622 112102
rect 525678 112046 525774 112102
rect 525154 111978 525774 112046
rect 525154 111922 525250 111978
rect 525306 111922 525374 111978
rect 525430 111922 525498 111978
rect 525554 111922 525622 111978
rect 525678 111922 525774 111978
rect 524448 94350 524768 94384
rect 524448 94294 524518 94350
rect 524574 94294 524642 94350
rect 524698 94294 524768 94350
rect 524448 94226 524768 94294
rect 524448 94170 524518 94226
rect 524574 94170 524642 94226
rect 524698 94170 524768 94226
rect 524448 94102 524768 94170
rect 524448 94046 524518 94102
rect 524574 94046 524642 94102
rect 524698 94046 524768 94102
rect 524448 93978 524768 94046
rect 524448 93922 524518 93978
rect 524574 93922 524642 93978
rect 524698 93922 524768 93978
rect 524448 93888 524768 93922
rect 525154 94350 525774 111922
rect 525154 94294 525250 94350
rect 525306 94294 525374 94350
rect 525430 94294 525498 94350
rect 525554 94294 525622 94350
rect 525678 94294 525774 94350
rect 525154 94226 525774 94294
rect 525154 94170 525250 94226
rect 525306 94170 525374 94226
rect 525430 94170 525498 94226
rect 525554 94170 525622 94226
rect 525678 94170 525774 94226
rect 525154 94102 525774 94170
rect 525154 94046 525250 94102
rect 525306 94046 525374 94102
rect 525430 94046 525498 94102
rect 525554 94046 525622 94102
rect 525678 94046 525774 94102
rect 525154 93978 525774 94046
rect 525154 93922 525250 93978
rect 525306 93922 525374 93978
rect 525430 93922 525498 93978
rect 525554 93922 525622 93978
rect 525678 93922 525774 93978
rect 510874 82294 510970 82350
rect 511026 82294 511094 82350
rect 511150 82294 511218 82350
rect 511274 82294 511342 82350
rect 511398 82294 511494 82350
rect 510874 82226 511494 82294
rect 510874 82170 510970 82226
rect 511026 82170 511094 82226
rect 511150 82170 511218 82226
rect 511274 82170 511342 82226
rect 511398 82170 511494 82226
rect 510874 82102 511494 82170
rect 510874 82046 510970 82102
rect 511026 82046 511094 82102
rect 511150 82046 511218 82102
rect 511274 82046 511342 82102
rect 511398 82046 511494 82102
rect 510874 81978 511494 82046
rect 510874 81922 510970 81978
rect 511026 81922 511094 81978
rect 511150 81922 511218 81978
rect 511274 81922 511342 81978
rect 511398 81922 511494 81978
rect 510874 64350 511494 81922
rect 524448 76350 524768 76384
rect 524448 76294 524518 76350
rect 524574 76294 524642 76350
rect 524698 76294 524768 76350
rect 524448 76226 524768 76294
rect 524448 76170 524518 76226
rect 524574 76170 524642 76226
rect 524698 76170 524768 76226
rect 524448 76102 524768 76170
rect 524448 76046 524518 76102
rect 524574 76046 524642 76102
rect 524698 76046 524768 76102
rect 524448 75978 524768 76046
rect 524448 75922 524518 75978
rect 524574 75922 524642 75978
rect 524698 75922 524768 75978
rect 524448 75888 524768 75922
rect 525154 76350 525774 93922
rect 525154 76294 525250 76350
rect 525306 76294 525374 76350
rect 525430 76294 525498 76350
rect 525554 76294 525622 76350
rect 525678 76294 525774 76350
rect 525154 76226 525774 76294
rect 525154 76170 525250 76226
rect 525306 76170 525374 76226
rect 525430 76170 525498 76226
rect 525554 76170 525622 76226
rect 525678 76170 525774 76226
rect 525154 76102 525774 76170
rect 525154 76046 525250 76102
rect 525306 76046 525374 76102
rect 525430 76046 525498 76102
rect 525554 76046 525622 76102
rect 525678 76046 525774 76102
rect 525154 75978 525774 76046
rect 525154 75922 525250 75978
rect 525306 75922 525374 75978
rect 525430 75922 525498 75978
rect 525554 75922 525622 75978
rect 525678 75922 525774 75978
rect 510874 64294 510970 64350
rect 511026 64294 511094 64350
rect 511150 64294 511218 64350
rect 511274 64294 511342 64350
rect 511398 64294 511494 64350
rect 510874 64226 511494 64294
rect 510874 64170 510970 64226
rect 511026 64170 511094 64226
rect 511150 64170 511218 64226
rect 511274 64170 511342 64226
rect 511398 64170 511494 64226
rect 510874 64102 511494 64170
rect 510874 64046 510970 64102
rect 511026 64046 511094 64102
rect 511150 64046 511218 64102
rect 511274 64046 511342 64102
rect 511398 64046 511494 64102
rect 510874 63978 511494 64046
rect 510874 63922 510970 63978
rect 511026 63922 511094 63978
rect 511150 63922 511218 63978
rect 511274 63922 511342 63978
rect 511398 63922 511494 63978
rect 510874 46350 511494 63922
rect 510874 46294 510970 46350
rect 511026 46294 511094 46350
rect 511150 46294 511218 46350
rect 511274 46294 511342 46350
rect 511398 46294 511494 46350
rect 510874 46226 511494 46294
rect 510874 46170 510970 46226
rect 511026 46170 511094 46226
rect 511150 46170 511218 46226
rect 511274 46170 511342 46226
rect 511398 46170 511494 46226
rect 510874 46102 511494 46170
rect 510874 46046 510970 46102
rect 511026 46046 511094 46102
rect 511150 46046 511218 46102
rect 511274 46046 511342 46102
rect 511398 46046 511494 46102
rect 510874 45978 511494 46046
rect 510874 45922 510970 45978
rect 511026 45922 511094 45978
rect 511150 45922 511218 45978
rect 511274 45922 511342 45978
rect 511398 45922 511494 45978
rect 510874 28350 511494 45922
rect 510874 28294 510970 28350
rect 511026 28294 511094 28350
rect 511150 28294 511218 28350
rect 511274 28294 511342 28350
rect 511398 28294 511494 28350
rect 510874 28226 511494 28294
rect 510874 28170 510970 28226
rect 511026 28170 511094 28226
rect 511150 28170 511218 28226
rect 511274 28170 511342 28226
rect 511398 28170 511494 28226
rect 510874 28102 511494 28170
rect 510874 28046 510970 28102
rect 511026 28046 511094 28102
rect 511150 28046 511218 28102
rect 511274 28046 511342 28102
rect 511398 28046 511494 28102
rect 510874 27978 511494 28046
rect 510874 27922 510970 27978
rect 511026 27922 511094 27978
rect 511150 27922 511218 27978
rect 511274 27922 511342 27978
rect 511398 27922 511494 27978
rect 510874 10350 511494 27922
rect 510874 10294 510970 10350
rect 511026 10294 511094 10350
rect 511150 10294 511218 10350
rect 511274 10294 511342 10350
rect 511398 10294 511494 10350
rect 510874 10226 511494 10294
rect 510874 10170 510970 10226
rect 511026 10170 511094 10226
rect 511150 10170 511218 10226
rect 511274 10170 511342 10226
rect 511398 10170 511494 10226
rect 510874 10102 511494 10170
rect 510874 10046 510970 10102
rect 511026 10046 511094 10102
rect 511150 10046 511218 10102
rect 511274 10046 511342 10102
rect 511398 10046 511494 10102
rect 510874 9978 511494 10046
rect 510874 9922 510970 9978
rect 511026 9922 511094 9978
rect 511150 9922 511218 9978
rect 511274 9922 511342 9978
rect 511398 9922 511494 9978
rect 510874 -1120 511494 9922
rect 510874 -1176 510970 -1120
rect 511026 -1176 511094 -1120
rect 511150 -1176 511218 -1120
rect 511274 -1176 511342 -1120
rect 511398 -1176 511494 -1120
rect 510874 -1244 511494 -1176
rect 510874 -1300 510970 -1244
rect 511026 -1300 511094 -1244
rect 511150 -1300 511218 -1244
rect 511274 -1300 511342 -1244
rect 511398 -1300 511494 -1244
rect 510874 -1368 511494 -1300
rect 510874 -1424 510970 -1368
rect 511026 -1424 511094 -1368
rect 511150 -1424 511218 -1368
rect 511274 -1424 511342 -1368
rect 511398 -1424 511494 -1368
rect 510874 -1492 511494 -1424
rect 510874 -1548 510970 -1492
rect 511026 -1548 511094 -1492
rect 511150 -1548 511218 -1492
rect 511274 -1548 511342 -1492
rect 511398 -1548 511494 -1492
rect 510874 -1644 511494 -1548
rect 525154 58350 525774 75922
rect 525154 58294 525250 58350
rect 525306 58294 525374 58350
rect 525430 58294 525498 58350
rect 525554 58294 525622 58350
rect 525678 58294 525774 58350
rect 525154 58226 525774 58294
rect 525154 58170 525250 58226
rect 525306 58170 525374 58226
rect 525430 58170 525498 58226
rect 525554 58170 525622 58226
rect 525678 58170 525774 58226
rect 525154 58102 525774 58170
rect 525154 58046 525250 58102
rect 525306 58046 525374 58102
rect 525430 58046 525498 58102
rect 525554 58046 525622 58102
rect 525678 58046 525774 58102
rect 525154 57978 525774 58046
rect 525154 57922 525250 57978
rect 525306 57922 525374 57978
rect 525430 57922 525498 57978
rect 525554 57922 525622 57978
rect 525678 57922 525774 57978
rect 525154 40350 525774 57922
rect 525154 40294 525250 40350
rect 525306 40294 525374 40350
rect 525430 40294 525498 40350
rect 525554 40294 525622 40350
rect 525678 40294 525774 40350
rect 525154 40226 525774 40294
rect 525154 40170 525250 40226
rect 525306 40170 525374 40226
rect 525430 40170 525498 40226
rect 525554 40170 525622 40226
rect 525678 40170 525774 40226
rect 525154 40102 525774 40170
rect 525154 40046 525250 40102
rect 525306 40046 525374 40102
rect 525430 40046 525498 40102
rect 525554 40046 525622 40102
rect 525678 40046 525774 40102
rect 525154 39978 525774 40046
rect 525154 39922 525250 39978
rect 525306 39922 525374 39978
rect 525430 39922 525498 39978
rect 525554 39922 525622 39978
rect 525678 39922 525774 39978
rect 525154 22350 525774 39922
rect 525154 22294 525250 22350
rect 525306 22294 525374 22350
rect 525430 22294 525498 22350
rect 525554 22294 525622 22350
rect 525678 22294 525774 22350
rect 525154 22226 525774 22294
rect 525154 22170 525250 22226
rect 525306 22170 525374 22226
rect 525430 22170 525498 22226
rect 525554 22170 525622 22226
rect 525678 22170 525774 22226
rect 525154 22102 525774 22170
rect 525154 22046 525250 22102
rect 525306 22046 525374 22102
rect 525430 22046 525498 22102
rect 525554 22046 525622 22102
rect 525678 22046 525774 22102
rect 525154 21978 525774 22046
rect 525154 21922 525250 21978
rect 525306 21922 525374 21978
rect 525430 21922 525498 21978
rect 525554 21922 525622 21978
rect 525678 21922 525774 21978
rect 525154 4350 525774 21922
rect 525154 4294 525250 4350
rect 525306 4294 525374 4350
rect 525430 4294 525498 4350
rect 525554 4294 525622 4350
rect 525678 4294 525774 4350
rect 525154 4226 525774 4294
rect 525154 4170 525250 4226
rect 525306 4170 525374 4226
rect 525430 4170 525498 4226
rect 525554 4170 525622 4226
rect 525678 4170 525774 4226
rect 525154 4102 525774 4170
rect 528332 155204 528388 155214
rect 528332 4228 528388 155148
rect 528332 4162 528388 4172
rect 528874 154350 529494 158858
rect 528874 154294 528970 154350
rect 529026 154294 529094 154350
rect 529150 154294 529218 154350
rect 529274 154294 529342 154350
rect 529398 154294 529494 154350
rect 528874 154226 529494 154294
rect 528874 154170 528970 154226
rect 529026 154170 529094 154226
rect 529150 154170 529218 154226
rect 529274 154170 529342 154226
rect 529398 154170 529494 154226
rect 528874 154102 529494 154170
rect 528874 154046 528970 154102
rect 529026 154046 529094 154102
rect 529150 154046 529218 154102
rect 529274 154046 529342 154102
rect 529398 154046 529494 154102
rect 528874 153978 529494 154046
rect 528874 153922 528970 153978
rect 529026 153922 529094 153978
rect 529150 153922 529218 153978
rect 529274 153922 529342 153978
rect 529398 153922 529494 153978
rect 528874 136350 529494 153922
rect 528874 136294 528970 136350
rect 529026 136294 529094 136350
rect 529150 136294 529218 136350
rect 529274 136294 529342 136350
rect 529398 136294 529494 136350
rect 528874 136226 529494 136294
rect 528874 136170 528970 136226
rect 529026 136170 529094 136226
rect 529150 136170 529218 136226
rect 529274 136170 529342 136226
rect 529398 136170 529494 136226
rect 528874 136102 529494 136170
rect 528874 136046 528970 136102
rect 529026 136046 529094 136102
rect 529150 136046 529218 136102
rect 529274 136046 529342 136102
rect 529398 136046 529494 136102
rect 528874 135978 529494 136046
rect 528874 135922 528970 135978
rect 529026 135922 529094 135978
rect 529150 135922 529218 135978
rect 529274 135922 529342 135978
rect 529398 135922 529494 135978
rect 528874 118350 529494 135922
rect 528874 118294 528970 118350
rect 529026 118294 529094 118350
rect 529150 118294 529218 118350
rect 529274 118294 529342 118350
rect 529398 118294 529494 118350
rect 528874 118226 529494 118294
rect 528874 118170 528970 118226
rect 529026 118170 529094 118226
rect 529150 118170 529218 118226
rect 529274 118170 529342 118226
rect 529398 118170 529494 118226
rect 528874 118102 529494 118170
rect 528874 118046 528970 118102
rect 529026 118046 529094 118102
rect 529150 118046 529218 118102
rect 529274 118046 529342 118102
rect 529398 118046 529494 118102
rect 528874 117978 529494 118046
rect 528874 117922 528970 117978
rect 529026 117922 529094 117978
rect 529150 117922 529218 117978
rect 529274 117922 529342 117978
rect 529398 117922 529494 117978
rect 528874 100350 529494 117922
rect 543154 148350 543774 158858
rect 543154 148294 543250 148350
rect 543306 148294 543374 148350
rect 543430 148294 543498 148350
rect 543554 148294 543622 148350
rect 543678 148294 543774 148350
rect 543154 148226 543774 148294
rect 543154 148170 543250 148226
rect 543306 148170 543374 148226
rect 543430 148170 543498 148226
rect 543554 148170 543622 148226
rect 543678 148170 543774 148226
rect 543154 148102 543774 148170
rect 543154 148046 543250 148102
rect 543306 148046 543374 148102
rect 543430 148046 543498 148102
rect 543554 148046 543622 148102
rect 543678 148046 543774 148102
rect 543154 147978 543774 148046
rect 543154 147922 543250 147978
rect 543306 147922 543374 147978
rect 543430 147922 543498 147978
rect 543554 147922 543622 147978
rect 543678 147922 543774 147978
rect 543154 130350 543774 147922
rect 543154 130294 543250 130350
rect 543306 130294 543374 130350
rect 543430 130294 543498 130350
rect 543554 130294 543622 130350
rect 543678 130294 543774 130350
rect 543154 130226 543774 130294
rect 543154 130170 543250 130226
rect 543306 130170 543374 130226
rect 543430 130170 543498 130226
rect 543554 130170 543622 130226
rect 543678 130170 543774 130226
rect 543154 130102 543774 130170
rect 543154 130046 543250 130102
rect 543306 130046 543374 130102
rect 543430 130046 543498 130102
rect 543554 130046 543622 130102
rect 543678 130046 543774 130102
rect 543154 129978 543774 130046
rect 543154 129922 543250 129978
rect 543306 129922 543374 129978
rect 543430 129922 543498 129978
rect 543554 129922 543622 129978
rect 543678 129922 543774 129978
rect 543154 112350 543774 129922
rect 543154 112294 543250 112350
rect 543306 112294 543374 112350
rect 543430 112294 543498 112350
rect 543554 112294 543622 112350
rect 543678 112294 543774 112350
rect 543154 112226 543774 112294
rect 543154 112170 543250 112226
rect 543306 112170 543374 112226
rect 543430 112170 543498 112226
rect 543554 112170 543622 112226
rect 543678 112170 543774 112226
rect 543154 112102 543774 112170
rect 543154 112046 543250 112102
rect 543306 112046 543374 112102
rect 543430 112046 543498 112102
rect 543554 112046 543622 112102
rect 543678 112046 543774 112102
rect 543154 111978 543774 112046
rect 543154 111922 543250 111978
rect 543306 111922 543374 111978
rect 543430 111922 543498 111978
rect 543554 111922 543622 111978
rect 543678 111922 543774 111978
rect 528874 100294 528970 100350
rect 529026 100294 529094 100350
rect 529150 100294 529218 100350
rect 529274 100294 529342 100350
rect 529398 100294 529494 100350
rect 528874 100226 529494 100294
rect 528874 100170 528970 100226
rect 529026 100170 529094 100226
rect 529150 100170 529218 100226
rect 529274 100170 529342 100226
rect 529398 100170 529494 100226
rect 528874 100102 529494 100170
rect 528874 100046 528970 100102
rect 529026 100046 529094 100102
rect 529150 100046 529218 100102
rect 529274 100046 529342 100102
rect 529398 100046 529494 100102
rect 528874 99978 529494 100046
rect 528874 99922 528970 99978
rect 529026 99922 529094 99978
rect 529150 99922 529218 99978
rect 529274 99922 529342 99978
rect 529398 99922 529494 99978
rect 528874 82350 529494 99922
rect 539808 100350 540128 100384
rect 539808 100294 539878 100350
rect 539934 100294 540002 100350
rect 540058 100294 540128 100350
rect 539808 100226 540128 100294
rect 539808 100170 539878 100226
rect 539934 100170 540002 100226
rect 540058 100170 540128 100226
rect 539808 100102 540128 100170
rect 539808 100046 539878 100102
rect 539934 100046 540002 100102
rect 540058 100046 540128 100102
rect 539808 99978 540128 100046
rect 539808 99922 539878 99978
rect 539934 99922 540002 99978
rect 540058 99922 540128 99978
rect 539808 99888 540128 99922
rect 543154 94350 543774 111922
rect 543154 94294 543250 94350
rect 543306 94294 543374 94350
rect 543430 94294 543498 94350
rect 543554 94294 543622 94350
rect 543678 94294 543774 94350
rect 543154 94226 543774 94294
rect 543154 94170 543250 94226
rect 543306 94170 543374 94226
rect 543430 94170 543498 94226
rect 543554 94170 543622 94226
rect 543678 94170 543774 94226
rect 543154 94102 543774 94170
rect 543154 94046 543250 94102
rect 543306 94046 543374 94102
rect 543430 94046 543498 94102
rect 543554 94046 543622 94102
rect 543678 94046 543774 94102
rect 543154 93978 543774 94046
rect 543154 93922 543250 93978
rect 543306 93922 543374 93978
rect 543430 93922 543498 93978
rect 543554 93922 543622 93978
rect 543678 93922 543774 93978
rect 528874 82294 528970 82350
rect 529026 82294 529094 82350
rect 529150 82294 529218 82350
rect 529274 82294 529342 82350
rect 529398 82294 529494 82350
rect 528874 82226 529494 82294
rect 528874 82170 528970 82226
rect 529026 82170 529094 82226
rect 529150 82170 529218 82226
rect 529274 82170 529342 82226
rect 529398 82170 529494 82226
rect 528874 82102 529494 82170
rect 528874 82046 528970 82102
rect 529026 82046 529094 82102
rect 529150 82046 529218 82102
rect 529274 82046 529342 82102
rect 529398 82046 529494 82102
rect 528874 81978 529494 82046
rect 528874 81922 528970 81978
rect 529026 81922 529094 81978
rect 529150 81922 529218 81978
rect 529274 81922 529342 81978
rect 529398 81922 529494 81978
rect 528874 64350 529494 81922
rect 539808 82350 540128 82384
rect 539808 82294 539878 82350
rect 539934 82294 540002 82350
rect 540058 82294 540128 82350
rect 539808 82226 540128 82294
rect 539808 82170 539878 82226
rect 539934 82170 540002 82226
rect 540058 82170 540128 82226
rect 539808 82102 540128 82170
rect 539808 82046 539878 82102
rect 539934 82046 540002 82102
rect 540058 82046 540128 82102
rect 539808 81978 540128 82046
rect 539808 81922 539878 81978
rect 539934 81922 540002 81978
rect 540058 81922 540128 81978
rect 539808 81888 540128 81922
rect 543154 76350 543774 93922
rect 543154 76294 543250 76350
rect 543306 76294 543374 76350
rect 543430 76294 543498 76350
rect 543554 76294 543622 76350
rect 543678 76294 543774 76350
rect 543154 76226 543774 76294
rect 543154 76170 543250 76226
rect 543306 76170 543374 76226
rect 543430 76170 543498 76226
rect 543554 76170 543622 76226
rect 543678 76170 543774 76226
rect 543154 76102 543774 76170
rect 543154 76046 543250 76102
rect 543306 76046 543374 76102
rect 543430 76046 543498 76102
rect 543554 76046 543622 76102
rect 543678 76046 543774 76102
rect 543154 75978 543774 76046
rect 543154 75922 543250 75978
rect 543306 75922 543374 75978
rect 543430 75922 543498 75978
rect 543554 75922 543622 75978
rect 543678 75922 543774 75978
rect 528874 64294 528970 64350
rect 529026 64294 529094 64350
rect 529150 64294 529218 64350
rect 529274 64294 529342 64350
rect 529398 64294 529494 64350
rect 528874 64226 529494 64294
rect 528874 64170 528970 64226
rect 529026 64170 529094 64226
rect 529150 64170 529218 64226
rect 529274 64170 529342 64226
rect 529398 64170 529494 64226
rect 528874 64102 529494 64170
rect 528874 64046 528970 64102
rect 529026 64046 529094 64102
rect 529150 64046 529218 64102
rect 529274 64046 529342 64102
rect 529398 64046 529494 64102
rect 528874 63978 529494 64046
rect 528874 63922 528970 63978
rect 529026 63922 529094 63978
rect 529150 63922 529218 63978
rect 529274 63922 529342 63978
rect 529398 63922 529494 63978
rect 528874 46350 529494 63922
rect 539808 64350 540128 64384
rect 539808 64294 539878 64350
rect 539934 64294 540002 64350
rect 540058 64294 540128 64350
rect 539808 64226 540128 64294
rect 539808 64170 539878 64226
rect 539934 64170 540002 64226
rect 540058 64170 540128 64226
rect 539808 64102 540128 64170
rect 539808 64046 539878 64102
rect 539934 64046 540002 64102
rect 540058 64046 540128 64102
rect 539808 63978 540128 64046
rect 539808 63922 539878 63978
rect 539934 63922 540002 63978
rect 540058 63922 540128 63978
rect 539808 63888 540128 63922
rect 528874 46294 528970 46350
rect 529026 46294 529094 46350
rect 529150 46294 529218 46350
rect 529274 46294 529342 46350
rect 529398 46294 529494 46350
rect 528874 46226 529494 46294
rect 528874 46170 528970 46226
rect 529026 46170 529094 46226
rect 529150 46170 529218 46226
rect 529274 46170 529342 46226
rect 529398 46170 529494 46226
rect 528874 46102 529494 46170
rect 528874 46046 528970 46102
rect 529026 46046 529094 46102
rect 529150 46046 529218 46102
rect 529274 46046 529342 46102
rect 529398 46046 529494 46102
rect 528874 45978 529494 46046
rect 528874 45922 528970 45978
rect 529026 45922 529094 45978
rect 529150 45922 529218 45978
rect 529274 45922 529342 45978
rect 529398 45922 529494 45978
rect 528874 28350 529494 45922
rect 528874 28294 528970 28350
rect 529026 28294 529094 28350
rect 529150 28294 529218 28350
rect 529274 28294 529342 28350
rect 529398 28294 529494 28350
rect 528874 28226 529494 28294
rect 528874 28170 528970 28226
rect 529026 28170 529094 28226
rect 529150 28170 529218 28226
rect 529274 28170 529342 28226
rect 529398 28170 529494 28226
rect 528874 28102 529494 28170
rect 528874 28046 528970 28102
rect 529026 28046 529094 28102
rect 529150 28046 529218 28102
rect 529274 28046 529342 28102
rect 529398 28046 529494 28102
rect 528874 27978 529494 28046
rect 528874 27922 528970 27978
rect 529026 27922 529094 27978
rect 529150 27922 529218 27978
rect 529274 27922 529342 27978
rect 529398 27922 529494 27978
rect 528874 10350 529494 27922
rect 528874 10294 528970 10350
rect 529026 10294 529094 10350
rect 529150 10294 529218 10350
rect 529274 10294 529342 10350
rect 529398 10294 529494 10350
rect 528874 10226 529494 10294
rect 528874 10170 528970 10226
rect 529026 10170 529094 10226
rect 529150 10170 529218 10226
rect 529274 10170 529342 10226
rect 529398 10170 529494 10226
rect 528874 10102 529494 10170
rect 528874 10046 528970 10102
rect 529026 10046 529094 10102
rect 529150 10046 529218 10102
rect 529274 10046 529342 10102
rect 529398 10046 529494 10102
rect 528874 9978 529494 10046
rect 528874 9922 528970 9978
rect 529026 9922 529094 9978
rect 529150 9922 529218 9978
rect 529274 9922 529342 9978
rect 529398 9922 529494 9978
rect 525154 4046 525250 4102
rect 525306 4046 525374 4102
rect 525430 4046 525498 4102
rect 525554 4046 525622 4102
rect 525678 4046 525774 4102
rect 525154 3978 525774 4046
rect 525154 3922 525250 3978
rect 525306 3922 525374 3978
rect 525430 3922 525498 3978
rect 525554 3922 525622 3978
rect 525678 3922 525774 3978
rect 525154 -160 525774 3922
rect 525154 -216 525250 -160
rect 525306 -216 525374 -160
rect 525430 -216 525498 -160
rect 525554 -216 525622 -160
rect 525678 -216 525774 -160
rect 525154 -284 525774 -216
rect 525154 -340 525250 -284
rect 525306 -340 525374 -284
rect 525430 -340 525498 -284
rect 525554 -340 525622 -284
rect 525678 -340 525774 -284
rect 525154 -408 525774 -340
rect 525154 -464 525250 -408
rect 525306 -464 525374 -408
rect 525430 -464 525498 -408
rect 525554 -464 525622 -408
rect 525678 -464 525774 -408
rect 525154 -532 525774 -464
rect 525154 -588 525250 -532
rect 525306 -588 525374 -532
rect 525430 -588 525498 -532
rect 525554 -588 525622 -532
rect 525678 -588 525774 -532
rect 525154 -1644 525774 -588
rect 528874 -1120 529494 9922
rect 528874 -1176 528970 -1120
rect 529026 -1176 529094 -1120
rect 529150 -1176 529218 -1120
rect 529274 -1176 529342 -1120
rect 529398 -1176 529494 -1120
rect 528874 -1244 529494 -1176
rect 528874 -1300 528970 -1244
rect 529026 -1300 529094 -1244
rect 529150 -1300 529218 -1244
rect 529274 -1300 529342 -1244
rect 529398 -1300 529494 -1244
rect 528874 -1368 529494 -1300
rect 528874 -1424 528970 -1368
rect 529026 -1424 529094 -1368
rect 529150 -1424 529218 -1368
rect 529274 -1424 529342 -1368
rect 529398 -1424 529494 -1368
rect 528874 -1492 529494 -1424
rect 528874 -1548 528970 -1492
rect 529026 -1548 529094 -1492
rect 529150 -1548 529218 -1492
rect 529274 -1548 529342 -1492
rect 529398 -1548 529494 -1492
rect 528874 -1644 529494 -1548
rect 543154 58350 543774 75922
rect 543154 58294 543250 58350
rect 543306 58294 543374 58350
rect 543430 58294 543498 58350
rect 543554 58294 543622 58350
rect 543678 58294 543774 58350
rect 543154 58226 543774 58294
rect 543154 58170 543250 58226
rect 543306 58170 543374 58226
rect 543430 58170 543498 58226
rect 543554 58170 543622 58226
rect 543678 58170 543774 58226
rect 543154 58102 543774 58170
rect 543154 58046 543250 58102
rect 543306 58046 543374 58102
rect 543430 58046 543498 58102
rect 543554 58046 543622 58102
rect 543678 58046 543774 58102
rect 543154 57978 543774 58046
rect 543154 57922 543250 57978
rect 543306 57922 543374 57978
rect 543430 57922 543498 57978
rect 543554 57922 543622 57978
rect 543678 57922 543774 57978
rect 543154 40350 543774 57922
rect 543154 40294 543250 40350
rect 543306 40294 543374 40350
rect 543430 40294 543498 40350
rect 543554 40294 543622 40350
rect 543678 40294 543774 40350
rect 543154 40226 543774 40294
rect 543154 40170 543250 40226
rect 543306 40170 543374 40226
rect 543430 40170 543498 40226
rect 543554 40170 543622 40226
rect 543678 40170 543774 40226
rect 543154 40102 543774 40170
rect 543154 40046 543250 40102
rect 543306 40046 543374 40102
rect 543430 40046 543498 40102
rect 543554 40046 543622 40102
rect 543678 40046 543774 40102
rect 543154 39978 543774 40046
rect 543154 39922 543250 39978
rect 543306 39922 543374 39978
rect 543430 39922 543498 39978
rect 543554 39922 543622 39978
rect 543678 39922 543774 39978
rect 543154 22350 543774 39922
rect 543154 22294 543250 22350
rect 543306 22294 543374 22350
rect 543430 22294 543498 22350
rect 543554 22294 543622 22350
rect 543678 22294 543774 22350
rect 543154 22226 543774 22294
rect 543154 22170 543250 22226
rect 543306 22170 543374 22226
rect 543430 22170 543498 22226
rect 543554 22170 543622 22226
rect 543678 22170 543774 22226
rect 543154 22102 543774 22170
rect 543154 22046 543250 22102
rect 543306 22046 543374 22102
rect 543430 22046 543498 22102
rect 543554 22046 543622 22102
rect 543678 22046 543774 22102
rect 543154 21978 543774 22046
rect 543154 21922 543250 21978
rect 543306 21922 543374 21978
rect 543430 21922 543498 21978
rect 543554 21922 543622 21978
rect 543678 21922 543774 21978
rect 543154 4350 543774 21922
rect 543154 4294 543250 4350
rect 543306 4294 543374 4350
rect 543430 4294 543498 4350
rect 543554 4294 543622 4350
rect 543678 4294 543774 4350
rect 543154 4226 543774 4294
rect 543154 4170 543250 4226
rect 543306 4170 543374 4226
rect 543430 4170 543498 4226
rect 543554 4170 543622 4226
rect 543678 4170 543774 4226
rect 543154 4102 543774 4170
rect 543154 4046 543250 4102
rect 543306 4046 543374 4102
rect 543430 4046 543498 4102
rect 543554 4046 543622 4102
rect 543678 4046 543774 4102
rect 543154 3978 543774 4046
rect 543154 3922 543250 3978
rect 543306 3922 543374 3978
rect 543430 3922 543498 3978
rect 543554 3922 543622 3978
rect 543678 3922 543774 3978
rect 543154 -160 543774 3922
rect 543154 -216 543250 -160
rect 543306 -216 543374 -160
rect 543430 -216 543498 -160
rect 543554 -216 543622 -160
rect 543678 -216 543774 -160
rect 543154 -284 543774 -216
rect 543154 -340 543250 -284
rect 543306 -340 543374 -284
rect 543430 -340 543498 -284
rect 543554 -340 543622 -284
rect 543678 -340 543774 -284
rect 543154 -408 543774 -340
rect 543154 -464 543250 -408
rect 543306 -464 543374 -408
rect 543430 -464 543498 -408
rect 543554 -464 543622 -408
rect 543678 -464 543774 -408
rect 543154 -532 543774 -464
rect 543154 -588 543250 -532
rect 543306 -588 543374 -532
rect 543430 -588 543498 -532
rect 543554 -588 543622 -532
rect 543678 -588 543774 -532
rect 543154 -1644 543774 -588
rect 546874 154350 547494 158858
rect 546874 154294 546970 154350
rect 547026 154294 547094 154350
rect 547150 154294 547218 154350
rect 547274 154294 547342 154350
rect 547398 154294 547494 154350
rect 546874 154226 547494 154294
rect 546874 154170 546970 154226
rect 547026 154170 547094 154226
rect 547150 154170 547218 154226
rect 547274 154170 547342 154226
rect 547398 154170 547494 154226
rect 546874 154102 547494 154170
rect 546874 154046 546970 154102
rect 547026 154046 547094 154102
rect 547150 154046 547218 154102
rect 547274 154046 547342 154102
rect 547398 154046 547494 154102
rect 546874 153978 547494 154046
rect 546874 153922 546970 153978
rect 547026 153922 547094 153978
rect 547150 153922 547218 153978
rect 547274 153922 547342 153978
rect 547398 153922 547494 153978
rect 546874 136350 547494 153922
rect 546874 136294 546970 136350
rect 547026 136294 547094 136350
rect 547150 136294 547218 136350
rect 547274 136294 547342 136350
rect 547398 136294 547494 136350
rect 546874 136226 547494 136294
rect 546874 136170 546970 136226
rect 547026 136170 547094 136226
rect 547150 136170 547218 136226
rect 547274 136170 547342 136226
rect 547398 136170 547494 136226
rect 546874 136102 547494 136170
rect 546874 136046 546970 136102
rect 547026 136046 547094 136102
rect 547150 136046 547218 136102
rect 547274 136046 547342 136102
rect 547398 136046 547494 136102
rect 546874 135978 547494 136046
rect 546874 135922 546970 135978
rect 547026 135922 547094 135978
rect 547150 135922 547218 135978
rect 547274 135922 547342 135978
rect 547398 135922 547494 135978
rect 546874 118350 547494 135922
rect 546874 118294 546970 118350
rect 547026 118294 547094 118350
rect 547150 118294 547218 118350
rect 547274 118294 547342 118350
rect 547398 118294 547494 118350
rect 546874 118226 547494 118294
rect 546874 118170 546970 118226
rect 547026 118170 547094 118226
rect 547150 118170 547218 118226
rect 547274 118170 547342 118226
rect 547398 118170 547494 118226
rect 546874 118102 547494 118170
rect 546874 118046 546970 118102
rect 547026 118046 547094 118102
rect 547150 118046 547218 118102
rect 547274 118046 547342 118102
rect 547398 118046 547494 118102
rect 546874 117978 547494 118046
rect 546874 117922 546970 117978
rect 547026 117922 547094 117978
rect 547150 117922 547218 117978
rect 547274 117922 547342 117978
rect 547398 117922 547494 117978
rect 546874 100350 547494 117922
rect 546874 100294 546970 100350
rect 547026 100294 547094 100350
rect 547150 100294 547218 100350
rect 547274 100294 547342 100350
rect 547398 100294 547494 100350
rect 546874 100226 547494 100294
rect 546874 100170 546970 100226
rect 547026 100170 547094 100226
rect 547150 100170 547218 100226
rect 547274 100170 547342 100226
rect 547398 100170 547494 100226
rect 546874 100102 547494 100170
rect 546874 100046 546970 100102
rect 547026 100046 547094 100102
rect 547150 100046 547218 100102
rect 547274 100046 547342 100102
rect 547398 100046 547494 100102
rect 546874 99978 547494 100046
rect 546874 99922 546970 99978
rect 547026 99922 547094 99978
rect 547150 99922 547218 99978
rect 547274 99922 547342 99978
rect 547398 99922 547494 99978
rect 546874 82350 547494 99922
rect 546874 82294 546970 82350
rect 547026 82294 547094 82350
rect 547150 82294 547218 82350
rect 547274 82294 547342 82350
rect 547398 82294 547494 82350
rect 546874 82226 547494 82294
rect 546874 82170 546970 82226
rect 547026 82170 547094 82226
rect 547150 82170 547218 82226
rect 547274 82170 547342 82226
rect 547398 82170 547494 82226
rect 546874 82102 547494 82170
rect 546874 82046 546970 82102
rect 547026 82046 547094 82102
rect 547150 82046 547218 82102
rect 547274 82046 547342 82102
rect 547398 82046 547494 82102
rect 546874 81978 547494 82046
rect 546874 81922 546970 81978
rect 547026 81922 547094 81978
rect 547150 81922 547218 81978
rect 547274 81922 547342 81978
rect 547398 81922 547494 81978
rect 546874 64350 547494 81922
rect 546874 64294 546970 64350
rect 547026 64294 547094 64350
rect 547150 64294 547218 64350
rect 547274 64294 547342 64350
rect 547398 64294 547494 64350
rect 546874 64226 547494 64294
rect 546874 64170 546970 64226
rect 547026 64170 547094 64226
rect 547150 64170 547218 64226
rect 547274 64170 547342 64226
rect 547398 64170 547494 64226
rect 546874 64102 547494 64170
rect 546874 64046 546970 64102
rect 547026 64046 547094 64102
rect 547150 64046 547218 64102
rect 547274 64046 547342 64102
rect 547398 64046 547494 64102
rect 546874 63978 547494 64046
rect 546874 63922 546970 63978
rect 547026 63922 547094 63978
rect 547150 63922 547218 63978
rect 547274 63922 547342 63978
rect 547398 63922 547494 63978
rect 546874 46350 547494 63922
rect 546874 46294 546970 46350
rect 547026 46294 547094 46350
rect 547150 46294 547218 46350
rect 547274 46294 547342 46350
rect 547398 46294 547494 46350
rect 546874 46226 547494 46294
rect 546874 46170 546970 46226
rect 547026 46170 547094 46226
rect 547150 46170 547218 46226
rect 547274 46170 547342 46226
rect 547398 46170 547494 46226
rect 546874 46102 547494 46170
rect 546874 46046 546970 46102
rect 547026 46046 547094 46102
rect 547150 46046 547218 46102
rect 547274 46046 547342 46102
rect 547398 46046 547494 46102
rect 546874 45978 547494 46046
rect 546874 45922 546970 45978
rect 547026 45922 547094 45978
rect 547150 45922 547218 45978
rect 547274 45922 547342 45978
rect 547398 45922 547494 45978
rect 546874 28350 547494 45922
rect 546874 28294 546970 28350
rect 547026 28294 547094 28350
rect 547150 28294 547218 28350
rect 547274 28294 547342 28350
rect 547398 28294 547494 28350
rect 546874 28226 547494 28294
rect 546874 28170 546970 28226
rect 547026 28170 547094 28226
rect 547150 28170 547218 28226
rect 547274 28170 547342 28226
rect 547398 28170 547494 28226
rect 546874 28102 547494 28170
rect 546874 28046 546970 28102
rect 547026 28046 547094 28102
rect 547150 28046 547218 28102
rect 547274 28046 547342 28102
rect 547398 28046 547494 28102
rect 546874 27978 547494 28046
rect 546874 27922 546970 27978
rect 547026 27922 547094 27978
rect 547150 27922 547218 27978
rect 547274 27922 547342 27978
rect 547398 27922 547494 27978
rect 546874 10350 547494 27922
rect 546874 10294 546970 10350
rect 547026 10294 547094 10350
rect 547150 10294 547218 10350
rect 547274 10294 547342 10350
rect 547398 10294 547494 10350
rect 546874 10226 547494 10294
rect 546874 10170 546970 10226
rect 547026 10170 547094 10226
rect 547150 10170 547218 10226
rect 547274 10170 547342 10226
rect 547398 10170 547494 10226
rect 546874 10102 547494 10170
rect 546874 10046 546970 10102
rect 547026 10046 547094 10102
rect 547150 10046 547218 10102
rect 547274 10046 547342 10102
rect 547398 10046 547494 10102
rect 546874 9978 547494 10046
rect 546874 9922 546970 9978
rect 547026 9922 547094 9978
rect 547150 9922 547218 9978
rect 547274 9922 547342 9978
rect 547398 9922 547494 9978
rect 546874 -1120 547494 9922
rect 551068 156324 551124 156334
rect 551068 3220 551124 156268
rect 561154 148350 561774 158858
rect 561154 148294 561250 148350
rect 561306 148294 561374 148350
rect 561430 148294 561498 148350
rect 561554 148294 561622 148350
rect 561678 148294 561774 148350
rect 561154 148226 561774 148294
rect 561154 148170 561250 148226
rect 561306 148170 561374 148226
rect 561430 148170 561498 148226
rect 561554 148170 561622 148226
rect 561678 148170 561774 148226
rect 561154 148102 561774 148170
rect 561154 148046 561250 148102
rect 561306 148046 561374 148102
rect 561430 148046 561498 148102
rect 561554 148046 561622 148102
rect 561678 148046 561774 148102
rect 561154 147978 561774 148046
rect 561154 147922 561250 147978
rect 561306 147922 561374 147978
rect 561430 147922 561498 147978
rect 561554 147922 561622 147978
rect 561678 147922 561774 147978
rect 561154 130350 561774 147922
rect 561154 130294 561250 130350
rect 561306 130294 561374 130350
rect 561430 130294 561498 130350
rect 561554 130294 561622 130350
rect 561678 130294 561774 130350
rect 561154 130226 561774 130294
rect 561154 130170 561250 130226
rect 561306 130170 561374 130226
rect 561430 130170 561498 130226
rect 561554 130170 561622 130226
rect 561678 130170 561774 130226
rect 561154 130102 561774 130170
rect 561154 130046 561250 130102
rect 561306 130046 561374 130102
rect 561430 130046 561498 130102
rect 561554 130046 561622 130102
rect 561678 130046 561774 130102
rect 561154 129978 561774 130046
rect 561154 129922 561250 129978
rect 561306 129922 561374 129978
rect 561430 129922 561498 129978
rect 561554 129922 561622 129978
rect 561678 129922 561774 129978
rect 561154 112350 561774 129922
rect 561154 112294 561250 112350
rect 561306 112294 561374 112350
rect 561430 112294 561498 112350
rect 561554 112294 561622 112350
rect 561678 112294 561774 112350
rect 561154 112226 561774 112294
rect 561154 112170 561250 112226
rect 561306 112170 561374 112226
rect 561430 112170 561498 112226
rect 561554 112170 561622 112226
rect 561678 112170 561774 112226
rect 561154 112102 561774 112170
rect 561154 112046 561250 112102
rect 561306 112046 561374 112102
rect 561430 112046 561498 112102
rect 561554 112046 561622 112102
rect 561678 112046 561774 112102
rect 561154 111978 561774 112046
rect 561154 111922 561250 111978
rect 561306 111922 561374 111978
rect 561430 111922 561498 111978
rect 561554 111922 561622 111978
rect 561678 111922 561774 111978
rect 555168 94350 555488 94384
rect 555168 94294 555238 94350
rect 555294 94294 555362 94350
rect 555418 94294 555488 94350
rect 555168 94226 555488 94294
rect 555168 94170 555238 94226
rect 555294 94170 555362 94226
rect 555418 94170 555488 94226
rect 555168 94102 555488 94170
rect 555168 94046 555238 94102
rect 555294 94046 555362 94102
rect 555418 94046 555488 94102
rect 555168 93978 555488 94046
rect 555168 93922 555238 93978
rect 555294 93922 555362 93978
rect 555418 93922 555488 93978
rect 555168 93888 555488 93922
rect 561154 94350 561774 111922
rect 561154 94294 561250 94350
rect 561306 94294 561374 94350
rect 561430 94294 561498 94350
rect 561554 94294 561622 94350
rect 561678 94294 561774 94350
rect 561154 94226 561774 94294
rect 561154 94170 561250 94226
rect 561306 94170 561374 94226
rect 561430 94170 561498 94226
rect 561554 94170 561622 94226
rect 561678 94170 561774 94226
rect 561154 94102 561774 94170
rect 561154 94046 561250 94102
rect 561306 94046 561374 94102
rect 561430 94046 561498 94102
rect 561554 94046 561622 94102
rect 561678 94046 561774 94102
rect 561154 93978 561774 94046
rect 561154 93922 561250 93978
rect 561306 93922 561374 93978
rect 561430 93922 561498 93978
rect 561554 93922 561622 93978
rect 561678 93922 561774 93978
rect 555168 76350 555488 76384
rect 555168 76294 555238 76350
rect 555294 76294 555362 76350
rect 555418 76294 555488 76350
rect 555168 76226 555488 76294
rect 555168 76170 555238 76226
rect 555294 76170 555362 76226
rect 555418 76170 555488 76226
rect 555168 76102 555488 76170
rect 555168 76046 555238 76102
rect 555294 76046 555362 76102
rect 555418 76046 555488 76102
rect 555168 75978 555488 76046
rect 555168 75922 555238 75978
rect 555294 75922 555362 75978
rect 555418 75922 555488 75978
rect 555168 75888 555488 75922
rect 561154 76350 561774 93922
rect 561154 76294 561250 76350
rect 561306 76294 561374 76350
rect 561430 76294 561498 76350
rect 561554 76294 561622 76350
rect 561678 76294 561774 76350
rect 561154 76226 561774 76294
rect 561154 76170 561250 76226
rect 561306 76170 561374 76226
rect 561430 76170 561498 76226
rect 561554 76170 561622 76226
rect 561678 76170 561774 76226
rect 561154 76102 561774 76170
rect 561154 76046 561250 76102
rect 561306 76046 561374 76102
rect 561430 76046 561498 76102
rect 561554 76046 561622 76102
rect 561678 76046 561774 76102
rect 561154 75978 561774 76046
rect 561154 75922 561250 75978
rect 561306 75922 561374 75978
rect 561430 75922 561498 75978
rect 561554 75922 561622 75978
rect 561678 75922 561774 75978
rect 551068 3154 551124 3164
rect 561154 58350 561774 75922
rect 561154 58294 561250 58350
rect 561306 58294 561374 58350
rect 561430 58294 561498 58350
rect 561554 58294 561622 58350
rect 561678 58294 561774 58350
rect 561154 58226 561774 58294
rect 561154 58170 561250 58226
rect 561306 58170 561374 58226
rect 561430 58170 561498 58226
rect 561554 58170 561622 58226
rect 561678 58170 561774 58226
rect 561154 58102 561774 58170
rect 561154 58046 561250 58102
rect 561306 58046 561374 58102
rect 561430 58046 561498 58102
rect 561554 58046 561622 58102
rect 561678 58046 561774 58102
rect 561154 57978 561774 58046
rect 561154 57922 561250 57978
rect 561306 57922 561374 57978
rect 561430 57922 561498 57978
rect 561554 57922 561622 57978
rect 561678 57922 561774 57978
rect 561154 40350 561774 57922
rect 561154 40294 561250 40350
rect 561306 40294 561374 40350
rect 561430 40294 561498 40350
rect 561554 40294 561622 40350
rect 561678 40294 561774 40350
rect 561154 40226 561774 40294
rect 561154 40170 561250 40226
rect 561306 40170 561374 40226
rect 561430 40170 561498 40226
rect 561554 40170 561622 40226
rect 561678 40170 561774 40226
rect 561154 40102 561774 40170
rect 561154 40046 561250 40102
rect 561306 40046 561374 40102
rect 561430 40046 561498 40102
rect 561554 40046 561622 40102
rect 561678 40046 561774 40102
rect 561154 39978 561774 40046
rect 561154 39922 561250 39978
rect 561306 39922 561374 39978
rect 561430 39922 561498 39978
rect 561554 39922 561622 39978
rect 561678 39922 561774 39978
rect 561154 22350 561774 39922
rect 561154 22294 561250 22350
rect 561306 22294 561374 22350
rect 561430 22294 561498 22350
rect 561554 22294 561622 22350
rect 561678 22294 561774 22350
rect 561154 22226 561774 22294
rect 561154 22170 561250 22226
rect 561306 22170 561374 22226
rect 561430 22170 561498 22226
rect 561554 22170 561622 22226
rect 561678 22170 561774 22226
rect 561154 22102 561774 22170
rect 561154 22046 561250 22102
rect 561306 22046 561374 22102
rect 561430 22046 561498 22102
rect 561554 22046 561622 22102
rect 561678 22046 561774 22102
rect 561154 21978 561774 22046
rect 561154 21922 561250 21978
rect 561306 21922 561374 21978
rect 561430 21922 561498 21978
rect 561554 21922 561622 21978
rect 561678 21922 561774 21978
rect 561154 4350 561774 21922
rect 561154 4294 561250 4350
rect 561306 4294 561374 4350
rect 561430 4294 561498 4350
rect 561554 4294 561622 4350
rect 561678 4294 561774 4350
rect 561154 4226 561774 4294
rect 561154 4170 561250 4226
rect 561306 4170 561374 4226
rect 561430 4170 561498 4226
rect 561554 4170 561622 4226
rect 561678 4170 561774 4226
rect 561154 4102 561774 4170
rect 561154 4046 561250 4102
rect 561306 4046 561374 4102
rect 561430 4046 561498 4102
rect 561554 4046 561622 4102
rect 561678 4046 561774 4102
rect 561154 3978 561774 4046
rect 561154 3922 561250 3978
rect 561306 3922 561374 3978
rect 561430 3922 561498 3978
rect 561554 3922 561622 3978
rect 561678 3922 561774 3978
rect 546874 -1176 546970 -1120
rect 547026 -1176 547094 -1120
rect 547150 -1176 547218 -1120
rect 547274 -1176 547342 -1120
rect 547398 -1176 547494 -1120
rect 546874 -1244 547494 -1176
rect 546874 -1300 546970 -1244
rect 547026 -1300 547094 -1244
rect 547150 -1300 547218 -1244
rect 547274 -1300 547342 -1244
rect 547398 -1300 547494 -1244
rect 546874 -1368 547494 -1300
rect 546874 -1424 546970 -1368
rect 547026 -1424 547094 -1368
rect 547150 -1424 547218 -1368
rect 547274 -1424 547342 -1368
rect 547398 -1424 547494 -1368
rect 546874 -1492 547494 -1424
rect 546874 -1548 546970 -1492
rect 547026 -1548 547094 -1492
rect 547150 -1548 547218 -1492
rect 547274 -1548 547342 -1492
rect 547398 -1548 547494 -1492
rect 546874 -1644 547494 -1548
rect 561154 -160 561774 3922
rect 563612 156324 563668 156334
rect 563612 756 563668 156268
rect 563612 690 563668 700
rect 564874 154350 565494 158858
rect 564874 154294 564970 154350
rect 565026 154294 565094 154350
rect 565150 154294 565218 154350
rect 565274 154294 565342 154350
rect 565398 154294 565494 154350
rect 564874 154226 565494 154294
rect 564874 154170 564970 154226
rect 565026 154170 565094 154226
rect 565150 154170 565218 154226
rect 565274 154170 565342 154226
rect 565398 154170 565494 154226
rect 564874 154102 565494 154170
rect 564874 154046 564970 154102
rect 565026 154046 565094 154102
rect 565150 154046 565218 154102
rect 565274 154046 565342 154102
rect 565398 154046 565494 154102
rect 564874 153978 565494 154046
rect 564874 153922 564970 153978
rect 565026 153922 565094 153978
rect 565150 153922 565218 153978
rect 565274 153922 565342 153978
rect 565398 153922 565494 153978
rect 564874 136350 565494 153922
rect 564874 136294 564970 136350
rect 565026 136294 565094 136350
rect 565150 136294 565218 136350
rect 565274 136294 565342 136350
rect 565398 136294 565494 136350
rect 564874 136226 565494 136294
rect 564874 136170 564970 136226
rect 565026 136170 565094 136226
rect 565150 136170 565218 136226
rect 565274 136170 565342 136226
rect 565398 136170 565494 136226
rect 564874 136102 565494 136170
rect 564874 136046 564970 136102
rect 565026 136046 565094 136102
rect 565150 136046 565218 136102
rect 565274 136046 565342 136102
rect 565398 136046 565494 136102
rect 564874 135978 565494 136046
rect 564874 135922 564970 135978
rect 565026 135922 565094 135978
rect 565150 135922 565218 135978
rect 565274 135922 565342 135978
rect 565398 135922 565494 135978
rect 564874 118350 565494 135922
rect 564874 118294 564970 118350
rect 565026 118294 565094 118350
rect 565150 118294 565218 118350
rect 565274 118294 565342 118350
rect 565398 118294 565494 118350
rect 564874 118226 565494 118294
rect 564874 118170 564970 118226
rect 565026 118170 565094 118226
rect 565150 118170 565218 118226
rect 565274 118170 565342 118226
rect 565398 118170 565494 118226
rect 564874 118102 565494 118170
rect 564874 118046 564970 118102
rect 565026 118046 565094 118102
rect 565150 118046 565218 118102
rect 565274 118046 565342 118102
rect 565398 118046 565494 118102
rect 564874 117978 565494 118046
rect 564874 117922 564970 117978
rect 565026 117922 565094 117978
rect 565150 117922 565218 117978
rect 565274 117922 565342 117978
rect 565398 117922 565494 117978
rect 564874 100350 565494 117922
rect 564874 100294 564970 100350
rect 565026 100294 565094 100350
rect 565150 100294 565218 100350
rect 565274 100294 565342 100350
rect 565398 100294 565494 100350
rect 564874 100226 565494 100294
rect 564874 100170 564970 100226
rect 565026 100170 565094 100226
rect 565150 100170 565218 100226
rect 565274 100170 565342 100226
rect 565398 100170 565494 100226
rect 564874 100102 565494 100170
rect 564874 100046 564970 100102
rect 565026 100046 565094 100102
rect 565150 100046 565218 100102
rect 565274 100046 565342 100102
rect 565398 100046 565494 100102
rect 564874 99978 565494 100046
rect 564874 99922 564970 99978
rect 565026 99922 565094 99978
rect 565150 99922 565218 99978
rect 565274 99922 565342 99978
rect 565398 99922 565494 99978
rect 564874 82350 565494 99922
rect 564874 82294 564970 82350
rect 565026 82294 565094 82350
rect 565150 82294 565218 82350
rect 565274 82294 565342 82350
rect 565398 82294 565494 82350
rect 564874 82226 565494 82294
rect 564874 82170 564970 82226
rect 565026 82170 565094 82226
rect 565150 82170 565218 82226
rect 565274 82170 565342 82226
rect 565398 82170 565494 82226
rect 564874 82102 565494 82170
rect 564874 82046 564970 82102
rect 565026 82046 565094 82102
rect 565150 82046 565218 82102
rect 565274 82046 565342 82102
rect 565398 82046 565494 82102
rect 564874 81978 565494 82046
rect 564874 81922 564970 81978
rect 565026 81922 565094 81978
rect 565150 81922 565218 81978
rect 565274 81922 565342 81978
rect 565398 81922 565494 81978
rect 564874 64350 565494 81922
rect 564874 64294 564970 64350
rect 565026 64294 565094 64350
rect 565150 64294 565218 64350
rect 565274 64294 565342 64350
rect 565398 64294 565494 64350
rect 564874 64226 565494 64294
rect 564874 64170 564970 64226
rect 565026 64170 565094 64226
rect 565150 64170 565218 64226
rect 565274 64170 565342 64226
rect 565398 64170 565494 64226
rect 564874 64102 565494 64170
rect 564874 64046 564970 64102
rect 565026 64046 565094 64102
rect 565150 64046 565218 64102
rect 565274 64046 565342 64102
rect 565398 64046 565494 64102
rect 564874 63978 565494 64046
rect 564874 63922 564970 63978
rect 565026 63922 565094 63978
rect 565150 63922 565218 63978
rect 565274 63922 565342 63978
rect 565398 63922 565494 63978
rect 564874 46350 565494 63922
rect 564874 46294 564970 46350
rect 565026 46294 565094 46350
rect 565150 46294 565218 46350
rect 565274 46294 565342 46350
rect 565398 46294 565494 46350
rect 564874 46226 565494 46294
rect 564874 46170 564970 46226
rect 565026 46170 565094 46226
rect 565150 46170 565218 46226
rect 565274 46170 565342 46226
rect 565398 46170 565494 46226
rect 564874 46102 565494 46170
rect 564874 46046 564970 46102
rect 565026 46046 565094 46102
rect 565150 46046 565218 46102
rect 565274 46046 565342 46102
rect 565398 46046 565494 46102
rect 564874 45978 565494 46046
rect 564874 45922 564970 45978
rect 565026 45922 565094 45978
rect 565150 45922 565218 45978
rect 565274 45922 565342 45978
rect 565398 45922 565494 45978
rect 564874 28350 565494 45922
rect 564874 28294 564970 28350
rect 565026 28294 565094 28350
rect 565150 28294 565218 28350
rect 565274 28294 565342 28350
rect 565398 28294 565494 28350
rect 564874 28226 565494 28294
rect 564874 28170 564970 28226
rect 565026 28170 565094 28226
rect 565150 28170 565218 28226
rect 565274 28170 565342 28226
rect 565398 28170 565494 28226
rect 564874 28102 565494 28170
rect 564874 28046 564970 28102
rect 565026 28046 565094 28102
rect 565150 28046 565218 28102
rect 565274 28046 565342 28102
rect 565398 28046 565494 28102
rect 564874 27978 565494 28046
rect 564874 27922 564970 27978
rect 565026 27922 565094 27978
rect 565150 27922 565218 27978
rect 565274 27922 565342 27978
rect 565398 27922 565494 27978
rect 564874 10350 565494 27922
rect 564874 10294 564970 10350
rect 565026 10294 565094 10350
rect 565150 10294 565218 10350
rect 565274 10294 565342 10350
rect 565398 10294 565494 10350
rect 564874 10226 565494 10294
rect 564874 10170 564970 10226
rect 565026 10170 565094 10226
rect 565150 10170 565218 10226
rect 565274 10170 565342 10226
rect 565398 10170 565494 10226
rect 564874 10102 565494 10170
rect 564874 10046 564970 10102
rect 565026 10046 565094 10102
rect 565150 10046 565218 10102
rect 565274 10046 565342 10102
rect 565398 10046 565494 10102
rect 564874 9978 565494 10046
rect 564874 9922 564970 9978
rect 565026 9922 565094 9978
rect 565150 9922 565218 9978
rect 565274 9922 565342 9978
rect 565398 9922 565494 9978
rect 561154 -216 561250 -160
rect 561306 -216 561374 -160
rect 561430 -216 561498 -160
rect 561554 -216 561622 -160
rect 561678 -216 561774 -160
rect 561154 -284 561774 -216
rect 561154 -340 561250 -284
rect 561306 -340 561374 -284
rect 561430 -340 561498 -284
rect 561554 -340 561622 -284
rect 561678 -340 561774 -284
rect 561154 -408 561774 -340
rect 561154 -464 561250 -408
rect 561306 -464 561374 -408
rect 561430 -464 561498 -408
rect 561554 -464 561622 -408
rect 561678 -464 561774 -408
rect 561154 -532 561774 -464
rect 561154 -588 561250 -532
rect 561306 -588 561374 -532
rect 561430 -588 561498 -532
rect 561554 -588 561622 -532
rect 561678 -588 561774 -532
rect 561154 -1644 561774 -588
rect 564874 -1120 565494 9922
rect 564874 -1176 564970 -1120
rect 565026 -1176 565094 -1120
rect 565150 -1176 565218 -1120
rect 565274 -1176 565342 -1120
rect 565398 -1176 565494 -1120
rect 564874 -1244 565494 -1176
rect 564874 -1300 564970 -1244
rect 565026 -1300 565094 -1244
rect 565150 -1300 565218 -1244
rect 565274 -1300 565342 -1244
rect 565398 -1300 565494 -1244
rect 564874 -1368 565494 -1300
rect 564874 -1424 564970 -1368
rect 565026 -1424 565094 -1368
rect 565150 -1424 565218 -1368
rect 565274 -1424 565342 -1368
rect 565398 -1424 565494 -1368
rect 564874 -1492 565494 -1424
rect 564874 -1548 564970 -1492
rect 565026 -1548 565094 -1492
rect 565150 -1548 565218 -1492
rect 565274 -1548 565342 -1492
rect 565398 -1548 565494 -1492
rect 564874 -1644 565494 -1548
rect 579154 148350 579774 165922
rect 579154 148294 579250 148350
rect 579306 148294 579374 148350
rect 579430 148294 579498 148350
rect 579554 148294 579622 148350
rect 579678 148294 579774 148350
rect 579154 148226 579774 148294
rect 579154 148170 579250 148226
rect 579306 148170 579374 148226
rect 579430 148170 579498 148226
rect 579554 148170 579622 148226
rect 579678 148170 579774 148226
rect 579154 148102 579774 148170
rect 579154 148046 579250 148102
rect 579306 148046 579374 148102
rect 579430 148046 579498 148102
rect 579554 148046 579622 148102
rect 579678 148046 579774 148102
rect 579154 147978 579774 148046
rect 579154 147922 579250 147978
rect 579306 147922 579374 147978
rect 579430 147922 579498 147978
rect 579554 147922 579622 147978
rect 579678 147922 579774 147978
rect 579154 130350 579774 147922
rect 579154 130294 579250 130350
rect 579306 130294 579374 130350
rect 579430 130294 579498 130350
rect 579554 130294 579622 130350
rect 579678 130294 579774 130350
rect 579154 130226 579774 130294
rect 579154 130170 579250 130226
rect 579306 130170 579374 130226
rect 579430 130170 579498 130226
rect 579554 130170 579622 130226
rect 579678 130170 579774 130226
rect 579154 130102 579774 130170
rect 579154 130046 579250 130102
rect 579306 130046 579374 130102
rect 579430 130046 579498 130102
rect 579554 130046 579622 130102
rect 579678 130046 579774 130102
rect 579154 129978 579774 130046
rect 579154 129922 579250 129978
rect 579306 129922 579374 129978
rect 579430 129922 579498 129978
rect 579554 129922 579622 129978
rect 579678 129922 579774 129978
rect 579154 112350 579774 129922
rect 579154 112294 579250 112350
rect 579306 112294 579374 112350
rect 579430 112294 579498 112350
rect 579554 112294 579622 112350
rect 579678 112294 579774 112350
rect 579154 112226 579774 112294
rect 579154 112170 579250 112226
rect 579306 112170 579374 112226
rect 579430 112170 579498 112226
rect 579554 112170 579622 112226
rect 579678 112170 579774 112226
rect 579154 112102 579774 112170
rect 579154 112046 579250 112102
rect 579306 112046 579374 112102
rect 579430 112046 579498 112102
rect 579554 112046 579622 112102
rect 579678 112046 579774 112102
rect 579154 111978 579774 112046
rect 579154 111922 579250 111978
rect 579306 111922 579374 111978
rect 579430 111922 579498 111978
rect 579554 111922 579622 111978
rect 579678 111922 579774 111978
rect 579154 94350 579774 111922
rect 579154 94294 579250 94350
rect 579306 94294 579374 94350
rect 579430 94294 579498 94350
rect 579554 94294 579622 94350
rect 579678 94294 579774 94350
rect 579154 94226 579774 94294
rect 579154 94170 579250 94226
rect 579306 94170 579374 94226
rect 579430 94170 579498 94226
rect 579554 94170 579622 94226
rect 579678 94170 579774 94226
rect 579154 94102 579774 94170
rect 579154 94046 579250 94102
rect 579306 94046 579374 94102
rect 579430 94046 579498 94102
rect 579554 94046 579622 94102
rect 579678 94046 579774 94102
rect 579154 93978 579774 94046
rect 579154 93922 579250 93978
rect 579306 93922 579374 93978
rect 579430 93922 579498 93978
rect 579554 93922 579622 93978
rect 579678 93922 579774 93978
rect 579154 76350 579774 93922
rect 579154 76294 579250 76350
rect 579306 76294 579374 76350
rect 579430 76294 579498 76350
rect 579554 76294 579622 76350
rect 579678 76294 579774 76350
rect 579154 76226 579774 76294
rect 579154 76170 579250 76226
rect 579306 76170 579374 76226
rect 579430 76170 579498 76226
rect 579554 76170 579622 76226
rect 579678 76170 579774 76226
rect 579154 76102 579774 76170
rect 579154 76046 579250 76102
rect 579306 76046 579374 76102
rect 579430 76046 579498 76102
rect 579554 76046 579622 76102
rect 579678 76046 579774 76102
rect 579154 75978 579774 76046
rect 579154 75922 579250 75978
rect 579306 75922 579374 75978
rect 579430 75922 579498 75978
rect 579554 75922 579622 75978
rect 579678 75922 579774 75978
rect 579154 58350 579774 75922
rect 579154 58294 579250 58350
rect 579306 58294 579374 58350
rect 579430 58294 579498 58350
rect 579554 58294 579622 58350
rect 579678 58294 579774 58350
rect 579154 58226 579774 58294
rect 579154 58170 579250 58226
rect 579306 58170 579374 58226
rect 579430 58170 579498 58226
rect 579554 58170 579622 58226
rect 579678 58170 579774 58226
rect 579154 58102 579774 58170
rect 579154 58046 579250 58102
rect 579306 58046 579374 58102
rect 579430 58046 579498 58102
rect 579554 58046 579622 58102
rect 579678 58046 579774 58102
rect 579154 57978 579774 58046
rect 579154 57922 579250 57978
rect 579306 57922 579374 57978
rect 579430 57922 579498 57978
rect 579554 57922 579622 57978
rect 579678 57922 579774 57978
rect 579154 40350 579774 57922
rect 579154 40294 579250 40350
rect 579306 40294 579374 40350
rect 579430 40294 579498 40350
rect 579554 40294 579622 40350
rect 579678 40294 579774 40350
rect 579154 40226 579774 40294
rect 579154 40170 579250 40226
rect 579306 40170 579374 40226
rect 579430 40170 579498 40226
rect 579554 40170 579622 40226
rect 579678 40170 579774 40226
rect 579154 40102 579774 40170
rect 579154 40046 579250 40102
rect 579306 40046 579374 40102
rect 579430 40046 579498 40102
rect 579554 40046 579622 40102
rect 579678 40046 579774 40102
rect 579154 39978 579774 40046
rect 579154 39922 579250 39978
rect 579306 39922 579374 39978
rect 579430 39922 579498 39978
rect 579554 39922 579622 39978
rect 579678 39922 579774 39978
rect 579154 22350 579774 39922
rect 579154 22294 579250 22350
rect 579306 22294 579374 22350
rect 579430 22294 579498 22350
rect 579554 22294 579622 22350
rect 579678 22294 579774 22350
rect 579154 22226 579774 22294
rect 579154 22170 579250 22226
rect 579306 22170 579374 22226
rect 579430 22170 579498 22226
rect 579554 22170 579622 22226
rect 579678 22170 579774 22226
rect 579154 22102 579774 22170
rect 579154 22046 579250 22102
rect 579306 22046 579374 22102
rect 579430 22046 579498 22102
rect 579554 22046 579622 22102
rect 579678 22046 579774 22102
rect 579154 21978 579774 22046
rect 579154 21922 579250 21978
rect 579306 21922 579374 21978
rect 579430 21922 579498 21978
rect 579554 21922 579622 21978
rect 579678 21922 579774 21978
rect 579154 4350 579774 21922
rect 579154 4294 579250 4350
rect 579306 4294 579374 4350
rect 579430 4294 579498 4350
rect 579554 4294 579622 4350
rect 579678 4294 579774 4350
rect 579154 4226 579774 4294
rect 579154 4170 579250 4226
rect 579306 4170 579374 4226
rect 579430 4170 579498 4226
rect 579554 4170 579622 4226
rect 579678 4170 579774 4226
rect 579154 4102 579774 4170
rect 579154 4046 579250 4102
rect 579306 4046 579374 4102
rect 579430 4046 579498 4102
rect 579554 4046 579622 4102
rect 579678 4046 579774 4102
rect 579154 3978 579774 4046
rect 579154 3922 579250 3978
rect 579306 3922 579374 3978
rect 579430 3922 579498 3978
rect 579554 3922 579622 3978
rect 579678 3922 579774 3978
rect 579154 -160 579774 3922
rect 579154 -216 579250 -160
rect 579306 -216 579374 -160
rect 579430 -216 579498 -160
rect 579554 -216 579622 -160
rect 579678 -216 579774 -160
rect 579154 -284 579774 -216
rect 579154 -340 579250 -284
rect 579306 -340 579374 -284
rect 579430 -340 579498 -284
rect 579554 -340 579622 -284
rect 579678 -340 579774 -284
rect 579154 -408 579774 -340
rect 579154 -464 579250 -408
rect 579306 -464 579374 -408
rect 579430 -464 579498 -408
rect 579554 -464 579622 -408
rect 579678 -464 579774 -408
rect 579154 -532 579774 -464
rect 579154 -588 579250 -532
rect 579306 -588 579374 -532
rect 579430 -588 579498 -532
rect 579554 -588 579622 -532
rect 579678 -588 579774 -532
rect 579154 -1644 579774 -588
rect 582874 598172 583494 598268
rect 582874 598116 582970 598172
rect 583026 598116 583094 598172
rect 583150 598116 583218 598172
rect 583274 598116 583342 598172
rect 583398 598116 583494 598172
rect 582874 598048 583494 598116
rect 582874 597992 582970 598048
rect 583026 597992 583094 598048
rect 583150 597992 583218 598048
rect 583274 597992 583342 598048
rect 583398 597992 583494 598048
rect 582874 597924 583494 597992
rect 582874 597868 582970 597924
rect 583026 597868 583094 597924
rect 583150 597868 583218 597924
rect 583274 597868 583342 597924
rect 583398 597868 583494 597924
rect 582874 597800 583494 597868
rect 582874 597744 582970 597800
rect 583026 597744 583094 597800
rect 583150 597744 583218 597800
rect 583274 597744 583342 597800
rect 583398 597744 583494 597800
rect 582874 586350 583494 597744
rect 597360 598172 597980 598268
rect 597360 598116 597456 598172
rect 597512 598116 597580 598172
rect 597636 598116 597704 598172
rect 597760 598116 597828 598172
rect 597884 598116 597980 598172
rect 597360 598048 597980 598116
rect 597360 597992 597456 598048
rect 597512 597992 597580 598048
rect 597636 597992 597704 598048
rect 597760 597992 597828 598048
rect 597884 597992 597980 598048
rect 597360 597924 597980 597992
rect 597360 597868 597456 597924
rect 597512 597868 597580 597924
rect 597636 597868 597704 597924
rect 597760 597868 597828 597924
rect 597884 597868 597980 597924
rect 597360 597800 597980 597868
rect 597360 597744 597456 597800
rect 597512 597744 597580 597800
rect 597636 597744 597704 597800
rect 597760 597744 597828 597800
rect 597884 597744 597980 597800
rect 582874 586294 582970 586350
rect 583026 586294 583094 586350
rect 583150 586294 583218 586350
rect 583274 586294 583342 586350
rect 583398 586294 583494 586350
rect 582874 586226 583494 586294
rect 582874 586170 582970 586226
rect 583026 586170 583094 586226
rect 583150 586170 583218 586226
rect 583274 586170 583342 586226
rect 583398 586170 583494 586226
rect 582874 586102 583494 586170
rect 582874 586046 582970 586102
rect 583026 586046 583094 586102
rect 583150 586046 583218 586102
rect 583274 586046 583342 586102
rect 583398 586046 583494 586102
rect 582874 585978 583494 586046
rect 582874 585922 582970 585978
rect 583026 585922 583094 585978
rect 583150 585922 583218 585978
rect 583274 585922 583342 585978
rect 583398 585922 583494 585978
rect 582874 568350 583494 585922
rect 582874 568294 582970 568350
rect 583026 568294 583094 568350
rect 583150 568294 583218 568350
rect 583274 568294 583342 568350
rect 583398 568294 583494 568350
rect 582874 568226 583494 568294
rect 582874 568170 582970 568226
rect 583026 568170 583094 568226
rect 583150 568170 583218 568226
rect 583274 568170 583342 568226
rect 583398 568170 583494 568226
rect 582874 568102 583494 568170
rect 582874 568046 582970 568102
rect 583026 568046 583094 568102
rect 583150 568046 583218 568102
rect 583274 568046 583342 568102
rect 583398 568046 583494 568102
rect 582874 567978 583494 568046
rect 582874 567922 582970 567978
rect 583026 567922 583094 567978
rect 583150 567922 583218 567978
rect 583274 567922 583342 567978
rect 583398 567922 583494 567978
rect 582874 550350 583494 567922
rect 582874 550294 582970 550350
rect 583026 550294 583094 550350
rect 583150 550294 583218 550350
rect 583274 550294 583342 550350
rect 583398 550294 583494 550350
rect 582874 550226 583494 550294
rect 582874 550170 582970 550226
rect 583026 550170 583094 550226
rect 583150 550170 583218 550226
rect 583274 550170 583342 550226
rect 583398 550170 583494 550226
rect 582874 550102 583494 550170
rect 582874 550046 582970 550102
rect 583026 550046 583094 550102
rect 583150 550046 583218 550102
rect 583274 550046 583342 550102
rect 583398 550046 583494 550102
rect 582874 549978 583494 550046
rect 582874 549922 582970 549978
rect 583026 549922 583094 549978
rect 583150 549922 583218 549978
rect 583274 549922 583342 549978
rect 583398 549922 583494 549978
rect 582874 532350 583494 549922
rect 582874 532294 582970 532350
rect 583026 532294 583094 532350
rect 583150 532294 583218 532350
rect 583274 532294 583342 532350
rect 583398 532294 583494 532350
rect 582874 532226 583494 532294
rect 582874 532170 582970 532226
rect 583026 532170 583094 532226
rect 583150 532170 583218 532226
rect 583274 532170 583342 532226
rect 583398 532170 583494 532226
rect 582874 532102 583494 532170
rect 582874 532046 582970 532102
rect 583026 532046 583094 532102
rect 583150 532046 583218 532102
rect 583274 532046 583342 532102
rect 583398 532046 583494 532102
rect 582874 531978 583494 532046
rect 582874 531922 582970 531978
rect 583026 531922 583094 531978
rect 583150 531922 583218 531978
rect 583274 531922 583342 531978
rect 583398 531922 583494 531978
rect 582874 514350 583494 531922
rect 582874 514294 582970 514350
rect 583026 514294 583094 514350
rect 583150 514294 583218 514350
rect 583274 514294 583342 514350
rect 583398 514294 583494 514350
rect 582874 514226 583494 514294
rect 582874 514170 582970 514226
rect 583026 514170 583094 514226
rect 583150 514170 583218 514226
rect 583274 514170 583342 514226
rect 583398 514170 583494 514226
rect 582874 514102 583494 514170
rect 582874 514046 582970 514102
rect 583026 514046 583094 514102
rect 583150 514046 583218 514102
rect 583274 514046 583342 514102
rect 583398 514046 583494 514102
rect 582874 513978 583494 514046
rect 582874 513922 582970 513978
rect 583026 513922 583094 513978
rect 583150 513922 583218 513978
rect 583274 513922 583342 513978
rect 583398 513922 583494 513978
rect 582874 496350 583494 513922
rect 582874 496294 582970 496350
rect 583026 496294 583094 496350
rect 583150 496294 583218 496350
rect 583274 496294 583342 496350
rect 583398 496294 583494 496350
rect 582874 496226 583494 496294
rect 582874 496170 582970 496226
rect 583026 496170 583094 496226
rect 583150 496170 583218 496226
rect 583274 496170 583342 496226
rect 583398 496170 583494 496226
rect 582874 496102 583494 496170
rect 582874 496046 582970 496102
rect 583026 496046 583094 496102
rect 583150 496046 583218 496102
rect 583274 496046 583342 496102
rect 583398 496046 583494 496102
rect 582874 495978 583494 496046
rect 582874 495922 582970 495978
rect 583026 495922 583094 495978
rect 583150 495922 583218 495978
rect 583274 495922 583342 495978
rect 583398 495922 583494 495978
rect 582874 478350 583494 495922
rect 582874 478294 582970 478350
rect 583026 478294 583094 478350
rect 583150 478294 583218 478350
rect 583274 478294 583342 478350
rect 583398 478294 583494 478350
rect 582874 478226 583494 478294
rect 582874 478170 582970 478226
rect 583026 478170 583094 478226
rect 583150 478170 583218 478226
rect 583274 478170 583342 478226
rect 583398 478170 583494 478226
rect 582874 478102 583494 478170
rect 582874 478046 582970 478102
rect 583026 478046 583094 478102
rect 583150 478046 583218 478102
rect 583274 478046 583342 478102
rect 583398 478046 583494 478102
rect 582874 477978 583494 478046
rect 582874 477922 582970 477978
rect 583026 477922 583094 477978
rect 583150 477922 583218 477978
rect 583274 477922 583342 477978
rect 583398 477922 583494 477978
rect 582874 460350 583494 477922
rect 582874 460294 582970 460350
rect 583026 460294 583094 460350
rect 583150 460294 583218 460350
rect 583274 460294 583342 460350
rect 583398 460294 583494 460350
rect 582874 460226 583494 460294
rect 582874 460170 582970 460226
rect 583026 460170 583094 460226
rect 583150 460170 583218 460226
rect 583274 460170 583342 460226
rect 583398 460170 583494 460226
rect 582874 460102 583494 460170
rect 582874 460046 582970 460102
rect 583026 460046 583094 460102
rect 583150 460046 583218 460102
rect 583274 460046 583342 460102
rect 583398 460046 583494 460102
rect 582874 459978 583494 460046
rect 582874 459922 582970 459978
rect 583026 459922 583094 459978
rect 583150 459922 583218 459978
rect 583274 459922 583342 459978
rect 583398 459922 583494 459978
rect 582874 442350 583494 459922
rect 582874 442294 582970 442350
rect 583026 442294 583094 442350
rect 583150 442294 583218 442350
rect 583274 442294 583342 442350
rect 583398 442294 583494 442350
rect 582874 442226 583494 442294
rect 582874 442170 582970 442226
rect 583026 442170 583094 442226
rect 583150 442170 583218 442226
rect 583274 442170 583342 442226
rect 583398 442170 583494 442226
rect 582874 442102 583494 442170
rect 582874 442046 582970 442102
rect 583026 442046 583094 442102
rect 583150 442046 583218 442102
rect 583274 442046 583342 442102
rect 583398 442046 583494 442102
rect 582874 441978 583494 442046
rect 582874 441922 582970 441978
rect 583026 441922 583094 441978
rect 583150 441922 583218 441978
rect 583274 441922 583342 441978
rect 583398 441922 583494 441978
rect 582874 424350 583494 441922
rect 582874 424294 582970 424350
rect 583026 424294 583094 424350
rect 583150 424294 583218 424350
rect 583274 424294 583342 424350
rect 583398 424294 583494 424350
rect 582874 424226 583494 424294
rect 582874 424170 582970 424226
rect 583026 424170 583094 424226
rect 583150 424170 583218 424226
rect 583274 424170 583342 424226
rect 583398 424170 583494 424226
rect 582874 424102 583494 424170
rect 582874 424046 582970 424102
rect 583026 424046 583094 424102
rect 583150 424046 583218 424102
rect 583274 424046 583342 424102
rect 583398 424046 583494 424102
rect 582874 423978 583494 424046
rect 582874 423922 582970 423978
rect 583026 423922 583094 423978
rect 583150 423922 583218 423978
rect 583274 423922 583342 423978
rect 583398 423922 583494 423978
rect 582874 406350 583494 423922
rect 582874 406294 582970 406350
rect 583026 406294 583094 406350
rect 583150 406294 583218 406350
rect 583274 406294 583342 406350
rect 583398 406294 583494 406350
rect 582874 406226 583494 406294
rect 582874 406170 582970 406226
rect 583026 406170 583094 406226
rect 583150 406170 583218 406226
rect 583274 406170 583342 406226
rect 583398 406170 583494 406226
rect 582874 406102 583494 406170
rect 582874 406046 582970 406102
rect 583026 406046 583094 406102
rect 583150 406046 583218 406102
rect 583274 406046 583342 406102
rect 583398 406046 583494 406102
rect 582874 405978 583494 406046
rect 582874 405922 582970 405978
rect 583026 405922 583094 405978
rect 583150 405922 583218 405978
rect 583274 405922 583342 405978
rect 583398 405922 583494 405978
rect 582874 388350 583494 405922
rect 582874 388294 582970 388350
rect 583026 388294 583094 388350
rect 583150 388294 583218 388350
rect 583274 388294 583342 388350
rect 583398 388294 583494 388350
rect 582874 388226 583494 388294
rect 582874 388170 582970 388226
rect 583026 388170 583094 388226
rect 583150 388170 583218 388226
rect 583274 388170 583342 388226
rect 583398 388170 583494 388226
rect 582874 388102 583494 388170
rect 582874 388046 582970 388102
rect 583026 388046 583094 388102
rect 583150 388046 583218 388102
rect 583274 388046 583342 388102
rect 583398 388046 583494 388102
rect 582874 387978 583494 388046
rect 582874 387922 582970 387978
rect 583026 387922 583094 387978
rect 583150 387922 583218 387978
rect 583274 387922 583342 387978
rect 583398 387922 583494 387978
rect 582874 370350 583494 387922
rect 582874 370294 582970 370350
rect 583026 370294 583094 370350
rect 583150 370294 583218 370350
rect 583274 370294 583342 370350
rect 583398 370294 583494 370350
rect 582874 370226 583494 370294
rect 582874 370170 582970 370226
rect 583026 370170 583094 370226
rect 583150 370170 583218 370226
rect 583274 370170 583342 370226
rect 583398 370170 583494 370226
rect 582874 370102 583494 370170
rect 582874 370046 582970 370102
rect 583026 370046 583094 370102
rect 583150 370046 583218 370102
rect 583274 370046 583342 370102
rect 583398 370046 583494 370102
rect 582874 369978 583494 370046
rect 582874 369922 582970 369978
rect 583026 369922 583094 369978
rect 583150 369922 583218 369978
rect 583274 369922 583342 369978
rect 583398 369922 583494 369978
rect 582874 352350 583494 369922
rect 582874 352294 582970 352350
rect 583026 352294 583094 352350
rect 583150 352294 583218 352350
rect 583274 352294 583342 352350
rect 583398 352294 583494 352350
rect 582874 352226 583494 352294
rect 582874 352170 582970 352226
rect 583026 352170 583094 352226
rect 583150 352170 583218 352226
rect 583274 352170 583342 352226
rect 583398 352170 583494 352226
rect 582874 352102 583494 352170
rect 582874 352046 582970 352102
rect 583026 352046 583094 352102
rect 583150 352046 583218 352102
rect 583274 352046 583342 352102
rect 583398 352046 583494 352102
rect 582874 351978 583494 352046
rect 582874 351922 582970 351978
rect 583026 351922 583094 351978
rect 583150 351922 583218 351978
rect 583274 351922 583342 351978
rect 583398 351922 583494 351978
rect 582874 334350 583494 351922
rect 582874 334294 582970 334350
rect 583026 334294 583094 334350
rect 583150 334294 583218 334350
rect 583274 334294 583342 334350
rect 583398 334294 583494 334350
rect 582874 334226 583494 334294
rect 582874 334170 582970 334226
rect 583026 334170 583094 334226
rect 583150 334170 583218 334226
rect 583274 334170 583342 334226
rect 583398 334170 583494 334226
rect 582874 334102 583494 334170
rect 582874 334046 582970 334102
rect 583026 334046 583094 334102
rect 583150 334046 583218 334102
rect 583274 334046 583342 334102
rect 583398 334046 583494 334102
rect 582874 333978 583494 334046
rect 582874 333922 582970 333978
rect 583026 333922 583094 333978
rect 583150 333922 583218 333978
rect 583274 333922 583342 333978
rect 583398 333922 583494 333978
rect 582874 316350 583494 333922
rect 582874 316294 582970 316350
rect 583026 316294 583094 316350
rect 583150 316294 583218 316350
rect 583274 316294 583342 316350
rect 583398 316294 583494 316350
rect 582874 316226 583494 316294
rect 582874 316170 582970 316226
rect 583026 316170 583094 316226
rect 583150 316170 583218 316226
rect 583274 316170 583342 316226
rect 583398 316170 583494 316226
rect 582874 316102 583494 316170
rect 582874 316046 582970 316102
rect 583026 316046 583094 316102
rect 583150 316046 583218 316102
rect 583274 316046 583342 316102
rect 583398 316046 583494 316102
rect 582874 315978 583494 316046
rect 582874 315922 582970 315978
rect 583026 315922 583094 315978
rect 583150 315922 583218 315978
rect 583274 315922 583342 315978
rect 583398 315922 583494 315978
rect 582874 298350 583494 315922
rect 582874 298294 582970 298350
rect 583026 298294 583094 298350
rect 583150 298294 583218 298350
rect 583274 298294 583342 298350
rect 583398 298294 583494 298350
rect 582874 298226 583494 298294
rect 582874 298170 582970 298226
rect 583026 298170 583094 298226
rect 583150 298170 583218 298226
rect 583274 298170 583342 298226
rect 583398 298170 583494 298226
rect 582874 298102 583494 298170
rect 582874 298046 582970 298102
rect 583026 298046 583094 298102
rect 583150 298046 583218 298102
rect 583274 298046 583342 298102
rect 583398 298046 583494 298102
rect 582874 297978 583494 298046
rect 582874 297922 582970 297978
rect 583026 297922 583094 297978
rect 583150 297922 583218 297978
rect 583274 297922 583342 297978
rect 583398 297922 583494 297978
rect 582874 280350 583494 297922
rect 582874 280294 582970 280350
rect 583026 280294 583094 280350
rect 583150 280294 583218 280350
rect 583274 280294 583342 280350
rect 583398 280294 583494 280350
rect 582874 280226 583494 280294
rect 582874 280170 582970 280226
rect 583026 280170 583094 280226
rect 583150 280170 583218 280226
rect 583274 280170 583342 280226
rect 583398 280170 583494 280226
rect 582874 280102 583494 280170
rect 582874 280046 582970 280102
rect 583026 280046 583094 280102
rect 583150 280046 583218 280102
rect 583274 280046 583342 280102
rect 583398 280046 583494 280102
rect 582874 279978 583494 280046
rect 582874 279922 582970 279978
rect 583026 279922 583094 279978
rect 583150 279922 583218 279978
rect 583274 279922 583342 279978
rect 583398 279922 583494 279978
rect 582874 262350 583494 279922
rect 582874 262294 582970 262350
rect 583026 262294 583094 262350
rect 583150 262294 583218 262350
rect 583274 262294 583342 262350
rect 583398 262294 583494 262350
rect 582874 262226 583494 262294
rect 582874 262170 582970 262226
rect 583026 262170 583094 262226
rect 583150 262170 583218 262226
rect 583274 262170 583342 262226
rect 583398 262170 583494 262226
rect 582874 262102 583494 262170
rect 582874 262046 582970 262102
rect 583026 262046 583094 262102
rect 583150 262046 583218 262102
rect 583274 262046 583342 262102
rect 583398 262046 583494 262102
rect 582874 261978 583494 262046
rect 582874 261922 582970 261978
rect 583026 261922 583094 261978
rect 583150 261922 583218 261978
rect 583274 261922 583342 261978
rect 583398 261922 583494 261978
rect 582874 244350 583494 261922
rect 582874 244294 582970 244350
rect 583026 244294 583094 244350
rect 583150 244294 583218 244350
rect 583274 244294 583342 244350
rect 583398 244294 583494 244350
rect 582874 244226 583494 244294
rect 582874 244170 582970 244226
rect 583026 244170 583094 244226
rect 583150 244170 583218 244226
rect 583274 244170 583342 244226
rect 583398 244170 583494 244226
rect 582874 244102 583494 244170
rect 582874 244046 582970 244102
rect 583026 244046 583094 244102
rect 583150 244046 583218 244102
rect 583274 244046 583342 244102
rect 583398 244046 583494 244102
rect 582874 243978 583494 244046
rect 582874 243922 582970 243978
rect 583026 243922 583094 243978
rect 583150 243922 583218 243978
rect 583274 243922 583342 243978
rect 583398 243922 583494 243978
rect 582874 226350 583494 243922
rect 582874 226294 582970 226350
rect 583026 226294 583094 226350
rect 583150 226294 583218 226350
rect 583274 226294 583342 226350
rect 583398 226294 583494 226350
rect 582874 226226 583494 226294
rect 582874 226170 582970 226226
rect 583026 226170 583094 226226
rect 583150 226170 583218 226226
rect 583274 226170 583342 226226
rect 583398 226170 583494 226226
rect 582874 226102 583494 226170
rect 582874 226046 582970 226102
rect 583026 226046 583094 226102
rect 583150 226046 583218 226102
rect 583274 226046 583342 226102
rect 583398 226046 583494 226102
rect 582874 225978 583494 226046
rect 582874 225922 582970 225978
rect 583026 225922 583094 225978
rect 583150 225922 583218 225978
rect 583274 225922 583342 225978
rect 583398 225922 583494 225978
rect 582874 208350 583494 225922
rect 582874 208294 582970 208350
rect 583026 208294 583094 208350
rect 583150 208294 583218 208350
rect 583274 208294 583342 208350
rect 583398 208294 583494 208350
rect 582874 208226 583494 208294
rect 582874 208170 582970 208226
rect 583026 208170 583094 208226
rect 583150 208170 583218 208226
rect 583274 208170 583342 208226
rect 583398 208170 583494 208226
rect 582874 208102 583494 208170
rect 582874 208046 582970 208102
rect 583026 208046 583094 208102
rect 583150 208046 583218 208102
rect 583274 208046 583342 208102
rect 583398 208046 583494 208102
rect 582874 207978 583494 208046
rect 582874 207922 582970 207978
rect 583026 207922 583094 207978
rect 583150 207922 583218 207978
rect 583274 207922 583342 207978
rect 583398 207922 583494 207978
rect 582874 190350 583494 207922
rect 582874 190294 582970 190350
rect 583026 190294 583094 190350
rect 583150 190294 583218 190350
rect 583274 190294 583342 190350
rect 583398 190294 583494 190350
rect 582874 190226 583494 190294
rect 582874 190170 582970 190226
rect 583026 190170 583094 190226
rect 583150 190170 583218 190226
rect 583274 190170 583342 190226
rect 583398 190170 583494 190226
rect 582874 190102 583494 190170
rect 582874 190046 582970 190102
rect 583026 190046 583094 190102
rect 583150 190046 583218 190102
rect 583274 190046 583342 190102
rect 583398 190046 583494 190102
rect 582874 189978 583494 190046
rect 582874 189922 582970 189978
rect 583026 189922 583094 189978
rect 583150 189922 583218 189978
rect 583274 189922 583342 189978
rect 583398 189922 583494 189978
rect 582874 172350 583494 189922
rect 582874 172294 582970 172350
rect 583026 172294 583094 172350
rect 583150 172294 583218 172350
rect 583274 172294 583342 172350
rect 583398 172294 583494 172350
rect 582874 172226 583494 172294
rect 582874 172170 582970 172226
rect 583026 172170 583094 172226
rect 583150 172170 583218 172226
rect 583274 172170 583342 172226
rect 583398 172170 583494 172226
rect 582874 172102 583494 172170
rect 582874 172046 582970 172102
rect 583026 172046 583094 172102
rect 583150 172046 583218 172102
rect 583274 172046 583342 172102
rect 583398 172046 583494 172102
rect 582874 171978 583494 172046
rect 582874 171922 582970 171978
rect 583026 171922 583094 171978
rect 583150 171922 583218 171978
rect 583274 171922 583342 171978
rect 583398 171922 583494 171978
rect 582874 154350 583494 171922
rect 582874 154294 582970 154350
rect 583026 154294 583094 154350
rect 583150 154294 583218 154350
rect 583274 154294 583342 154350
rect 583398 154294 583494 154350
rect 582874 154226 583494 154294
rect 582874 154170 582970 154226
rect 583026 154170 583094 154226
rect 583150 154170 583218 154226
rect 583274 154170 583342 154226
rect 583398 154170 583494 154226
rect 582874 154102 583494 154170
rect 582874 154046 582970 154102
rect 583026 154046 583094 154102
rect 583150 154046 583218 154102
rect 583274 154046 583342 154102
rect 583398 154046 583494 154102
rect 582874 153978 583494 154046
rect 582874 153922 582970 153978
rect 583026 153922 583094 153978
rect 583150 153922 583218 153978
rect 583274 153922 583342 153978
rect 583398 153922 583494 153978
rect 582874 136350 583494 153922
rect 582874 136294 582970 136350
rect 583026 136294 583094 136350
rect 583150 136294 583218 136350
rect 583274 136294 583342 136350
rect 583398 136294 583494 136350
rect 582874 136226 583494 136294
rect 582874 136170 582970 136226
rect 583026 136170 583094 136226
rect 583150 136170 583218 136226
rect 583274 136170 583342 136226
rect 583398 136170 583494 136226
rect 582874 136102 583494 136170
rect 582874 136046 582970 136102
rect 583026 136046 583094 136102
rect 583150 136046 583218 136102
rect 583274 136046 583342 136102
rect 583398 136046 583494 136102
rect 582874 135978 583494 136046
rect 582874 135922 582970 135978
rect 583026 135922 583094 135978
rect 583150 135922 583218 135978
rect 583274 135922 583342 135978
rect 583398 135922 583494 135978
rect 582874 118350 583494 135922
rect 582874 118294 582970 118350
rect 583026 118294 583094 118350
rect 583150 118294 583218 118350
rect 583274 118294 583342 118350
rect 583398 118294 583494 118350
rect 582874 118226 583494 118294
rect 582874 118170 582970 118226
rect 583026 118170 583094 118226
rect 583150 118170 583218 118226
rect 583274 118170 583342 118226
rect 583398 118170 583494 118226
rect 582874 118102 583494 118170
rect 582874 118046 582970 118102
rect 583026 118046 583094 118102
rect 583150 118046 583218 118102
rect 583274 118046 583342 118102
rect 583398 118046 583494 118102
rect 582874 117978 583494 118046
rect 582874 117922 582970 117978
rect 583026 117922 583094 117978
rect 583150 117922 583218 117978
rect 583274 117922 583342 117978
rect 583398 117922 583494 117978
rect 582874 100350 583494 117922
rect 582874 100294 582970 100350
rect 583026 100294 583094 100350
rect 583150 100294 583218 100350
rect 583274 100294 583342 100350
rect 583398 100294 583494 100350
rect 582874 100226 583494 100294
rect 582874 100170 582970 100226
rect 583026 100170 583094 100226
rect 583150 100170 583218 100226
rect 583274 100170 583342 100226
rect 583398 100170 583494 100226
rect 582874 100102 583494 100170
rect 582874 100046 582970 100102
rect 583026 100046 583094 100102
rect 583150 100046 583218 100102
rect 583274 100046 583342 100102
rect 583398 100046 583494 100102
rect 582874 99978 583494 100046
rect 582874 99922 582970 99978
rect 583026 99922 583094 99978
rect 583150 99922 583218 99978
rect 583274 99922 583342 99978
rect 583398 99922 583494 99978
rect 582874 82350 583494 99922
rect 582874 82294 582970 82350
rect 583026 82294 583094 82350
rect 583150 82294 583218 82350
rect 583274 82294 583342 82350
rect 583398 82294 583494 82350
rect 582874 82226 583494 82294
rect 582874 82170 582970 82226
rect 583026 82170 583094 82226
rect 583150 82170 583218 82226
rect 583274 82170 583342 82226
rect 583398 82170 583494 82226
rect 582874 82102 583494 82170
rect 582874 82046 582970 82102
rect 583026 82046 583094 82102
rect 583150 82046 583218 82102
rect 583274 82046 583342 82102
rect 583398 82046 583494 82102
rect 582874 81978 583494 82046
rect 582874 81922 582970 81978
rect 583026 81922 583094 81978
rect 583150 81922 583218 81978
rect 583274 81922 583342 81978
rect 583398 81922 583494 81978
rect 582874 64350 583494 81922
rect 582874 64294 582970 64350
rect 583026 64294 583094 64350
rect 583150 64294 583218 64350
rect 583274 64294 583342 64350
rect 583398 64294 583494 64350
rect 582874 64226 583494 64294
rect 582874 64170 582970 64226
rect 583026 64170 583094 64226
rect 583150 64170 583218 64226
rect 583274 64170 583342 64226
rect 583398 64170 583494 64226
rect 582874 64102 583494 64170
rect 582874 64046 582970 64102
rect 583026 64046 583094 64102
rect 583150 64046 583218 64102
rect 583274 64046 583342 64102
rect 583398 64046 583494 64102
rect 582874 63978 583494 64046
rect 582874 63922 582970 63978
rect 583026 63922 583094 63978
rect 583150 63922 583218 63978
rect 583274 63922 583342 63978
rect 583398 63922 583494 63978
rect 582874 46350 583494 63922
rect 582874 46294 582970 46350
rect 583026 46294 583094 46350
rect 583150 46294 583218 46350
rect 583274 46294 583342 46350
rect 583398 46294 583494 46350
rect 582874 46226 583494 46294
rect 582874 46170 582970 46226
rect 583026 46170 583094 46226
rect 583150 46170 583218 46226
rect 583274 46170 583342 46226
rect 583398 46170 583494 46226
rect 582874 46102 583494 46170
rect 582874 46046 582970 46102
rect 583026 46046 583094 46102
rect 583150 46046 583218 46102
rect 583274 46046 583342 46102
rect 583398 46046 583494 46102
rect 582874 45978 583494 46046
rect 582874 45922 582970 45978
rect 583026 45922 583094 45978
rect 583150 45922 583218 45978
rect 583274 45922 583342 45978
rect 583398 45922 583494 45978
rect 582874 28350 583494 45922
rect 582874 28294 582970 28350
rect 583026 28294 583094 28350
rect 583150 28294 583218 28350
rect 583274 28294 583342 28350
rect 583398 28294 583494 28350
rect 582874 28226 583494 28294
rect 582874 28170 582970 28226
rect 583026 28170 583094 28226
rect 583150 28170 583218 28226
rect 583274 28170 583342 28226
rect 583398 28170 583494 28226
rect 582874 28102 583494 28170
rect 582874 28046 582970 28102
rect 583026 28046 583094 28102
rect 583150 28046 583218 28102
rect 583274 28046 583342 28102
rect 583398 28046 583494 28102
rect 582874 27978 583494 28046
rect 582874 27922 582970 27978
rect 583026 27922 583094 27978
rect 583150 27922 583218 27978
rect 583274 27922 583342 27978
rect 583398 27922 583494 27978
rect 582874 10350 583494 27922
rect 582874 10294 582970 10350
rect 583026 10294 583094 10350
rect 583150 10294 583218 10350
rect 583274 10294 583342 10350
rect 583398 10294 583494 10350
rect 582874 10226 583494 10294
rect 582874 10170 582970 10226
rect 583026 10170 583094 10226
rect 583150 10170 583218 10226
rect 583274 10170 583342 10226
rect 583398 10170 583494 10226
rect 582874 10102 583494 10170
rect 582874 10046 582970 10102
rect 583026 10046 583094 10102
rect 583150 10046 583218 10102
rect 583274 10046 583342 10102
rect 583398 10046 583494 10102
rect 582874 9978 583494 10046
rect 582874 9922 582970 9978
rect 583026 9922 583094 9978
rect 583150 9922 583218 9978
rect 583274 9922 583342 9978
rect 583398 9922 583494 9978
rect 582874 -1120 583494 9922
rect 596400 597212 597020 597308
rect 596400 597156 596496 597212
rect 596552 597156 596620 597212
rect 596676 597156 596744 597212
rect 596800 597156 596868 597212
rect 596924 597156 597020 597212
rect 596400 597088 597020 597156
rect 596400 597032 596496 597088
rect 596552 597032 596620 597088
rect 596676 597032 596744 597088
rect 596800 597032 596868 597088
rect 596924 597032 597020 597088
rect 596400 596964 597020 597032
rect 596400 596908 596496 596964
rect 596552 596908 596620 596964
rect 596676 596908 596744 596964
rect 596800 596908 596868 596964
rect 596924 596908 597020 596964
rect 596400 596840 597020 596908
rect 596400 596784 596496 596840
rect 596552 596784 596620 596840
rect 596676 596784 596744 596840
rect 596800 596784 596868 596840
rect 596924 596784 597020 596840
rect 596400 580350 597020 596784
rect 596400 580294 596496 580350
rect 596552 580294 596620 580350
rect 596676 580294 596744 580350
rect 596800 580294 596868 580350
rect 596924 580294 597020 580350
rect 596400 580226 597020 580294
rect 596400 580170 596496 580226
rect 596552 580170 596620 580226
rect 596676 580170 596744 580226
rect 596800 580170 596868 580226
rect 596924 580170 597020 580226
rect 596400 580102 597020 580170
rect 596400 580046 596496 580102
rect 596552 580046 596620 580102
rect 596676 580046 596744 580102
rect 596800 580046 596868 580102
rect 596924 580046 597020 580102
rect 596400 579978 597020 580046
rect 596400 579922 596496 579978
rect 596552 579922 596620 579978
rect 596676 579922 596744 579978
rect 596800 579922 596868 579978
rect 596924 579922 597020 579978
rect 596400 562350 597020 579922
rect 596400 562294 596496 562350
rect 596552 562294 596620 562350
rect 596676 562294 596744 562350
rect 596800 562294 596868 562350
rect 596924 562294 597020 562350
rect 596400 562226 597020 562294
rect 596400 562170 596496 562226
rect 596552 562170 596620 562226
rect 596676 562170 596744 562226
rect 596800 562170 596868 562226
rect 596924 562170 597020 562226
rect 596400 562102 597020 562170
rect 596400 562046 596496 562102
rect 596552 562046 596620 562102
rect 596676 562046 596744 562102
rect 596800 562046 596868 562102
rect 596924 562046 597020 562102
rect 596400 561978 597020 562046
rect 596400 561922 596496 561978
rect 596552 561922 596620 561978
rect 596676 561922 596744 561978
rect 596800 561922 596868 561978
rect 596924 561922 597020 561978
rect 596400 544350 597020 561922
rect 596400 544294 596496 544350
rect 596552 544294 596620 544350
rect 596676 544294 596744 544350
rect 596800 544294 596868 544350
rect 596924 544294 597020 544350
rect 596400 544226 597020 544294
rect 596400 544170 596496 544226
rect 596552 544170 596620 544226
rect 596676 544170 596744 544226
rect 596800 544170 596868 544226
rect 596924 544170 597020 544226
rect 596400 544102 597020 544170
rect 596400 544046 596496 544102
rect 596552 544046 596620 544102
rect 596676 544046 596744 544102
rect 596800 544046 596868 544102
rect 596924 544046 597020 544102
rect 596400 543978 597020 544046
rect 596400 543922 596496 543978
rect 596552 543922 596620 543978
rect 596676 543922 596744 543978
rect 596800 543922 596868 543978
rect 596924 543922 597020 543978
rect 596400 526350 597020 543922
rect 596400 526294 596496 526350
rect 596552 526294 596620 526350
rect 596676 526294 596744 526350
rect 596800 526294 596868 526350
rect 596924 526294 597020 526350
rect 596400 526226 597020 526294
rect 596400 526170 596496 526226
rect 596552 526170 596620 526226
rect 596676 526170 596744 526226
rect 596800 526170 596868 526226
rect 596924 526170 597020 526226
rect 596400 526102 597020 526170
rect 596400 526046 596496 526102
rect 596552 526046 596620 526102
rect 596676 526046 596744 526102
rect 596800 526046 596868 526102
rect 596924 526046 597020 526102
rect 596400 525978 597020 526046
rect 596400 525922 596496 525978
rect 596552 525922 596620 525978
rect 596676 525922 596744 525978
rect 596800 525922 596868 525978
rect 596924 525922 597020 525978
rect 596400 508350 597020 525922
rect 596400 508294 596496 508350
rect 596552 508294 596620 508350
rect 596676 508294 596744 508350
rect 596800 508294 596868 508350
rect 596924 508294 597020 508350
rect 596400 508226 597020 508294
rect 596400 508170 596496 508226
rect 596552 508170 596620 508226
rect 596676 508170 596744 508226
rect 596800 508170 596868 508226
rect 596924 508170 597020 508226
rect 596400 508102 597020 508170
rect 596400 508046 596496 508102
rect 596552 508046 596620 508102
rect 596676 508046 596744 508102
rect 596800 508046 596868 508102
rect 596924 508046 597020 508102
rect 596400 507978 597020 508046
rect 596400 507922 596496 507978
rect 596552 507922 596620 507978
rect 596676 507922 596744 507978
rect 596800 507922 596868 507978
rect 596924 507922 597020 507978
rect 596400 490350 597020 507922
rect 596400 490294 596496 490350
rect 596552 490294 596620 490350
rect 596676 490294 596744 490350
rect 596800 490294 596868 490350
rect 596924 490294 597020 490350
rect 596400 490226 597020 490294
rect 596400 490170 596496 490226
rect 596552 490170 596620 490226
rect 596676 490170 596744 490226
rect 596800 490170 596868 490226
rect 596924 490170 597020 490226
rect 596400 490102 597020 490170
rect 596400 490046 596496 490102
rect 596552 490046 596620 490102
rect 596676 490046 596744 490102
rect 596800 490046 596868 490102
rect 596924 490046 597020 490102
rect 596400 489978 597020 490046
rect 596400 489922 596496 489978
rect 596552 489922 596620 489978
rect 596676 489922 596744 489978
rect 596800 489922 596868 489978
rect 596924 489922 597020 489978
rect 596400 472350 597020 489922
rect 596400 472294 596496 472350
rect 596552 472294 596620 472350
rect 596676 472294 596744 472350
rect 596800 472294 596868 472350
rect 596924 472294 597020 472350
rect 596400 472226 597020 472294
rect 596400 472170 596496 472226
rect 596552 472170 596620 472226
rect 596676 472170 596744 472226
rect 596800 472170 596868 472226
rect 596924 472170 597020 472226
rect 596400 472102 597020 472170
rect 596400 472046 596496 472102
rect 596552 472046 596620 472102
rect 596676 472046 596744 472102
rect 596800 472046 596868 472102
rect 596924 472046 597020 472102
rect 596400 471978 597020 472046
rect 596400 471922 596496 471978
rect 596552 471922 596620 471978
rect 596676 471922 596744 471978
rect 596800 471922 596868 471978
rect 596924 471922 597020 471978
rect 596400 454350 597020 471922
rect 596400 454294 596496 454350
rect 596552 454294 596620 454350
rect 596676 454294 596744 454350
rect 596800 454294 596868 454350
rect 596924 454294 597020 454350
rect 596400 454226 597020 454294
rect 596400 454170 596496 454226
rect 596552 454170 596620 454226
rect 596676 454170 596744 454226
rect 596800 454170 596868 454226
rect 596924 454170 597020 454226
rect 596400 454102 597020 454170
rect 596400 454046 596496 454102
rect 596552 454046 596620 454102
rect 596676 454046 596744 454102
rect 596800 454046 596868 454102
rect 596924 454046 597020 454102
rect 596400 453978 597020 454046
rect 596400 453922 596496 453978
rect 596552 453922 596620 453978
rect 596676 453922 596744 453978
rect 596800 453922 596868 453978
rect 596924 453922 597020 453978
rect 596400 436350 597020 453922
rect 596400 436294 596496 436350
rect 596552 436294 596620 436350
rect 596676 436294 596744 436350
rect 596800 436294 596868 436350
rect 596924 436294 597020 436350
rect 596400 436226 597020 436294
rect 596400 436170 596496 436226
rect 596552 436170 596620 436226
rect 596676 436170 596744 436226
rect 596800 436170 596868 436226
rect 596924 436170 597020 436226
rect 596400 436102 597020 436170
rect 596400 436046 596496 436102
rect 596552 436046 596620 436102
rect 596676 436046 596744 436102
rect 596800 436046 596868 436102
rect 596924 436046 597020 436102
rect 596400 435978 597020 436046
rect 596400 435922 596496 435978
rect 596552 435922 596620 435978
rect 596676 435922 596744 435978
rect 596800 435922 596868 435978
rect 596924 435922 597020 435978
rect 596400 418350 597020 435922
rect 596400 418294 596496 418350
rect 596552 418294 596620 418350
rect 596676 418294 596744 418350
rect 596800 418294 596868 418350
rect 596924 418294 597020 418350
rect 596400 418226 597020 418294
rect 596400 418170 596496 418226
rect 596552 418170 596620 418226
rect 596676 418170 596744 418226
rect 596800 418170 596868 418226
rect 596924 418170 597020 418226
rect 596400 418102 597020 418170
rect 596400 418046 596496 418102
rect 596552 418046 596620 418102
rect 596676 418046 596744 418102
rect 596800 418046 596868 418102
rect 596924 418046 597020 418102
rect 596400 417978 597020 418046
rect 596400 417922 596496 417978
rect 596552 417922 596620 417978
rect 596676 417922 596744 417978
rect 596800 417922 596868 417978
rect 596924 417922 597020 417978
rect 596400 400350 597020 417922
rect 596400 400294 596496 400350
rect 596552 400294 596620 400350
rect 596676 400294 596744 400350
rect 596800 400294 596868 400350
rect 596924 400294 597020 400350
rect 596400 400226 597020 400294
rect 596400 400170 596496 400226
rect 596552 400170 596620 400226
rect 596676 400170 596744 400226
rect 596800 400170 596868 400226
rect 596924 400170 597020 400226
rect 596400 400102 597020 400170
rect 596400 400046 596496 400102
rect 596552 400046 596620 400102
rect 596676 400046 596744 400102
rect 596800 400046 596868 400102
rect 596924 400046 597020 400102
rect 596400 399978 597020 400046
rect 596400 399922 596496 399978
rect 596552 399922 596620 399978
rect 596676 399922 596744 399978
rect 596800 399922 596868 399978
rect 596924 399922 597020 399978
rect 596400 382350 597020 399922
rect 596400 382294 596496 382350
rect 596552 382294 596620 382350
rect 596676 382294 596744 382350
rect 596800 382294 596868 382350
rect 596924 382294 597020 382350
rect 596400 382226 597020 382294
rect 596400 382170 596496 382226
rect 596552 382170 596620 382226
rect 596676 382170 596744 382226
rect 596800 382170 596868 382226
rect 596924 382170 597020 382226
rect 596400 382102 597020 382170
rect 596400 382046 596496 382102
rect 596552 382046 596620 382102
rect 596676 382046 596744 382102
rect 596800 382046 596868 382102
rect 596924 382046 597020 382102
rect 596400 381978 597020 382046
rect 596400 381922 596496 381978
rect 596552 381922 596620 381978
rect 596676 381922 596744 381978
rect 596800 381922 596868 381978
rect 596924 381922 597020 381978
rect 596400 364350 597020 381922
rect 596400 364294 596496 364350
rect 596552 364294 596620 364350
rect 596676 364294 596744 364350
rect 596800 364294 596868 364350
rect 596924 364294 597020 364350
rect 596400 364226 597020 364294
rect 596400 364170 596496 364226
rect 596552 364170 596620 364226
rect 596676 364170 596744 364226
rect 596800 364170 596868 364226
rect 596924 364170 597020 364226
rect 596400 364102 597020 364170
rect 596400 364046 596496 364102
rect 596552 364046 596620 364102
rect 596676 364046 596744 364102
rect 596800 364046 596868 364102
rect 596924 364046 597020 364102
rect 596400 363978 597020 364046
rect 596400 363922 596496 363978
rect 596552 363922 596620 363978
rect 596676 363922 596744 363978
rect 596800 363922 596868 363978
rect 596924 363922 597020 363978
rect 596400 346350 597020 363922
rect 596400 346294 596496 346350
rect 596552 346294 596620 346350
rect 596676 346294 596744 346350
rect 596800 346294 596868 346350
rect 596924 346294 597020 346350
rect 596400 346226 597020 346294
rect 596400 346170 596496 346226
rect 596552 346170 596620 346226
rect 596676 346170 596744 346226
rect 596800 346170 596868 346226
rect 596924 346170 597020 346226
rect 596400 346102 597020 346170
rect 596400 346046 596496 346102
rect 596552 346046 596620 346102
rect 596676 346046 596744 346102
rect 596800 346046 596868 346102
rect 596924 346046 597020 346102
rect 596400 345978 597020 346046
rect 596400 345922 596496 345978
rect 596552 345922 596620 345978
rect 596676 345922 596744 345978
rect 596800 345922 596868 345978
rect 596924 345922 597020 345978
rect 596400 328350 597020 345922
rect 596400 328294 596496 328350
rect 596552 328294 596620 328350
rect 596676 328294 596744 328350
rect 596800 328294 596868 328350
rect 596924 328294 597020 328350
rect 596400 328226 597020 328294
rect 596400 328170 596496 328226
rect 596552 328170 596620 328226
rect 596676 328170 596744 328226
rect 596800 328170 596868 328226
rect 596924 328170 597020 328226
rect 596400 328102 597020 328170
rect 596400 328046 596496 328102
rect 596552 328046 596620 328102
rect 596676 328046 596744 328102
rect 596800 328046 596868 328102
rect 596924 328046 597020 328102
rect 596400 327978 597020 328046
rect 596400 327922 596496 327978
rect 596552 327922 596620 327978
rect 596676 327922 596744 327978
rect 596800 327922 596868 327978
rect 596924 327922 597020 327978
rect 596400 310350 597020 327922
rect 596400 310294 596496 310350
rect 596552 310294 596620 310350
rect 596676 310294 596744 310350
rect 596800 310294 596868 310350
rect 596924 310294 597020 310350
rect 596400 310226 597020 310294
rect 596400 310170 596496 310226
rect 596552 310170 596620 310226
rect 596676 310170 596744 310226
rect 596800 310170 596868 310226
rect 596924 310170 597020 310226
rect 596400 310102 597020 310170
rect 596400 310046 596496 310102
rect 596552 310046 596620 310102
rect 596676 310046 596744 310102
rect 596800 310046 596868 310102
rect 596924 310046 597020 310102
rect 596400 309978 597020 310046
rect 596400 309922 596496 309978
rect 596552 309922 596620 309978
rect 596676 309922 596744 309978
rect 596800 309922 596868 309978
rect 596924 309922 597020 309978
rect 596400 292350 597020 309922
rect 596400 292294 596496 292350
rect 596552 292294 596620 292350
rect 596676 292294 596744 292350
rect 596800 292294 596868 292350
rect 596924 292294 597020 292350
rect 596400 292226 597020 292294
rect 596400 292170 596496 292226
rect 596552 292170 596620 292226
rect 596676 292170 596744 292226
rect 596800 292170 596868 292226
rect 596924 292170 597020 292226
rect 596400 292102 597020 292170
rect 596400 292046 596496 292102
rect 596552 292046 596620 292102
rect 596676 292046 596744 292102
rect 596800 292046 596868 292102
rect 596924 292046 597020 292102
rect 596400 291978 597020 292046
rect 596400 291922 596496 291978
rect 596552 291922 596620 291978
rect 596676 291922 596744 291978
rect 596800 291922 596868 291978
rect 596924 291922 597020 291978
rect 596400 274350 597020 291922
rect 596400 274294 596496 274350
rect 596552 274294 596620 274350
rect 596676 274294 596744 274350
rect 596800 274294 596868 274350
rect 596924 274294 597020 274350
rect 596400 274226 597020 274294
rect 596400 274170 596496 274226
rect 596552 274170 596620 274226
rect 596676 274170 596744 274226
rect 596800 274170 596868 274226
rect 596924 274170 597020 274226
rect 596400 274102 597020 274170
rect 596400 274046 596496 274102
rect 596552 274046 596620 274102
rect 596676 274046 596744 274102
rect 596800 274046 596868 274102
rect 596924 274046 597020 274102
rect 596400 273978 597020 274046
rect 596400 273922 596496 273978
rect 596552 273922 596620 273978
rect 596676 273922 596744 273978
rect 596800 273922 596868 273978
rect 596924 273922 597020 273978
rect 596400 256350 597020 273922
rect 596400 256294 596496 256350
rect 596552 256294 596620 256350
rect 596676 256294 596744 256350
rect 596800 256294 596868 256350
rect 596924 256294 597020 256350
rect 596400 256226 597020 256294
rect 596400 256170 596496 256226
rect 596552 256170 596620 256226
rect 596676 256170 596744 256226
rect 596800 256170 596868 256226
rect 596924 256170 597020 256226
rect 596400 256102 597020 256170
rect 596400 256046 596496 256102
rect 596552 256046 596620 256102
rect 596676 256046 596744 256102
rect 596800 256046 596868 256102
rect 596924 256046 597020 256102
rect 596400 255978 597020 256046
rect 596400 255922 596496 255978
rect 596552 255922 596620 255978
rect 596676 255922 596744 255978
rect 596800 255922 596868 255978
rect 596924 255922 597020 255978
rect 596400 238350 597020 255922
rect 596400 238294 596496 238350
rect 596552 238294 596620 238350
rect 596676 238294 596744 238350
rect 596800 238294 596868 238350
rect 596924 238294 597020 238350
rect 596400 238226 597020 238294
rect 596400 238170 596496 238226
rect 596552 238170 596620 238226
rect 596676 238170 596744 238226
rect 596800 238170 596868 238226
rect 596924 238170 597020 238226
rect 596400 238102 597020 238170
rect 596400 238046 596496 238102
rect 596552 238046 596620 238102
rect 596676 238046 596744 238102
rect 596800 238046 596868 238102
rect 596924 238046 597020 238102
rect 596400 237978 597020 238046
rect 596400 237922 596496 237978
rect 596552 237922 596620 237978
rect 596676 237922 596744 237978
rect 596800 237922 596868 237978
rect 596924 237922 597020 237978
rect 596400 220350 597020 237922
rect 596400 220294 596496 220350
rect 596552 220294 596620 220350
rect 596676 220294 596744 220350
rect 596800 220294 596868 220350
rect 596924 220294 597020 220350
rect 596400 220226 597020 220294
rect 596400 220170 596496 220226
rect 596552 220170 596620 220226
rect 596676 220170 596744 220226
rect 596800 220170 596868 220226
rect 596924 220170 597020 220226
rect 596400 220102 597020 220170
rect 596400 220046 596496 220102
rect 596552 220046 596620 220102
rect 596676 220046 596744 220102
rect 596800 220046 596868 220102
rect 596924 220046 597020 220102
rect 596400 219978 597020 220046
rect 596400 219922 596496 219978
rect 596552 219922 596620 219978
rect 596676 219922 596744 219978
rect 596800 219922 596868 219978
rect 596924 219922 597020 219978
rect 596400 202350 597020 219922
rect 596400 202294 596496 202350
rect 596552 202294 596620 202350
rect 596676 202294 596744 202350
rect 596800 202294 596868 202350
rect 596924 202294 597020 202350
rect 596400 202226 597020 202294
rect 596400 202170 596496 202226
rect 596552 202170 596620 202226
rect 596676 202170 596744 202226
rect 596800 202170 596868 202226
rect 596924 202170 597020 202226
rect 596400 202102 597020 202170
rect 596400 202046 596496 202102
rect 596552 202046 596620 202102
rect 596676 202046 596744 202102
rect 596800 202046 596868 202102
rect 596924 202046 597020 202102
rect 596400 201978 597020 202046
rect 596400 201922 596496 201978
rect 596552 201922 596620 201978
rect 596676 201922 596744 201978
rect 596800 201922 596868 201978
rect 596924 201922 597020 201978
rect 596400 184350 597020 201922
rect 596400 184294 596496 184350
rect 596552 184294 596620 184350
rect 596676 184294 596744 184350
rect 596800 184294 596868 184350
rect 596924 184294 597020 184350
rect 596400 184226 597020 184294
rect 596400 184170 596496 184226
rect 596552 184170 596620 184226
rect 596676 184170 596744 184226
rect 596800 184170 596868 184226
rect 596924 184170 597020 184226
rect 596400 184102 597020 184170
rect 596400 184046 596496 184102
rect 596552 184046 596620 184102
rect 596676 184046 596744 184102
rect 596800 184046 596868 184102
rect 596924 184046 597020 184102
rect 596400 183978 597020 184046
rect 596400 183922 596496 183978
rect 596552 183922 596620 183978
rect 596676 183922 596744 183978
rect 596800 183922 596868 183978
rect 596924 183922 597020 183978
rect 596400 166350 597020 183922
rect 596400 166294 596496 166350
rect 596552 166294 596620 166350
rect 596676 166294 596744 166350
rect 596800 166294 596868 166350
rect 596924 166294 597020 166350
rect 596400 166226 597020 166294
rect 596400 166170 596496 166226
rect 596552 166170 596620 166226
rect 596676 166170 596744 166226
rect 596800 166170 596868 166226
rect 596924 166170 597020 166226
rect 596400 166102 597020 166170
rect 596400 166046 596496 166102
rect 596552 166046 596620 166102
rect 596676 166046 596744 166102
rect 596800 166046 596868 166102
rect 596924 166046 597020 166102
rect 596400 165978 597020 166046
rect 596400 165922 596496 165978
rect 596552 165922 596620 165978
rect 596676 165922 596744 165978
rect 596800 165922 596868 165978
rect 596924 165922 597020 165978
rect 596400 148350 597020 165922
rect 596400 148294 596496 148350
rect 596552 148294 596620 148350
rect 596676 148294 596744 148350
rect 596800 148294 596868 148350
rect 596924 148294 597020 148350
rect 596400 148226 597020 148294
rect 596400 148170 596496 148226
rect 596552 148170 596620 148226
rect 596676 148170 596744 148226
rect 596800 148170 596868 148226
rect 596924 148170 597020 148226
rect 596400 148102 597020 148170
rect 596400 148046 596496 148102
rect 596552 148046 596620 148102
rect 596676 148046 596744 148102
rect 596800 148046 596868 148102
rect 596924 148046 597020 148102
rect 596400 147978 597020 148046
rect 596400 147922 596496 147978
rect 596552 147922 596620 147978
rect 596676 147922 596744 147978
rect 596800 147922 596868 147978
rect 596924 147922 597020 147978
rect 596400 130350 597020 147922
rect 596400 130294 596496 130350
rect 596552 130294 596620 130350
rect 596676 130294 596744 130350
rect 596800 130294 596868 130350
rect 596924 130294 597020 130350
rect 596400 130226 597020 130294
rect 596400 130170 596496 130226
rect 596552 130170 596620 130226
rect 596676 130170 596744 130226
rect 596800 130170 596868 130226
rect 596924 130170 597020 130226
rect 596400 130102 597020 130170
rect 596400 130046 596496 130102
rect 596552 130046 596620 130102
rect 596676 130046 596744 130102
rect 596800 130046 596868 130102
rect 596924 130046 597020 130102
rect 596400 129978 597020 130046
rect 596400 129922 596496 129978
rect 596552 129922 596620 129978
rect 596676 129922 596744 129978
rect 596800 129922 596868 129978
rect 596924 129922 597020 129978
rect 596400 112350 597020 129922
rect 596400 112294 596496 112350
rect 596552 112294 596620 112350
rect 596676 112294 596744 112350
rect 596800 112294 596868 112350
rect 596924 112294 597020 112350
rect 596400 112226 597020 112294
rect 596400 112170 596496 112226
rect 596552 112170 596620 112226
rect 596676 112170 596744 112226
rect 596800 112170 596868 112226
rect 596924 112170 597020 112226
rect 596400 112102 597020 112170
rect 596400 112046 596496 112102
rect 596552 112046 596620 112102
rect 596676 112046 596744 112102
rect 596800 112046 596868 112102
rect 596924 112046 597020 112102
rect 596400 111978 597020 112046
rect 596400 111922 596496 111978
rect 596552 111922 596620 111978
rect 596676 111922 596744 111978
rect 596800 111922 596868 111978
rect 596924 111922 597020 111978
rect 596400 94350 597020 111922
rect 596400 94294 596496 94350
rect 596552 94294 596620 94350
rect 596676 94294 596744 94350
rect 596800 94294 596868 94350
rect 596924 94294 597020 94350
rect 596400 94226 597020 94294
rect 596400 94170 596496 94226
rect 596552 94170 596620 94226
rect 596676 94170 596744 94226
rect 596800 94170 596868 94226
rect 596924 94170 597020 94226
rect 596400 94102 597020 94170
rect 596400 94046 596496 94102
rect 596552 94046 596620 94102
rect 596676 94046 596744 94102
rect 596800 94046 596868 94102
rect 596924 94046 597020 94102
rect 596400 93978 597020 94046
rect 596400 93922 596496 93978
rect 596552 93922 596620 93978
rect 596676 93922 596744 93978
rect 596800 93922 596868 93978
rect 596924 93922 597020 93978
rect 596400 76350 597020 93922
rect 596400 76294 596496 76350
rect 596552 76294 596620 76350
rect 596676 76294 596744 76350
rect 596800 76294 596868 76350
rect 596924 76294 597020 76350
rect 596400 76226 597020 76294
rect 596400 76170 596496 76226
rect 596552 76170 596620 76226
rect 596676 76170 596744 76226
rect 596800 76170 596868 76226
rect 596924 76170 597020 76226
rect 596400 76102 597020 76170
rect 596400 76046 596496 76102
rect 596552 76046 596620 76102
rect 596676 76046 596744 76102
rect 596800 76046 596868 76102
rect 596924 76046 597020 76102
rect 596400 75978 597020 76046
rect 596400 75922 596496 75978
rect 596552 75922 596620 75978
rect 596676 75922 596744 75978
rect 596800 75922 596868 75978
rect 596924 75922 597020 75978
rect 596400 58350 597020 75922
rect 596400 58294 596496 58350
rect 596552 58294 596620 58350
rect 596676 58294 596744 58350
rect 596800 58294 596868 58350
rect 596924 58294 597020 58350
rect 596400 58226 597020 58294
rect 596400 58170 596496 58226
rect 596552 58170 596620 58226
rect 596676 58170 596744 58226
rect 596800 58170 596868 58226
rect 596924 58170 597020 58226
rect 596400 58102 597020 58170
rect 596400 58046 596496 58102
rect 596552 58046 596620 58102
rect 596676 58046 596744 58102
rect 596800 58046 596868 58102
rect 596924 58046 597020 58102
rect 596400 57978 597020 58046
rect 596400 57922 596496 57978
rect 596552 57922 596620 57978
rect 596676 57922 596744 57978
rect 596800 57922 596868 57978
rect 596924 57922 597020 57978
rect 596400 40350 597020 57922
rect 596400 40294 596496 40350
rect 596552 40294 596620 40350
rect 596676 40294 596744 40350
rect 596800 40294 596868 40350
rect 596924 40294 597020 40350
rect 596400 40226 597020 40294
rect 596400 40170 596496 40226
rect 596552 40170 596620 40226
rect 596676 40170 596744 40226
rect 596800 40170 596868 40226
rect 596924 40170 597020 40226
rect 596400 40102 597020 40170
rect 596400 40046 596496 40102
rect 596552 40046 596620 40102
rect 596676 40046 596744 40102
rect 596800 40046 596868 40102
rect 596924 40046 597020 40102
rect 596400 39978 597020 40046
rect 596400 39922 596496 39978
rect 596552 39922 596620 39978
rect 596676 39922 596744 39978
rect 596800 39922 596868 39978
rect 596924 39922 597020 39978
rect 596400 22350 597020 39922
rect 596400 22294 596496 22350
rect 596552 22294 596620 22350
rect 596676 22294 596744 22350
rect 596800 22294 596868 22350
rect 596924 22294 597020 22350
rect 596400 22226 597020 22294
rect 596400 22170 596496 22226
rect 596552 22170 596620 22226
rect 596676 22170 596744 22226
rect 596800 22170 596868 22226
rect 596924 22170 597020 22226
rect 596400 22102 597020 22170
rect 596400 22046 596496 22102
rect 596552 22046 596620 22102
rect 596676 22046 596744 22102
rect 596800 22046 596868 22102
rect 596924 22046 597020 22102
rect 596400 21978 597020 22046
rect 596400 21922 596496 21978
rect 596552 21922 596620 21978
rect 596676 21922 596744 21978
rect 596800 21922 596868 21978
rect 596924 21922 597020 21978
rect 596400 4350 597020 21922
rect 596400 4294 596496 4350
rect 596552 4294 596620 4350
rect 596676 4294 596744 4350
rect 596800 4294 596868 4350
rect 596924 4294 597020 4350
rect 596400 4226 597020 4294
rect 596400 4170 596496 4226
rect 596552 4170 596620 4226
rect 596676 4170 596744 4226
rect 596800 4170 596868 4226
rect 596924 4170 597020 4226
rect 596400 4102 597020 4170
rect 596400 4046 596496 4102
rect 596552 4046 596620 4102
rect 596676 4046 596744 4102
rect 596800 4046 596868 4102
rect 596924 4046 597020 4102
rect 596400 3978 597020 4046
rect 596400 3922 596496 3978
rect 596552 3922 596620 3978
rect 596676 3922 596744 3978
rect 596800 3922 596868 3978
rect 596924 3922 597020 3978
rect 596400 -160 597020 3922
rect 596400 -216 596496 -160
rect 596552 -216 596620 -160
rect 596676 -216 596744 -160
rect 596800 -216 596868 -160
rect 596924 -216 597020 -160
rect 596400 -284 597020 -216
rect 596400 -340 596496 -284
rect 596552 -340 596620 -284
rect 596676 -340 596744 -284
rect 596800 -340 596868 -284
rect 596924 -340 597020 -284
rect 596400 -408 597020 -340
rect 596400 -464 596496 -408
rect 596552 -464 596620 -408
rect 596676 -464 596744 -408
rect 596800 -464 596868 -408
rect 596924 -464 597020 -408
rect 596400 -532 597020 -464
rect 596400 -588 596496 -532
rect 596552 -588 596620 -532
rect 596676 -588 596744 -532
rect 596800 -588 596868 -532
rect 596924 -588 597020 -532
rect 596400 -684 597020 -588
rect 597360 586350 597980 597744
rect 597360 586294 597456 586350
rect 597512 586294 597580 586350
rect 597636 586294 597704 586350
rect 597760 586294 597828 586350
rect 597884 586294 597980 586350
rect 597360 586226 597980 586294
rect 597360 586170 597456 586226
rect 597512 586170 597580 586226
rect 597636 586170 597704 586226
rect 597760 586170 597828 586226
rect 597884 586170 597980 586226
rect 597360 586102 597980 586170
rect 597360 586046 597456 586102
rect 597512 586046 597580 586102
rect 597636 586046 597704 586102
rect 597760 586046 597828 586102
rect 597884 586046 597980 586102
rect 597360 585978 597980 586046
rect 597360 585922 597456 585978
rect 597512 585922 597580 585978
rect 597636 585922 597704 585978
rect 597760 585922 597828 585978
rect 597884 585922 597980 585978
rect 597360 568350 597980 585922
rect 597360 568294 597456 568350
rect 597512 568294 597580 568350
rect 597636 568294 597704 568350
rect 597760 568294 597828 568350
rect 597884 568294 597980 568350
rect 597360 568226 597980 568294
rect 597360 568170 597456 568226
rect 597512 568170 597580 568226
rect 597636 568170 597704 568226
rect 597760 568170 597828 568226
rect 597884 568170 597980 568226
rect 597360 568102 597980 568170
rect 597360 568046 597456 568102
rect 597512 568046 597580 568102
rect 597636 568046 597704 568102
rect 597760 568046 597828 568102
rect 597884 568046 597980 568102
rect 597360 567978 597980 568046
rect 597360 567922 597456 567978
rect 597512 567922 597580 567978
rect 597636 567922 597704 567978
rect 597760 567922 597828 567978
rect 597884 567922 597980 567978
rect 597360 550350 597980 567922
rect 597360 550294 597456 550350
rect 597512 550294 597580 550350
rect 597636 550294 597704 550350
rect 597760 550294 597828 550350
rect 597884 550294 597980 550350
rect 597360 550226 597980 550294
rect 597360 550170 597456 550226
rect 597512 550170 597580 550226
rect 597636 550170 597704 550226
rect 597760 550170 597828 550226
rect 597884 550170 597980 550226
rect 597360 550102 597980 550170
rect 597360 550046 597456 550102
rect 597512 550046 597580 550102
rect 597636 550046 597704 550102
rect 597760 550046 597828 550102
rect 597884 550046 597980 550102
rect 597360 549978 597980 550046
rect 597360 549922 597456 549978
rect 597512 549922 597580 549978
rect 597636 549922 597704 549978
rect 597760 549922 597828 549978
rect 597884 549922 597980 549978
rect 597360 532350 597980 549922
rect 597360 532294 597456 532350
rect 597512 532294 597580 532350
rect 597636 532294 597704 532350
rect 597760 532294 597828 532350
rect 597884 532294 597980 532350
rect 597360 532226 597980 532294
rect 597360 532170 597456 532226
rect 597512 532170 597580 532226
rect 597636 532170 597704 532226
rect 597760 532170 597828 532226
rect 597884 532170 597980 532226
rect 597360 532102 597980 532170
rect 597360 532046 597456 532102
rect 597512 532046 597580 532102
rect 597636 532046 597704 532102
rect 597760 532046 597828 532102
rect 597884 532046 597980 532102
rect 597360 531978 597980 532046
rect 597360 531922 597456 531978
rect 597512 531922 597580 531978
rect 597636 531922 597704 531978
rect 597760 531922 597828 531978
rect 597884 531922 597980 531978
rect 597360 514350 597980 531922
rect 597360 514294 597456 514350
rect 597512 514294 597580 514350
rect 597636 514294 597704 514350
rect 597760 514294 597828 514350
rect 597884 514294 597980 514350
rect 597360 514226 597980 514294
rect 597360 514170 597456 514226
rect 597512 514170 597580 514226
rect 597636 514170 597704 514226
rect 597760 514170 597828 514226
rect 597884 514170 597980 514226
rect 597360 514102 597980 514170
rect 597360 514046 597456 514102
rect 597512 514046 597580 514102
rect 597636 514046 597704 514102
rect 597760 514046 597828 514102
rect 597884 514046 597980 514102
rect 597360 513978 597980 514046
rect 597360 513922 597456 513978
rect 597512 513922 597580 513978
rect 597636 513922 597704 513978
rect 597760 513922 597828 513978
rect 597884 513922 597980 513978
rect 597360 496350 597980 513922
rect 597360 496294 597456 496350
rect 597512 496294 597580 496350
rect 597636 496294 597704 496350
rect 597760 496294 597828 496350
rect 597884 496294 597980 496350
rect 597360 496226 597980 496294
rect 597360 496170 597456 496226
rect 597512 496170 597580 496226
rect 597636 496170 597704 496226
rect 597760 496170 597828 496226
rect 597884 496170 597980 496226
rect 597360 496102 597980 496170
rect 597360 496046 597456 496102
rect 597512 496046 597580 496102
rect 597636 496046 597704 496102
rect 597760 496046 597828 496102
rect 597884 496046 597980 496102
rect 597360 495978 597980 496046
rect 597360 495922 597456 495978
rect 597512 495922 597580 495978
rect 597636 495922 597704 495978
rect 597760 495922 597828 495978
rect 597884 495922 597980 495978
rect 597360 478350 597980 495922
rect 597360 478294 597456 478350
rect 597512 478294 597580 478350
rect 597636 478294 597704 478350
rect 597760 478294 597828 478350
rect 597884 478294 597980 478350
rect 597360 478226 597980 478294
rect 597360 478170 597456 478226
rect 597512 478170 597580 478226
rect 597636 478170 597704 478226
rect 597760 478170 597828 478226
rect 597884 478170 597980 478226
rect 597360 478102 597980 478170
rect 597360 478046 597456 478102
rect 597512 478046 597580 478102
rect 597636 478046 597704 478102
rect 597760 478046 597828 478102
rect 597884 478046 597980 478102
rect 597360 477978 597980 478046
rect 597360 477922 597456 477978
rect 597512 477922 597580 477978
rect 597636 477922 597704 477978
rect 597760 477922 597828 477978
rect 597884 477922 597980 477978
rect 597360 460350 597980 477922
rect 597360 460294 597456 460350
rect 597512 460294 597580 460350
rect 597636 460294 597704 460350
rect 597760 460294 597828 460350
rect 597884 460294 597980 460350
rect 597360 460226 597980 460294
rect 597360 460170 597456 460226
rect 597512 460170 597580 460226
rect 597636 460170 597704 460226
rect 597760 460170 597828 460226
rect 597884 460170 597980 460226
rect 597360 460102 597980 460170
rect 597360 460046 597456 460102
rect 597512 460046 597580 460102
rect 597636 460046 597704 460102
rect 597760 460046 597828 460102
rect 597884 460046 597980 460102
rect 597360 459978 597980 460046
rect 597360 459922 597456 459978
rect 597512 459922 597580 459978
rect 597636 459922 597704 459978
rect 597760 459922 597828 459978
rect 597884 459922 597980 459978
rect 597360 442350 597980 459922
rect 597360 442294 597456 442350
rect 597512 442294 597580 442350
rect 597636 442294 597704 442350
rect 597760 442294 597828 442350
rect 597884 442294 597980 442350
rect 597360 442226 597980 442294
rect 597360 442170 597456 442226
rect 597512 442170 597580 442226
rect 597636 442170 597704 442226
rect 597760 442170 597828 442226
rect 597884 442170 597980 442226
rect 597360 442102 597980 442170
rect 597360 442046 597456 442102
rect 597512 442046 597580 442102
rect 597636 442046 597704 442102
rect 597760 442046 597828 442102
rect 597884 442046 597980 442102
rect 597360 441978 597980 442046
rect 597360 441922 597456 441978
rect 597512 441922 597580 441978
rect 597636 441922 597704 441978
rect 597760 441922 597828 441978
rect 597884 441922 597980 441978
rect 597360 424350 597980 441922
rect 597360 424294 597456 424350
rect 597512 424294 597580 424350
rect 597636 424294 597704 424350
rect 597760 424294 597828 424350
rect 597884 424294 597980 424350
rect 597360 424226 597980 424294
rect 597360 424170 597456 424226
rect 597512 424170 597580 424226
rect 597636 424170 597704 424226
rect 597760 424170 597828 424226
rect 597884 424170 597980 424226
rect 597360 424102 597980 424170
rect 597360 424046 597456 424102
rect 597512 424046 597580 424102
rect 597636 424046 597704 424102
rect 597760 424046 597828 424102
rect 597884 424046 597980 424102
rect 597360 423978 597980 424046
rect 597360 423922 597456 423978
rect 597512 423922 597580 423978
rect 597636 423922 597704 423978
rect 597760 423922 597828 423978
rect 597884 423922 597980 423978
rect 597360 406350 597980 423922
rect 597360 406294 597456 406350
rect 597512 406294 597580 406350
rect 597636 406294 597704 406350
rect 597760 406294 597828 406350
rect 597884 406294 597980 406350
rect 597360 406226 597980 406294
rect 597360 406170 597456 406226
rect 597512 406170 597580 406226
rect 597636 406170 597704 406226
rect 597760 406170 597828 406226
rect 597884 406170 597980 406226
rect 597360 406102 597980 406170
rect 597360 406046 597456 406102
rect 597512 406046 597580 406102
rect 597636 406046 597704 406102
rect 597760 406046 597828 406102
rect 597884 406046 597980 406102
rect 597360 405978 597980 406046
rect 597360 405922 597456 405978
rect 597512 405922 597580 405978
rect 597636 405922 597704 405978
rect 597760 405922 597828 405978
rect 597884 405922 597980 405978
rect 597360 388350 597980 405922
rect 597360 388294 597456 388350
rect 597512 388294 597580 388350
rect 597636 388294 597704 388350
rect 597760 388294 597828 388350
rect 597884 388294 597980 388350
rect 597360 388226 597980 388294
rect 597360 388170 597456 388226
rect 597512 388170 597580 388226
rect 597636 388170 597704 388226
rect 597760 388170 597828 388226
rect 597884 388170 597980 388226
rect 597360 388102 597980 388170
rect 597360 388046 597456 388102
rect 597512 388046 597580 388102
rect 597636 388046 597704 388102
rect 597760 388046 597828 388102
rect 597884 388046 597980 388102
rect 597360 387978 597980 388046
rect 597360 387922 597456 387978
rect 597512 387922 597580 387978
rect 597636 387922 597704 387978
rect 597760 387922 597828 387978
rect 597884 387922 597980 387978
rect 597360 370350 597980 387922
rect 597360 370294 597456 370350
rect 597512 370294 597580 370350
rect 597636 370294 597704 370350
rect 597760 370294 597828 370350
rect 597884 370294 597980 370350
rect 597360 370226 597980 370294
rect 597360 370170 597456 370226
rect 597512 370170 597580 370226
rect 597636 370170 597704 370226
rect 597760 370170 597828 370226
rect 597884 370170 597980 370226
rect 597360 370102 597980 370170
rect 597360 370046 597456 370102
rect 597512 370046 597580 370102
rect 597636 370046 597704 370102
rect 597760 370046 597828 370102
rect 597884 370046 597980 370102
rect 597360 369978 597980 370046
rect 597360 369922 597456 369978
rect 597512 369922 597580 369978
rect 597636 369922 597704 369978
rect 597760 369922 597828 369978
rect 597884 369922 597980 369978
rect 597360 352350 597980 369922
rect 597360 352294 597456 352350
rect 597512 352294 597580 352350
rect 597636 352294 597704 352350
rect 597760 352294 597828 352350
rect 597884 352294 597980 352350
rect 597360 352226 597980 352294
rect 597360 352170 597456 352226
rect 597512 352170 597580 352226
rect 597636 352170 597704 352226
rect 597760 352170 597828 352226
rect 597884 352170 597980 352226
rect 597360 352102 597980 352170
rect 597360 352046 597456 352102
rect 597512 352046 597580 352102
rect 597636 352046 597704 352102
rect 597760 352046 597828 352102
rect 597884 352046 597980 352102
rect 597360 351978 597980 352046
rect 597360 351922 597456 351978
rect 597512 351922 597580 351978
rect 597636 351922 597704 351978
rect 597760 351922 597828 351978
rect 597884 351922 597980 351978
rect 597360 334350 597980 351922
rect 597360 334294 597456 334350
rect 597512 334294 597580 334350
rect 597636 334294 597704 334350
rect 597760 334294 597828 334350
rect 597884 334294 597980 334350
rect 597360 334226 597980 334294
rect 597360 334170 597456 334226
rect 597512 334170 597580 334226
rect 597636 334170 597704 334226
rect 597760 334170 597828 334226
rect 597884 334170 597980 334226
rect 597360 334102 597980 334170
rect 597360 334046 597456 334102
rect 597512 334046 597580 334102
rect 597636 334046 597704 334102
rect 597760 334046 597828 334102
rect 597884 334046 597980 334102
rect 597360 333978 597980 334046
rect 597360 333922 597456 333978
rect 597512 333922 597580 333978
rect 597636 333922 597704 333978
rect 597760 333922 597828 333978
rect 597884 333922 597980 333978
rect 597360 316350 597980 333922
rect 597360 316294 597456 316350
rect 597512 316294 597580 316350
rect 597636 316294 597704 316350
rect 597760 316294 597828 316350
rect 597884 316294 597980 316350
rect 597360 316226 597980 316294
rect 597360 316170 597456 316226
rect 597512 316170 597580 316226
rect 597636 316170 597704 316226
rect 597760 316170 597828 316226
rect 597884 316170 597980 316226
rect 597360 316102 597980 316170
rect 597360 316046 597456 316102
rect 597512 316046 597580 316102
rect 597636 316046 597704 316102
rect 597760 316046 597828 316102
rect 597884 316046 597980 316102
rect 597360 315978 597980 316046
rect 597360 315922 597456 315978
rect 597512 315922 597580 315978
rect 597636 315922 597704 315978
rect 597760 315922 597828 315978
rect 597884 315922 597980 315978
rect 597360 298350 597980 315922
rect 597360 298294 597456 298350
rect 597512 298294 597580 298350
rect 597636 298294 597704 298350
rect 597760 298294 597828 298350
rect 597884 298294 597980 298350
rect 597360 298226 597980 298294
rect 597360 298170 597456 298226
rect 597512 298170 597580 298226
rect 597636 298170 597704 298226
rect 597760 298170 597828 298226
rect 597884 298170 597980 298226
rect 597360 298102 597980 298170
rect 597360 298046 597456 298102
rect 597512 298046 597580 298102
rect 597636 298046 597704 298102
rect 597760 298046 597828 298102
rect 597884 298046 597980 298102
rect 597360 297978 597980 298046
rect 597360 297922 597456 297978
rect 597512 297922 597580 297978
rect 597636 297922 597704 297978
rect 597760 297922 597828 297978
rect 597884 297922 597980 297978
rect 597360 280350 597980 297922
rect 597360 280294 597456 280350
rect 597512 280294 597580 280350
rect 597636 280294 597704 280350
rect 597760 280294 597828 280350
rect 597884 280294 597980 280350
rect 597360 280226 597980 280294
rect 597360 280170 597456 280226
rect 597512 280170 597580 280226
rect 597636 280170 597704 280226
rect 597760 280170 597828 280226
rect 597884 280170 597980 280226
rect 597360 280102 597980 280170
rect 597360 280046 597456 280102
rect 597512 280046 597580 280102
rect 597636 280046 597704 280102
rect 597760 280046 597828 280102
rect 597884 280046 597980 280102
rect 597360 279978 597980 280046
rect 597360 279922 597456 279978
rect 597512 279922 597580 279978
rect 597636 279922 597704 279978
rect 597760 279922 597828 279978
rect 597884 279922 597980 279978
rect 597360 262350 597980 279922
rect 597360 262294 597456 262350
rect 597512 262294 597580 262350
rect 597636 262294 597704 262350
rect 597760 262294 597828 262350
rect 597884 262294 597980 262350
rect 597360 262226 597980 262294
rect 597360 262170 597456 262226
rect 597512 262170 597580 262226
rect 597636 262170 597704 262226
rect 597760 262170 597828 262226
rect 597884 262170 597980 262226
rect 597360 262102 597980 262170
rect 597360 262046 597456 262102
rect 597512 262046 597580 262102
rect 597636 262046 597704 262102
rect 597760 262046 597828 262102
rect 597884 262046 597980 262102
rect 597360 261978 597980 262046
rect 597360 261922 597456 261978
rect 597512 261922 597580 261978
rect 597636 261922 597704 261978
rect 597760 261922 597828 261978
rect 597884 261922 597980 261978
rect 597360 244350 597980 261922
rect 597360 244294 597456 244350
rect 597512 244294 597580 244350
rect 597636 244294 597704 244350
rect 597760 244294 597828 244350
rect 597884 244294 597980 244350
rect 597360 244226 597980 244294
rect 597360 244170 597456 244226
rect 597512 244170 597580 244226
rect 597636 244170 597704 244226
rect 597760 244170 597828 244226
rect 597884 244170 597980 244226
rect 597360 244102 597980 244170
rect 597360 244046 597456 244102
rect 597512 244046 597580 244102
rect 597636 244046 597704 244102
rect 597760 244046 597828 244102
rect 597884 244046 597980 244102
rect 597360 243978 597980 244046
rect 597360 243922 597456 243978
rect 597512 243922 597580 243978
rect 597636 243922 597704 243978
rect 597760 243922 597828 243978
rect 597884 243922 597980 243978
rect 597360 226350 597980 243922
rect 597360 226294 597456 226350
rect 597512 226294 597580 226350
rect 597636 226294 597704 226350
rect 597760 226294 597828 226350
rect 597884 226294 597980 226350
rect 597360 226226 597980 226294
rect 597360 226170 597456 226226
rect 597512 226170 597580 226226
rect 597636 226170 597704 226226
rect 597760 226170 597828 226226
rect 597884 226170 597980 226226
rect 597360 226102 597980 226170
rect 597360 226046 597456 226102
rect 597512 226046 597580 226102
rect 597636 226046 597704 226102
rect 597760 226046 597828 226102
rect 597884 226046 597980 226102
rect 597360 225978 597980 226046
rect 597360 225922 597456 225978
rect 597512 225922 597580 225978
rect 597636 225922 597704 225978
rect 597760 225922 597828 225978
rect 597884 225922 597980 225978
rect 597360 208350 597980 225922
rect 597360 208294 597456 208350
rect 597512 208294 597580 208350
rect 597636 208294 597704 208350
rect 597760 208294 597828 208350
rect 597884 208294 597980 208350
rect 597360 208226 597980 208294
rect 597360 208170 597456 208226
rect 597512 208170 597580 208226
rect 597636 208170 597704 208226
rect 597760 208170 597828 208226
rect 597884 208170 597980 208226
rect 597360 208102 597980 208170
rect 597360 208046 597456 208102
rect 597512 208046 597580 208102
rect 597636 208046 597704 208102
rect 597760 208046 597828 208102
rect 597884 208046 597980 208102
rect 597360 207978 597980 208046
rect 597360 207922 597456 207978
rect 597512 207922 597580 207978
rect 597636 207922 597704 207978
rect 597760 207922 597828 207978
rect 597884 207922 597980 207978
rect 597360 190350 597980 207922
rect 597360 190294 597456 190350
rect 597512 190294 597580 190350
rect 597636 190294 597704 190350
rect 597760 190294 597828 190350
rect 597884 190294 597980 190350
rect 597360 190226 597980 190294
rect 597360 190170 597456 190226
rect 597512 190170 597580 190226
rect 597636 190170 597704 190226
rect 597760 190170 597828 190226
rect 597884 190170 597980 190226
rect 597360 190102 597980 190170
rect 597360 190046 597456 190102
rect 597512 190046 597580 190102
rect 597636 190046 597704 190102
rect 597760 190046 597828 190102
rect 597884 190046 597980 190102
rect 597360 189978 597980 190046
rect 597360 189922 597456 189978
rect 597512 189922 597580 189978
rect 597636 189922 597704 189978
rect 597760 189922 597828 189978
rect 597884 189922 597980 189978
rect 597360 172350 597980 189922
rect 597360 172294 597456 172350
rect 597512 172294 597580 172350
rect 597636 172294 597704 172350
rect 597760 172294 597828 172350
rect 597884 172294 597980 172350
rect 597360 172226 597980 172294
rect 597360 172170 597456 172226
rect 597512 172170 597580 172226
rect 597636 172170 597704 172226
rect 597760 172170 597828 172226
rect 597884 172170 597980 172226
rect 597360 172102 597980 172170
rect 597360 172046 597456 172102
rect 597512 172046 597580 172102
rect 597636 172046 597704 172102
rect 597760 172046 597828 172102
rect 597884 172046 597980 172102
rect 597360 171978 597980 172046
rect 597360 171922 597456 171978
rect 597512 171922 597580 171978
rect 597636 171922 597704 171978
rect 597760 171922 597828 171978
rect 597884 171922 597980 171978
rect 597360 154350 597980 171922
rect 597360 154294 597456 154350
rect 597512 154294 597580 154350
rect 597636 154294 597704 154350
rect 597760 154294 597828 154350
rect 597884 154294 597980 154350
rect 597360 154226 597980 154294
rect 597360 154170 597456 154226
rect 597512 154170 597580 154226
rect 597636 154170 597704 154226
rect 597760 154170 597828 154226
rect 597884 154170 597980 154226
rect 597360 154102 597980 154170
rect 597360 154046 597456 154102
rect 597512 154046 597580 154102
rect 597636 154046 597704 154102
rect 597760 154046 597828 154102
rect 597884 154046 597980 154102
rect 597360 153978 597980 154046
rect 597360 153922 597456 153978
rect 597512 153922 597580 153978
rect 597636 153922 597704 153978
rect 597760 153922 597828 153978
rect 597884 153922 597980 153978
rect 597360 136350 597980 153922
rect 597360 136294 597456 136350
rect 597512 136294 597580 136350
rect 597636 136294 597704 136350
rect 597760 136294 597828 136350
rect 597884 136294 597980 136350
rect 597360 136226 597980 136294
rect 597360 136170 597456 136226
rect 597512 136170 597580 136226
rect 597636 136170 597704 136226
rect 597760 136170 597828 136226
rect 597884 136170 597980 136226
rect 597360 136102 597980 136170
rect 597360 136046 597456 136102
rect 597512 136046 597580 136102
rect 597636 136046 597704 136102
rect 597760 136046 597828 136102
rect 597884 136046 597980 136102
rect 597360 135978 597980 136046
rect 597360 135922 597456 135978
rect 597512 135922 597580 135978
rect 597636 135922 597704 135978
rect 597760 135922 597828 135978
rect 597884 135922 597980 135978
rect 597360 118350 597980 135922
rect 597360 118294 597456 118350
rect 597512 118294 597580 118350
rect 597636 118294 597704 118350
rect 597760 118294 597828 118350
rect 597884 118294 597980 118350
rect 597360 118226 597980 118294
rect 597360 118170 597456 118226
rect 597512 118170 597580 118226
rect 597636 118170 597704 118226
rect 597760 118170 597828 118226
rect 597884 118170 597980 118226
rect 597360 118102 597980 118170
rect 597360 118046 597456 118102
rect 597512 118046 597580 118102
rect 597636 118046 597704 118102
rect 597760 118046 597828 118102
rect 597884 118046 597980 118102
rect 597360 117978 597980 118046
rect 597360 117922 597456 117978
rect 597512 117922 597580 117978
rect 597636 117922 597704 117978
rect 597760 117922 597828 117978
rect 597884 117922 597980 117978
rect 597360 100350 597980 117922
rect 597360 100294 597456 100350
rect 597512 100294 597580 100350
rect 597636 100294 597704 100350
rect 597760 100294 597828 100350
rect 597884 100294 597980 100350
rect 597360 100226 597980 100294
rect 597360 100170 597456 100226
rect 597512 100170 597580 100226
rect 597636 100170 597704 100226
rect 597760 100170 597828 100226
rect 597884 100170 597980 100226
rect 597360 100102 597980 100170
rect 597360 100046 597456 100102
rect 597512 100046 597580 100102
rect 597636 100046 597704 100102
rect 597760 100046 597828 100102
rect 597884 100046 597980 100102
rect 597360 99978 597980 100046
rect 597360 99922 597456 99978
rect 597512 99922 597580 99978
rect 597636 99922 597704 99978
rect 597760 99922 597828 99978
rect 597884 99922 597980 99978
rect 597360 82350 597980 99922
rect 597360 82294 597456 82350
rect 597512 82294 597580 82350
rect 597636 82294 597704 82350
rect 597760 82294 597828 82350
rect 597884 82294 597980 82350
rect 597360 82226 597980 82294
rect 597360 82170 597456 82226
rect 597512 82170 597580 82226
rect 597636 82170 597704 82226
rect 597760 82170 597828 82226
rect 597884 82170 597980 82226
rect 597360 82102 597980 82170
rect 597360 82046 597456 82102
rect 597512 82046 597580 82102
rect 597636 82046 597704 82102
rect 597760 82046 597828 82102
rect 597884 82046 597980 82102
rect 597360 81978 597980 82046
rect 597360 81922 597456 81978
rect 597512 81922 597580 81978
rect 597636 81922 597704 81978
rect 597760 81922 597828 81978
rect 597884 81922 597980 81978
rect 597360 64350 597980 81922
rect 597360 64294 597456 64350
rect 597512 64294 597580 64350
rect 597636 64294 597704 64350
rect 597760 64294 597828 64350
rect 597884 64294 597980 64350
rect 597360 64226 597980 64294
rect 597360 64170 597456 64226
rect 597512 64170 597580 64226
rect 597636 64170 597704 64226
rect 597760 64170 597828 64226
rect 597884 64170 597980 64226
rect 597360 64102 597980 64170
rect 597360 64046 597456 64102
rect 597512 64046 597580 64102
rect 597636 64046 597704 64102
rect 597760 64046 597828 64102
rect 597884 64046 597980 64102
rect 597360 63978 597980 64046
rect 597360 63922 597456 63978
rect 597512 63922 597580 63978
rect 597636 63922 597704 63978
rect 597760 63922 597828 63978
rect 597884 63922 597980 63978
rect 597360 46350 597980 63922
rect 597360 46294 597456 46350
rect 597512 46294 597580 46350
rect 597636 46294 597704 46350
rect 597760 46294 597828 46350
rect 597884 46294 597980 46350
rect 597360 46226 597980 46294
rect 597360 46170 597456 46226
rect 597512 46170 597580 46226
rect 597636 46170 597704 46226
rect 597760 46170 597828 46226
rect 597884 46170 597980 46226
rect 597360 46102 597980 46170
rect 597360 46046 597456 46102
rect 597512 46046 597580 46102
rect 597636 46046 597704 46102
rect 597760 46046 597828 46102
rect 597884 46046 597980 46102
rect 597360 45978 597980 46046
rect 597360 45922 597456 45978
rect 597512 45922 597580 45978
rect 597636 45922 597704 45978
rect 597760 45922 597828 45978
rect 597884 45922 597980 45978
rect 597360 28350 597980 45922
rect 597360 28294 597456 28350
rect 597512 28294 597580 28350
rect 597636 28294 597704 28350
rect 597760 28294 597828 28350
rect 597884 28294 597980 28350
rect 597360 28226 597980 28294
rect 597360 28170 597456 28226
rect 597512 28170 597580 28226
rect 597636 28170 597704 28226
rect 597760 28170 597828 28226
rect 597884 28170 597980 28226
rect 597360 28102 597980 28170
rect 597360 28046 597456 28102
rect 597512 28046 597580 28102
rect 597636 28046 597704 28102
rect 597760 28046 597828 28102
rect 597884 28046 597980 28102
rect 597360 27978 597980 28046
rect 597360 27922 597456 27978
rect 597512 27922 597580 27978
rect 597636 27922 597704 27978
rect 597760 27922 597828 27978
rect 597884 27922 597980 27978
rect 597360 10350 597980 27922
rect 597360 10294 597456 10350
rect 597512 10294 597580 10350
rect 597636 10294 597704 10350
rect 597760 10294 597828 10350
rect 597884 10294 597980 10350
rect 597360 10226 597980 10294
rect 597360 10170 597456 10226
rect 597512 10170 597580 10226
rect 597636 10170 597704 10226
rect 597760 10170 597828 10226
rect 597884 10170 597980 10226
rect 597360 10102 597980 10170
rect 597360 10046 597456 10102
rect 597512 10046 597580 10102
rect 597636 10046 597704 10102
rect 597760 10046 597828 10102
rect 597884 10046 597980 10102
rect 597360 9978 597980 10046
rect 597360 9922 597456 9978
rect 597512 9922 597580 9978
rect 597636 9922 597704 9978
rect 597760 9922 597828 9978
rect 597884 9922 597980 9978
rect 582874 -1176 582970 -1120
rect 583026 -1176 583094 -1120
rect 583150 -1176 583218 -1120
rect 583274 -1176 583342 -1120
rect 583398 -1176 583494 -1120
rect 582874 -1244 583494 -1176
rect 582874 -1300 582970 -1244
rect 583026 -1300 583094 -1244
rect 583150 -1300 583218 -1244
rect 583274 -1300 583342 -1244
rect 583398 -1300 583494 -1244
rect 582874 -1368 583494 -1300
rect 582874 -1424 582970 -1368
rect 583026 -1424 583094 -1368
rect 583150 -1424 583218 -1368
rect 583274 -1424 583342 -1368
rect 583398 -1424 583494 -1368
rect 582874 -1492 583494 -1424
rect 582874 -1548 582970 -1492
rect 583026 -1548 583094 -1492
rect 583150 -1548 583218 -1492
rect 583274 -1548 583342 -1492
rect 583398 -1548 583494 -1492
rect 582874 -1644 583494 -1548
rect 597360 -1120 597980 9922
rect 597360 -1176 597456 -1120
rect 597512 -1176 597580 -1120
rect 597636 -1176 597704 -1120
rect 597760 -1176 597828 -1120
rect 597884 -1176 597980 -1120
rect 597360 -1244 597980 -1176
rect 597360 -1300 597456 -1244
rect 597512 -1300 597580 -1244
rect 597636 -1300 597704 -1244
rect 597760 -1300 597828 -1244
rect 597884 -1300 597980 -1244
rect 597360 -1368 597980 -1300
rect 597360 -1424 597456 -1368
rect 597512 -1424 597580 -1368
rect 597636 -1424 597704 -1368
rect 597760 -1424 597828 -1368
rect 597884 -1424 597980 -1368
rect 597360 -1492 597980 -1424
rect 597360 -1548 597456 -1492
rect 597512 -1548 597580 -1492
rect 597636 -1548 597704 -1492
rect 597760 -1548 597828 -1492
rect 597884 -1548 597980 -1492
rect 597360 -1644 597980 -1548
<< via4 >>
rect -1820 598116 -1764 598172
rect -1696 598116 -1640 598172
rect -1572 598116 -1516 598172
rect -1448 598116 -1392 598172
rect -1820 597992 -1764 598048
rect -1696 597992 -1640 598048
rect -1572 597992 -1516 598048
rect -1448 597992 -1392 598048
rect -1820 597868 -1764 597924
rect -1696 597868 -1640 597924
rect -1572 597868 -1516 597924
rect -1448 597868 -1392 597924
rect -1820 597744 -1764 597800
rect -1696 597744 -1640 597800
rect -1572 597744 -1516 597800
rect -1448 597744 -1392 597800
rect -1820 586294 -1764 586350
rect -1696 586294 -1640 586350
rect -1572 586294 -1516 586350
rect -1448 586294 -1392 586350
rect -1820 586170 -1764 586226
rect -1696 586170 -1640 586226
rect -1572 586170 -1516 586226
rect -1448 586170 -1392 586226
rect -1820 586046 -1764 586102
rect -1696 586046 -1640 586102
rect -1572 586046 -1516 586102
rect -1448 586046 -1392 586102
rect -1820 585922 -1764 585978
rect -1696 585922 -1640 585978
rect -1572 585922 -1516 585978
rect -1448 585922 -1392 585978
rect -1820 568294 -1764 568350
rect -1696 568294 -1640 568350
rect -1572 568294 -1516 568350
rect -1448 568294 -1392 568350
rect -1820 568170 -1764 568226
rect -1696 568170 -1640 568226
rect -1572 568170 -1516 568226
rect -1448 568170 -1392 568226
rect -1820 568046 -1764 568102
rect -1696 568046 -1640 568102
rect -1572 568046 -1516 568102
rect -1448 568046 -1392 568102
rect -1820 567922 -1764 567978
rect -1696 567922 -1640 567978
rect -1572 567922 -1516 567978
rect -1448 567922 -1392 567978
rect -1820 550294 -1764 550350
rect -1696 550294 -1640 550350
rect -1572 550294 -1516 550350
rect -1448 550294 -1392 550350
rect -1820 550170 -1764 550226
rect -1696 550170 -1640 550226
rect -1572 550170 -1516 550226
rect -1448 550170 -1392 550226
rect -1820 550046 -1764 550102
rect -1696 550046 -1640 550102
rect -1572 550046 -1516 550102
rect -1448 550046 -1392 550102
rect -1820 549922 -1764 549978
rect -1696 549922 -1640 549978
rect -1572 549922 -1516 549978
rect -1448 549922 -1392 549978
rect -1820 532294 -1764 532350
rect -1696 532294 -1640 532350
rect -1572 532294 -1516 532350
rect -1448 532294 -1392 532350
rect -1820 532170 -1764 532226
rect -1696 532170 -1640 532226
rect -1572 532170 -1516 532226
rect -1448 532170 -1392 532226
rect -1820 532046 -1764 532102
rect -1696 532046 -1640 532102
rect -1572 532046 -1516 532102
rect -1448 532046 -1392 532102
rect -1820 531922 -1764 531978
rect -1696 531922 -1640 531978
rect -1572 531922 -1516 531978
rect -1448 531922 -1392 531978
rect -1820 514294 -1764 514350
rect -1696 514294 -1640 514350
rect -1572 514294 -1516 514350
rect -1448 514294 -1392 514350
rect -1820 514170 -1764 514226
rect -1696 514170 -1640 514226
rect -1572 514170 -1516 514226
rect -1448 514170 -1392 514226
rect -1820 514046 -1764 514102
rect -1696 514046 -1640 514102
rect -1572 514046 -1516 514102
rect -1448 514046 -1392 514102
rect -1820 513922 -1764 513978
rect -1696 513922 -1640 513978
rect -1572 513922 -1516 513978
rect -1448 513922 -1392 513978
rect -1820 496294 -1764 496350
rect -1696 496294 -1640 496350
rect -1572 496294 -1516 496350
rect -1448 496294 -1392 496350
rect -1820 496170 -1764 496226
rect -1696 496170 -1640 496226
rect -1572 496170 -1516 496226
rect -1448 496170 -1392 496226
rect -1820 496046 -1764 496102
rect -1696 496046 -1640 496102
rect -1572 496046 -1516 496102
rect -1448 496046 -1392 496102
rect -1820 495922 -1764 495978
rect -1696 495922 -1640 495978
rect -1572 495922 -1516 495978
rect -1448 495922 -1392 495978
rect -1820 478294 -1764 478350
rect -1696 478294 -1640 478350
rect -1572 478294 -1516 478350
rect -1448 478294 -1392 478350
rect -1820 478170 -1764 478226
rect -1696 478170 -1640 478226
rect -1572 478170 -1516 478226
rect -1448 478170 -1392 478226
rect -1820 478046 -1764 478102
rect -1696 478046 -1640 478102
rect -1572 478046 -1516 478102
rect -1448 478046 -1392 478102
rect -1820 477922 -1764 477978
rect -1696 477922 -1640 477978
rect -1572 477922 -1516 477978
rect -1448 477922 -1392 477978
rect -1820 460294 -1764 460350
rect -1696 460294 -1640 460350
rect -1572 460294 -1516 460350
rect -1448 460294 -1392 460350
rect -1820 460170 -1764 460226
rect -1696 460170 -1640 460226
rect -1572 460170 -1516 460226
rect -1448 460170 -1392 460226
rect -1820 460046 -1764 460102
rect -1696 460046 -1640 460102
rect -1572 460046 -1516 460102
rect -1448 460046 -1392 460102
rect -1820 459922 -1764 459978
rect -1696 459922 -1640 459978
rect -1572 459922 -1516 459978
rect -1448 459922 -1392 459978
rect -1820 442294 -1764 442350
rect -1696 442294 -1640 442350
rect -1572 442294 -1516 442350
rect -1448 442294 -1392 442350
rect -1820 442170 -1764 442226
rect -1696 442170 -1640 442226
rect -1572 442170 -1516 442226
rect -1448 442170 -1392 442226
rect -1820 442046 -1764 442102
rect -1696 442046 -1640 442102
rect -1572 442046 -1516 442102
rect -1448 442046 -1392 442102
rect -1820 441922 -1764 441978
rect -1696 441922 -1640 441978
rect -1572 441922 -1516 441978
rect -1448 441922 -1392 441978
rect -1820 424294 -1764 424350
rect -1696 424294 -1640 424350
rect -1572 424294 -1516 424350
rect -1448 424294 -1392 424350
rect -1820 424170 -1764 424226
rect -1696 424170 -1640 424226
rect -1572 424170 -1516 424226
rect -1448 424170 -1392 424226
rect -1820 424046 -1764 424102
rect -1696 424046 -1640 424102
rect -1572 424046 -1516 424102
rect -1448 424046 -1392 424102
rect -1820 423922 -1764 423978
rect -1696 423922 -1640 423978
rect -1572 423922 -1516 423978
rect -1448 423922 -1392 423978
rect -1820 406294 -1764 406350
rect -1696 406294 -1640 406350
rect -1572 406294 -1516 406350
rect -1448 406294 -1392 406350
rect -1820 406170 -1764 406226
rect -1696 406170 -1640 406226
rect -1572 406170 -1516 406226
rect -1448 406170 -1392 406226
rect -1820 406046 -1764 406102
rect -1696 406046 -1640 406102
rect -1572 406046 -1516 406102
rect -1448 406046 -1392 406102
rect -1820 405922 -1764 405978
rect -1696 405922 -1640 405978
rect -1572 405922 -1516 405978
rect -1448 405922 -1392 405978
rect -1820 388294 -1764 388350
rect -1696 388294 -1640 388350
rect -1572 388294 -1516 388350
rect -1448 388294 -1392 388350
rect -1820 388170 -1764 388226
rect -1696 388170 -1640 388226
rect -1572 388170 -1516 388226
rect -1448 388170 -1392 388226
rect -1820 388046 -1764 388102
rect -1696 388046 -1640 388102
rect -1572 388046 -1516 388102
rect -1448 388046 -1392 388102
rect -1820 387922 -1764 387978
rect -1696 387922 -1640 387978
rect -1572 387922 -1516 387978
rect -1448 387922 -1392 387978
rect -1820 370294 -1764 370350
rect -1696 370294 -1640 370350
rect -1572 370294 -1516 370350
rect -1448 370294 -1392 370350
rect -1820 370170 -1764 370226
rect -1696 370170 -1640 370226
rect -1572 370170 -1516 370226
rect -1448 370170 -1392 370226
rect -1820 370046 -1764 370102
rect -1696 370046 -1640 370102
rect -1572 370046 -1516 370102
rect -1448 370046 -1392 370102
rect -1820 369922 -1764 369978
rect -1696 369922 -1640 369978
rect -1572 369922 -1516 369978
rect -1448 369922 -1392 369978
rect -1820 352294 -1764 352350
rect -1696 352294 -1640 352350
rect -1572 352294 -1516 352350
rect -1448 352294 -1392 352350
rect -1820 352170 -1764 352226
rect -1696 352170 -1640 352226
rect -1572 352170 -1516 352226
rect -1448 352170 -1392 352226
rect -1820 352046 -1764 352102
rect -1696 352046 -1640 352102
rect -1572 352046 -1516 352102
rect -1448 352046 -1392 352102
rect -1820 351922 -1764 351978
rect -1696 351922 -1640 351978
rect -1572 351922 -1516 351978
rect -1448 351922 -1392 351978
rect -1820 334294 -1764 334350
rect -1696 334294 -1640 334350
rect -1572 334294 -1516 334350
rect -1448 334294 -1392 334350
rect -1820 334170 -1764 334226
rect -1696 334170 -1640 334226
rect -1572 334170 -1516 334226
rect -1448 334170 -1392 334226
rect -1820 334046 -1764 334102
rect -1696 334046 -1640 334102
rect -1572 334046 -1516 334102
rect -1448 334046 -1392 334102
rect -1820 333922 -1764 333978
rect -1696 333922 -1640 333978
rect -1572 333922 -1516 333978
rect -1448 333922 -1392 333978
rect -1820 316294 -1764 316350
rect -1696 316294 -1640 316350
rect -1572 316294 -1516 316350
rect -1448 316294 -1392 316350
rect -1820 316170 -1764 316226
rect -1696 316170 -1640 316226
rect -1572 316170 -1516 316226
rect -1448 316170 -1392 316226
rect -1820 316046 -1764 316102
rect -1696 316046 -1640 316102
rect -1572 316046 -1516 316102
rect -1448 316046 -1392 316102
rect -1820 315922 -1764 315978
rect -1696 315922 -1640 315978
rect -1572 315922 -1516 315978
rect -1448 315922 -1392 315978
rect -1820 298294 -1764 298350
rect -1696 298294 -1640 298350
rect -1572 298294 -1516 298350
rect -1448 298294 -1392 298350
rect -1820 298170 -1764 298226
rect -1696 298170 -1640 298226
rect -1572 298170 -1516 298226
rect -1448 298170 -1392 298226
rect -1820 298046 -1764 298102
rect -1696 298046 -1640 298102
rect -1572 298046 -1516 298102
rect -1448 298046 -1392 298102
rect -1820 297922 -1764 297978
rect -1696 297922 -1640 297978
rect -1572 297922 -1516 297978
rect -1448 297922 -1392 297978
rect -1820 280294 -1764 280350
rect -1696 280294 -1640 280350
rect -1572 280294 -1516 280350
rect -1448 280294 -1392 280350
rect -1820 280170 -1764 280226
rect -1696 280170 -1640 280226
rect -1572 280170 -1516 280226
rect -1448 280170 -1392 280226
rect -1820 280046 -1764 280102
rect -1696 280046 -1640 280102
rect -1572 280046 -1516 280102
rect -1448 280046 -1392 280102
rect -1820 279922 -1764 279978
rect -1696 279922 -1640 279978
rect -1572 279922 -1516 279978
rect -1448 279922 -1392 279978
rect -1820 262294 -1764 262350
rect -1696 262294 -1640 262350
rect -1572 262294 -1516 262350
rect -1448 262294 -1392 262350
rect -1820 262170 -1764 262226
rect -1696 262170 -1640 262226
rect -1572 262170 -1516 262226
rect -1448 262170 -1392 262226
rect -1820 262046 -1764 262102
rect -1696 262046 -1640 262102
rect -1572 262046 -1516 262102
rect -1448 262046 -1392 262102
rect -1820 261922 -1764 261978
rect -1696 261922 -1640 261978
rect -1572 261922 -1516 261978
rect -1448 261922 -1392 261978
rect -1820 244294 -1764 244350
rect -1696 244294 -1640 244350
rect -1572 244294 -1516 244350
rect -1448 244294 -1392 244350
rect -1820 244170 -1764 244226
rect -1696 244170 -1640 244226
rect -1572 244170 -1516 244226
rect -1448 244170 -1392 244226
rect -1820 244046 -1764 244102
rect -1696 244046 -1640 244102
rect -1572 244046 -1516 244102
rect -1448 244046 -1392 244102
rect -1820 243922 -1764 243978
rect -1696 243922 -1640 243978
rect -1572 243922 -1516 243978
rect -1448 243922 -1392 243978
rect -1820 226294 -1764 226350
rect -1696 226294 -1640 226350
rect -1572 226294 -1516 226350
rect -1448 226294 -1392 226350
rect -1820 226170 -1764 226226
rect -1696 226170 -1640 226226
rect -1572 226170 -1516 226226
rect -1448 226170 -1392 226226
rect -1820 226046 -1764 226102
rect -1696 226046 -1640 226102
rect -1572 226046 -1516 226102
rect -1448 226046 -1392 226102
rect -1820 225922 -1764 225978
rect -1696 225922 -1640 225978
rect -1572 225922 -1516 225978
rect -1448 225922 -1392 225978
rect -1820 208294 -1764 208350
rect -1696 208294 -1640 208350
rect -1572 208294 -1516 208350
rect -1448 208294 -1392 208350
rect -1820 208170 -1764 208226
rect -1696 208170 -1640 208226
rect -1572 208170 -1516 208226
rect -1448 208170 -1392 208226
rect -1820 208046 -1764 208102
rect -1696 208046 -1640 208102
rect -1572 208046 -1516 208102
rect -1448 208046 -1392 208102
rect -1820 207922 -1764 207978
rect -1696 207922 -1640 207978
rect -1572 207922 -1516 207978
rect -1448 207922 -1392 207978
rect -1820 190294 -1764 190350
rect -1696 190294 -1640 190350
rect -1572 190294 -1516 190350
rect -1448 190294 -1392 190350
rect -1820 190170 -1764 190226
rect -1696 190170 -1640 190226
rect -1572 190170 -1516 190226
rect -1448 190170 -1392 190226
rect -1820 190046 -1764 190102
rect -1696 190046 -1640 190102
rect -1572 190046 -1516 190102
rect -1448 190046 -1392 190102
rect -1820 189922 -1764 189978
rect -1696 189922 -1640 189978
rect -1572 189922 -1516 189978
rect -1448 189922 -1392 189978
rect -1820 172294 -1764 172350
rect -1696 172294 -1640 172350
rect -1572 172294 -1516 172350
rect -1448 172294 -1392 172350
rect -1820 172170 -1764 172226
rect -1696 172170 -1640 172226
rect -1572 172170 -1516 172226
rect -1448 172170 -1392 172226
rect -1820 172046 -1764 172102
rect -1696 172046 -1640 172102
rect -1572 172046 -1516 172102
rect -1448 172046 -1392 172102
rect -1820 171922 -1764 171978
rect -1696 171922 -1640 171978
rect -1572 171922 -1516 171978
rect -1448 171922 -1392 171978
rect -1820 154294 -1764 154350
rect -1696 154294 -1640 154350
rect -1572 154294 -1516 154350
rect -1448 154294 -1392 154350
rect -1820 154170 -1764 154226
rect -1696 154170 -1640 154226
rect -1572 154170 -1516 154226
rect -1448 154170 -1392 154226
rect -1820 154046 -1764 154102
rect -1696 154046 -1640 154102
rect -1572 154046 -1516 154102
rect -1448 154046 -1392 154102
rect -1820 153922 -1764 153978
rect -1696 153922 -1640 153978
rect -1572 153922 -1516 153978
rect -1448 153922 -1392 153978
rect -1820 136294 -1764 136350
rect -1696 136294 -1640 136350
rect -1572 136294 -1516 136350
rect -1448 136294 -1392 136350
rect -1820 136170 -1764 136226
rect -1696 136170 -1640 136226
rect -1572 136170 -1516 136226
rect -1448 136170 -1392 136226
rect -1820 136046 -1764 136102
rect -1696 136046 -1640 136102
rect -1572 136046 -1516 136102
rect -1448 136046 -1392 136102
rect -1820 135922 -1764 135978
rect -1696 135922 -1640 135978
rect -1572 135922 -1516 135978
rect -1448 135922 -1392 135978
rect -1820 118294 -1764 118350
rect -1696 118294 -1640 118350
rect -1572 118294 -1516 118350
rect -1448 118294 -1392 118350
rect -1820 118170 -1764 118226
rect -1696 118170 -1640 118226
rect -1572 118170 -1516 118226
rect -1448 118170 -1392 118226
rect -1820 118046 -1764 118102
rect -1696 118046 -1640 118102
rect -1572 118046 -1516 118102
rect -1448 118046 -1392 118102
rect -1820 117922 -1764 117978
rect -1696 117922 -1640 117978
rect -1572 117922 -1516 117978
rect -1448 117922 -1392 117978
rect -1820 100294 -1764 100350
rect -1696 100294 -1640 100350
rect -1572 100294 -1516 100350
rect -1448 100294 -1392 100350
rect -1820 100170 -1764 100226
rect -1696 100170 -1640 100226
rect -1572 100170 -1516 100226
rect -1448 100170 -1392 100226
rect -1820 100046 -1764 100102
rect -1696 100046 -1640 100102
rect -1572 100046 -1516 100102
rect -1448 100046 -1392 100102
rect -1820 99922 -1764 99978
rect -1696 99922 -1640 99978
rect -1572 99922 -1516 99978
rect -1448 99922 -1392 99978
rect -1820 82294 -1764 82350
rect -1696 82294 -1640 82350
rect -1572 82294 -1516 82350
rect -1448 82294 -1392 82350
rect -1820 82170 -1764 82226
rect -1696 82170 -1640 82226
rect -1572 82170 -1516 82226
rect -1448 82170 -1392 82226
rect -1820 82046 -1764 82102
rect -1696 82046 -1640 82102
rect -1572 82046 -1516 82102
rect -1448 82046 -1392 82102
rect -1820 81922 -1764 81978
rect -1696 81922 -1640 81978
rect -1572 81922 -1516 81978
rect -1448 81922 -1392 81978
rect -1820 64294 -1764 64350
rect -1696 64294 -1640 64350
rect -1572 64294 -1516 64350
rect -1448 64294 -1392 64350
rect -1820 64170 -1764 64226
rect -1696 64170 -1640 64226
rect -1572 64170 -1516 64226
rect -1448 64170 -1392 64226
rect -1820 64046 -1764 64102
rect -1696 64046 -1640 64102
rect -1572 64046 -1516 64102
rect -1448 64046 -1392 64102
rect -1820 63922 -1764 63978
rect -1696 63922 -1640 63978
rect -1572 63922 -1516 63978
rect -1448 63922 -1392 63978
rect -1820 46294 -1764 46350
rect -1696 46294 -1640 46350
rect -1572 46294 -1516 46350
rect -1448 46294 -1392 46350
rect -1820 46170 -1764 46226
rect -1696 46170 -1640 46226
rect -1572 46170 -1516 46226
rect -1448 46170 -1392 46226
rect -1820 46046 -1764 46102
rect -1696 46046 -1640 46102
rect -1572 46046 -1516 46102
rect -1448 46046 -1392 46102
rect -1820 45922 -1764 45978
rect -1696 45922 -1640 45978
rect -1572 45922 -1516 45978
rect -1448 45922 -1392 45978
rect -1820 28294 -1764 28350
rect -1696 28294 -1640 28350
rect -1572 28294 -1516 28350
rect -1448 28294 -1392 28350
rect -1820 28170 -1764 28226
rect -1696 28170 -1640 28226
rect -1572 28170 -1516 28226
rect -1448 28170 -1392 28226
rect -1820 28046 -1764 28102
rect -1696 28046 -1640 28102
rect -1572 28046 -1516 28102
rect -1448 28046 -1392 28102
rect -1820 27922 -1764 27978
rect -1696 27922 -1640 27978
rect -1572 27922 -1516 27978
rect -1448 27922 -1392 27978
rect -1820 10294 -1764 10350
rect -1696 10294 -1640 10350
rect -1572 10294 -1516 10350
rect -1448 10294 -1392 10350
rect -1820 10170 -1764 10226
rect -1696 10170 -1640 10226
rect -1572 10170 -1516 10226
rect -1448 10170 -1392 10226
rect -1820 10046 -1764 10102
rect -1696 10046 -1640 10102
rect -1572 10046 -1516 10102
rect -1448 10046 -1392 10102
rect -1820 9922 -1764 9978
rect -1696 9922 -1640 9978
rect -1572 9922 -1516 9978
rect -1448 9922 -1392 9978
rect -860 597156 -804 597212
rect -736 597156 -680 597212
rect -612 597156 -556 597212
rect -488 597156 -432 597212
rect -860 597032 -804 597088
rect -736 597032 -680 597088
rect -612 597032 -556 597088
rect -488 597032 -432 597088
rect -860 596908 -804 596964
rect -736 596908 -680 596964
rect -612 596908 -556 596964
rect -488 596908 -432 596964
rect -860 596784 -804 596840
rect -736 596784 -680 596840
rect -612 596784 -556 596840
rect -488 596784 -432 596840
rect -860 580294 -804 580350
rect -736 580294 -680 580350
rect -612 580294 -556 580350
rect -488 580294 -432 580350
rect -860 580170 -804 580226
rect -736 580170 -680 580226
rect -612 580170 -556 580226
rect -488 580170 -432 580226
rect -860 580046 -804 580102
rect -736 580046 -680 580102
rect -612 580046 -556 580102
rect -488 580046 -432 580102
rect -860 579922 -804 579978
rect -736 579922 -680 579978
rect -612 579922 -556 579978
rect -488 579922 -432 579978
rect -860 562294 -804 562350
rect -736 562294 -680 562350
rect -612 562294 -556 562350
rect -488 562294 -432 562350
rect -860 562170 -804 562226
rect -736 562170 -680 562226
rect -612 562170 -556 562226
rect -488 562170 -432 562226
rect -860 562046 -804 562102
rect -736 562046 -680 562102
rect -612 562046 -556 562102
rect -488 562046 -432 562102
rect -860 561922 -804 561978
rect -736 561922 -680 561978
rect -612 561922 -556 561978
rect -488 561922 -432 561978
rect -860 544294 -804 544350
rect -736 544294 -680 544350
rect -612 544294 -556 544350
rect -488 544294 -432 544350
rect -860 544170 -804 544226
rect -736 544170 -680 544226
rect -612 544170 -556 544226
rect -488 544170 -432 544226
rect -860 544046 -804 544102
rect -736 544046 -680 544102
rect -612 544046 -556 544102
rect -488 544046 -432 544102
rect -860 543922 -804 543978
rect -736 543922 -680 543978
rect -612 543922 -556 543978
rect -488 543922 -432 543978
rect -860 526294 -804 526350
rect -736 526294 -680 526350
rect -612 526294 -556 526350
rect -488 526294 -432 526350
rect -860 526170 -804 526226
rect -736 526170 -680 526226
rect -612 526170 -556 526226
rect -488 526170 -432 526226
rect -860 526046 -804 526102
rect -736 526046 -680 526102
rect -612 526046 -556 526102
rect -488 526046 -432 526102
rect -860 525922 -804 525978
rect -736 525922 -680 525978
rect -612 525922 -556 525978
rect -488 525922 -432 525978
rect -860 508294 -804 508350
rect -736 508294 -680 508350
rect -612 508294 -556 508350
rect -488 508294 -432 508350
rect -860 508170 -804 508226
rect -736 508170 -680 508226
rect -612 508170 -556 508226
rect -488 508170 -432 508226
rect -860 508046 -804 508102
rect -736 508046 -680 508102
rect -612 508046 -556 508102
rect -488 508046 -432 508102
rect -860 507922 -804 507978
rect -736 507922 -680 507978
rect -612 507922 -556 507978
rect -488 507922 -432 507978
rect -860 490294 -804 490350
rect -736 490294 -680 490350
rect -612 490294 -556 490350
rect -488 490294 -432 490350
rect -860 490170 -804 490226
rect -736 490170 -680 490226
rect -612 490170 -556 490226
rect -488 490170 -432 490226
rect -860 490046 -804 490102
rect -736 490046 -680 490102
rect -612 490046 -556 490102
rect -488 490046 -432 490102
rect -860 489922 -804 489978
rect -736 489922 -680 489978
rect -612 489922 -556 489978
rect -488 489922 -432 489978
rect -860 472294 -804 472350
rect -736 472294 -680 472350
rect -612 472294 -556 472350
rect -488 472294 -432 472350
rect -860 472170 -804 472226
rect -736 472170 -680 472226
rect -612 472170 -556 472226
rect -488 472170 -432 472226
rect -860 472046 -804 472102
rect -736 472046 -680 472102
rect -612 472046 -556 472102
rect -488 472046 -432 472102
rect -860 471922 -804 471978
rect -736 471922 -680 471978
rect -612 471922 -556 471978
rect -488 471922 -432 471978
rect -860 454294 -804 454350
rect -736 454294 -680 454350
rect -612 454294 -556 454350
rect -488 454294 -432 454350
rect -860 454170 -804 454226
rect -736 454170 -680 454226
rect -612 454170 -556 454226
rect -488 454170 -432 454226
rect -860 454046 -804 454102
rect -736 454046 -680 454102
rect -612 454046 -556 454102
rect -488 454046 -432 454102
rect -860 453922 -804 453978
rect -736 453922 -680 453978
rect -612 453922 -556 453978
rect -488 453922 -432 453978
rect -860 436294 -804 436350
rect -736 436294 -680 436350
rect -612 436294 -556 436350
rect -488 436294 -432 436350
rect -860 436170 -804 436226
rect -736 436170 -680 436226
rect -612 436170 -556 436226
rect -488 436170 -432 436226
rect -860 436046 -804 436102
rect -736 436046 -680 436102
rect -612 436046 -556 436102
rect -488 436046 -432 436102
rect -860 435922 -804 435978
rect -736 435922 -680 435978
rect -612 435922 -556 435978
rect -488 435922 -432 435978
rect -860 418294 -804 418350
rect -736 418294 -680 418350
rect -612 418294 -556 418350
rect -488 418294 -432 418350
rect -860 418170 -804 418226
rect -736 418170 -680 418226
rect -612 418170 -556 418226
rect -488 418170 -432 418226
rect -860 418046 -804 418102
rect -736 418046 -680 418102
rect -612 418046 -556 418102
rect -488 418046 -432 418102
rect -860 417922 -804 417978
rect -736 417922 -680 417978
rect -612 417922 -556 417978
rect -488 417922 -432 417978
rect -860 400294 -804 400350
rect -736 400294 -680 400350
rect -612 400294 -556 400350
rect -488 400294 -432 400350
rect -860 400170 -804 400226
rect -736 400170 -680 400226
rect -612 400170 -556 400226
rect -488 400170 -432 400226
rect -860 400046 -804 400102
rect -736 400046 -680 400102
rect -612 400046 -556 400102
rect -488 400046 -432 400102
rect -860 399922 -804 399978
rect -736 399922 -680 399978
rect -612 399922 -556 399978
rect -488 399922 -432 399978
rect -860 382294 -804 382350
rect -736 382294 -680 382350
rect -612 382294 -556 382350
rect -488 382294 -432 382350
rect -860 382170 -804 382226
rect -736 382170 -680 382226
rect -612 382170 -556 382226
rect -488 382170 -432 382226
rect -860 382046 -804 382102
rect -736 382046 -680 382102
rect -612 382046 -556 382102
rect -488 382046 -432 382102
rect -860 381922 -804 381978
rect -736 381922 -680 381978
rect -612 381922 -556 381978
rect -488 381922 -432 381978
rect -860 364294 -804 364350
rect -736 364294 -680 364350
rect -612 364294 -556 364350
rect -488 364294 -432 364350
rect -860 364170 -804 364226
rect -736 364170 -680 364226
rect -612 364170 -556 364226
rect -488 364170 -432 364226
rect -860 364046 -804 364102
rect -736 364046 -680 364102
rect -612 364046 -556 364102
rect -488 364046 -432 364102
rect -860 363922 -804 363978
rect -736 363922 -680 363978
rect -612 363922 -556 363978
rect -488 363922 -432 363978
rect -860 346294 -804 346350
rect -736 346294 -680 346350
rect -612 346294 -556 346350
rect -488 346294 -432 346350
rect -860 346170 -804 346226
rect -736 346170 -680 346226
rect -612 346170 -556 346226
rect -488 346170 -432 346226
rect -860 346046 -804 346102
rect -736 346046 -680 346102
rect -612 346046 -556 346102
rect -488 346046 -432 346102
rect -860 345922 -804 345978
rect -736 345922 -680 345978
rect -612 345922 -556 345978
rect -488 345922 -432 345978
rect -860 328294 -804 328350
rect -736 328294 -680 328350
rect -612 328294 -556 328350
rect -488 328294 -432 328350
rect -860 328170 -804 328226
rect -736 328170 -680 328226
rect -612 328170 -556 328226
rect -488 328170 -432 328226
rect -860 328046 -804 328102
rect -736 328046 -680 328102
rect -612 328046 -556 328102
rect -488 328046 -432 328102
rect -860 327922 -804 327978
rect -736 327922 -680 327978
rect -612 327922 -556 327978
rect -488 327922 -432 327978
rect -860 310294 -804 310350
rect -736 310294 -680 310350
rect -612 310294 -556 310350
rect -488 310294 -432 310350
rect -860 310170 -804 310226
rect -736 310170 -680 310226
rect -612 310170 -556 310226
rect -488 310170 -432 310226
rect -860 310046 -804 310102
rect -736 310046 -680 310102
rect -612 310046 -556 310102
rect -488 310046 -432 310102
rect -860 309922 -804 309978
rect -736 309922 -680 309978
rect -612 309922 -556 309978
rect -488 309922 -432 309978
rect -860 292294 -804 292350
rect -736 292294 -680 292350
rect -612 292294 -556 292350
rect -488 292294 -432 292350
rect -860 292170 -804 292226
rect -736 292170 -680 292226
rect -612 292170 -556 292226
rect -488 292170 -432 292226
rect -860 292046 -804 292102
rect -736 292046 -680 292102
rect -612 292046 -556 292102
rect -488 292046 -432 292102
rect -860 291922 -804 291978
rect -736 291922 -680 291978
rect -612 291922 -556 291978
rect -488 291922 -432 291978
rect -860 274294 -804 274350
rect -736 274294 -680 274350
rect -612 274294 -556 274350
rect -488 274294 -432 274350
rect -860 274170 -804 274226
rect -736 274170 -680 274226
rect -612 274170 -556 274226
rect -488 274170 -432 274226
rect -860 274046 -804 274102
rect -736 274046 -680 274102
rect -612 274046 -556 274102
rect -488 274046 -432 274102
rect -860 273922 -804 273978
rect -736 273922 -680 273978
rect -612 273922 -556 273978
rect -488 273922 -432 273978
rect -860 256294 -804 256350
rect -736 256294 -680 256350
rect -612 256294 -556 256350
rect -488 256294 -432 256350
rect -860 256170 -804 256226
rect -736 256170 -680 256226
rect -612 256170 -556 256226
rect -488 256170 -432 256226
rect -860 256046 -804 256102
rect -736 256046 -680 256102
rect -612 256046 -556 256102
rect -488 256046 -432 256102
rect -860 255922 -804 255978
rect -736 255922 -680 255978
rect -612 255922 -556 255978
rect -488 255922 -432 255978
rect -860 238294 -804 238350
rect -736 238294 -680 238350
rect -612 238294 -556 238350
rect -488 238294 -432 238350
rect -860 238170 -804 238226
rect -736 238170 -680 238226
rect -612 238170 -556 238226
rect -488 238170 -432 238226
rect -860 238046 -804 238102
rect -736 238046 -680 238102
rect -612 238046 -556 238102
rect -488 238046 -432 238102
rect -860 237922 -804 237978
rect -736 237922 -680 237978
rect -612 237922 -556 237978
rect -488 237922 -432 237978
rect -860 220294 -804 220350
rect -736 220294 -680 220350
rect -612 220294 -556 220350
rect -488 220294 -432 220350
rect -860 220170 -804 220226
rect -736 220170 -680 220226
rect -612 220170 -556 220226
rect -488 220170 -432 220226
rect -860 220046 -804 220102
rect -736 220046 -680 220102
rect -612 220046 -556 220102
rect -488 220046 -432 220102
rect -860 219922 -804 219978
rect -736 219922 -680 219978
rect -612 219922 -556 219978
rect -488 219922 -432 219978
rect -860 202294 -804 202350
rect -736 202294 -680 202350
rect -612 202294 -556 202350
rect -488 202294 -432 202350
rect -860 202170 -804 202226
rect -736 202170 -680 202226
rect -612 202170 -556 202226
rect -488 202170 -432 202226
rect -860 202046 -804 202102
rect -736 202046 -680 202102
rect -612 202046 -556 202102
rect -488 202046 -432 202102
rect -860 201922 -804 201978
rect -736 201922 -680 201978
rect -612 201922 -556 201978
rect -488 201922 -432 201978
rect -860 184294 -804 184350
rect -736 184294 -680 184350
rect -612 184294 -556 184350
rect -488 184294 -432 184350
rect -860 184170 -804 184226
rect -736 184170 -680 184226
rect -612 184170 -556 184226
rect -488 184170 -432 184226
rect -860 184046 -804 184102
rect -736 184046 -680 184102
rect -612 184046 -556 184102
rect -488 184046 -432 184102
rect -860 183922 -804 183978
rect -736 183922 -680 183978
rect -612 183922 -556 183978
rect -488 183922 -432 183978
rect -860 166294 -804 166350
rect -736 166294 -680 166350
rect -612 166294 -556 166350
rect -488 166294 -432 166350
rect -860 166170 -804 166226
rect -736 166170 -680 166226
rect -612 166170 -556 166226
rect -488 166170 -432 166226
rect -860 166046 -804 166102
rect -736 166046 -680 166102
rect -612 166046 -556 166102
rect -488 166046 -432 166102
rect -860 165922 -804 165978
rect -736 165922 -680 165978
rect -612 165922 -556 165978
rect -488 165922 -432 165978
rect -860 148294 -804 148350
rect -736 148294 -680 148350
rect -612 148294 -556 148350
rect -488 148294 -432 148350
rect -860 148170 -804 148226
rect -736 148170 -680 148226
rect -612 148170 -556 148226
rect -488 148170 -432 148226
rect -860 148046 -804 148102
rect -736 148046 -680 148102
rect -612 148046 -556 148102
rect -488 148046 -432 148102
rect -860 147922 -804 147978
rect -736 147922 -680 147978
rect -612 147922 -556 147978
rect -488 147922 -432 147978
rect -860 130294 -804 130350
rect -736 130294 -680 130350
rect -612 130294 -556 130350
rect -488 130294 -432 130350
rect -860 130170 -804 130226
rect -736 130170 -680 130226
rect -612 130170 -556 130226
rect -488 130170 -432 130226
rect -860 130046 -804 130102
rect -736 130046 -680 130102
rect -612 130046 -556 130102
rect -488 130046 -432 130102
rect -860 129922 -804 129978
rect -736 129922 -680 129978
rect -612 129922 -556 129978
rect -488 129922 -432 129978
rect -860 112294 -804 112350
rect -736 112294 -680 112350
rect -612 112294 -556 112350
rect -488 112294 -432 112350
rect -860 112170 -804 112226
rect -736 112170 -680 112226
rect -612 112170 -556 112226
rect -488 112170 -432 112226
rect -860 112046 -804 112102
rect -736 112046 -680 112102
rect -612 112046 -556 112102
rect -488 112046 -432 112102
rect -860 111922 -804 111978
rect -736 111922 -680 111978
rect -612 111922 -556 111978
rect -488 111922 -432 111978
rect -860 94294 -804 94350
rect -736 94294 -680 94350
rect -612 94294 -556 94350
rect -488 94294 -432 94350
rect -860 94170 -804 94226
rect -736 94170 -680 94226
rect -612 94170 -556 94226
rect -488 94170 -432 94226
rect -860 94046 -804 94102
rect -736 94046 -680 94102
rect -612 94046 -556 94102
rect -488 94046 -432 94102
rect -860 93922 -804 93978
rect -736 93922 -680 93978
rect -612 93922 -556 93978
rect -488 93922 -432 93978
rect -860 76294 -804 76350
rect -736 76294 -680 76350
rect -612 76294 -556 76350
rect -488 76294 -432 76350
rect -860 76170 -804 76226
rect -736 76170 -680 76226
rect -612 76170 -556 76226
rect -488 76170 -432 76226
rect -860 76046 -804 76102
rect -736 76046 -680 76102
rect -612 76046 -556 76102
rect -488 76046 -432 76102
rect -860 75922 -804 75978
rect -736 75922 -680 75978
rect -612 75922 -556 75978
rect -488 75922 -432 75978
rect -860 58294 -804 58350
rect -736 58294 -680 58350
rect -612 58294 -556 58350
rect -488 58294 -432 58350
rect -860 58170 -804 58226
rect -736 58170 -680 58226
rect -612 58170 -556 58226
rect -488 58170 -432 58226
rect -860 58046 -804 58102
rect -736 58046 -680 58102
rect -612 58046 -556 58102
rect -488 58046 -432 58102
rect -860 57922 -804 57978
rect -736 57922 -680 57978
rect -612 57922 -556 57978
rect -488 57922 -432 57978
rect -860 40294 -804 40350
rect -736 40294 -680 40350
rect -612 40294 -556 40350
rect -488 40294 -432 40350
rect -860 40170 -804 40226
rect -736 40170 -680 40226
rect -612 40170 -556 40226
rect -488 40170 -432 40226
rect -860 40046 -804 40102
rect -736 40046 -680 40102
rect -612 40046 -556 40102
rect -488 40046 -432 40102
rect -860 39922 -804 39978
rect -736 39922 -680 39978
rect -612 39922 -556 39978
rect -488 39922 -432 39978
rect -860 22294 -804 22350
rect -736 22294 -680 22350
rect -612 22294 -556 22350
rect -488 22294 -432 22350
rect -860 22170 -804 22226
rect -736 22170 -680 22226
rect -612 22170 -556 22226
rect -488 22170 -432 22226
rect -860 22046 -804 22102
rect -736 22046 -680 22102
rect -612 22046 -556 22102
rect -488 22046 -432 22102
rect -860 21922 -804 21978
rect -736 21922 -680 21978
rect -612 21922 -556 21978
rect -488 21922 -432 21978
rect -860 4294 -804 4350
rect -736 4294 -680 4350
rect -612 4294 -556 4350
rect -488 4294 -432 4350
rect -860 4170 -804 4226
rect -736 4170 -680 4226
rect -612 4170 -556 4226
rect -488 4170 -432 4226
rect -860 4046 -804 4102
rect -736 4046 -680 4102
rect -612 4046 -556 4102
rect -488 4046 -432 4102
rect -860 3922 -804 3978
rect -736 3922 -680 3978
rect -612 3922 -556 3978
rect -488 3922 -432 3978
rect -860 -216 -804 -160
rect -736 -216 -680 -160
rect -612 -216 -556 -160
rect -488 -216 -432 -160
rect -860 -340 -804 -284
rect -736 -340 -680 -284
rect -612 -340 -556 -284
rect -488 -340 -432 -284
rect -860 -464 -804 -408
rect -736 -464 -680 -408
rect -612 -464 -556 -408
rect -488 -464 -432 -408
rect -860 -588 -804 -532
rect -736 -588 -680 -532
rect -612 -588 -556 -532
rect -488 -588 -432 -532
rect 3250 597156 3306 597212
rect 3374 597156 3430 597212
rect 3498 597156 3554 597212
rect 3622 597156 3678 597212
rect 3250 597032 3306 597088
rect 3374 597032 3430 597088
rect 3498 597032 3554 597088
rect 3622 597032 3678 597088
rect 3250 596908 3306 596964
rect 3374 596908 3430 596964
rect 3498 596908 3554 596964
rect 3622 596908 3678 596964
rect 3250 596784 3306 596840
rect 3374 596784 3430 596840
rect 3498 596784 3554 596840
rect 3622 596784 3678 596840
rect 3250 580294 3306 580350
rect 3374 580294 3430 580350
rect 3498 580294 3554 580350
rect 3622 580294 3678 580350
rect 3250 580170 3306 580226
rect 3374 580170 3430 580226
rect 3498 580170 3554 580226
rect 3622 580170 3678 580226
rect 3250 580046 3306 580102
rect 3374 580046 3430 580102
rect 3498 580046 3554 580102
rect 3622 580046 3678 580102
rect 3250 579922 3306 579978
rect 3374 579922 3430 579978
rect 3498 579922 3554 579978
rect 3622 579922 3678 579978
rect 3250 562294 3306 562350
rect 3374 562294 3430 562350
rect 3498 562294 3554 562350
rect 3622 562294 3678 562350
rect 3250 562170 3306 562226
rect 3374 562170 3430 562226
rect 3498 562170 3554 562226
rect 3622 562170 3678 562226
rect 3250 562046 3306 562102
rect 3374 562046 3430 562102
rect 3498 562046 3554 562102
rect 3622 562046 3678 562102
rect 3250 561922 3306 561978
rect 3374 561922 3430 561978
rect 3498 561922 3554 561978
rect 3622 561922 3678 561978
rect 3250 544294 3306 544350
rect 3374 544294 3430 544350
rect 3498 544294 3554 544350
rect 3622 544294 3678 544350
rect 3250 544170 3306 544226
rect 3374 544170 3430 544226
rect 3498 544170 3554 544226
rect 3622 544170 3678 544226
rect 3250 544046 3306 544102
rect 3374 544046 3430 544102
rect 3498 544046 3554 544102
rect 3622 544046 3678 544102
rect 3250 543922 3306 543978
rect 3374 543922 3430 543978
rect 3498 543922 3554 543978
rect 3622 543922 3678 543978
rect 3250 526294 3306 526350
rect 3374 526294 3430 526350
rect 3498 526294 3554 526350
rect 3622 526294 3678 526350
rect 3250 526170 3306 526226
rect 3374 526170 3430 526226
rect 3498 526170 3554 526226
rect 3622 526170 3678 526226
rect 3250 526046 3306 526102
rect 3374 526046 3430 526102
rect 3498 526046 3554 526102
rect 3622 526046 3678 526102
rect 3250 525922 3306 525978
rect 3374 525922 3430 525978
rect 3498 525922 3554 525978
rect 3622 525922 3678 525978
rect 3250 508294 3306 508350
rect 3374 508294 3430 508350
rect 3498 508294 3554 508350
rect 3622 508294 3678 508350
rect 3250 508170 3306 508226
rect 3374 508170 3430 508226
rect 3498 508170 3554 508226
rect 3622 508170 3678 508226
rect 3250 508046 3306 508102
rect 3374 508046 3430 508102
rect 3498 508046 3554 508102
rect 3622 508046 3678 508102
rect 3250 507922 3306 507978
rect 3374 507922 3430 507978
rect 3498 507922 3554 507978
rect 3622 507922 3678 507978
rect 3250 490294 3306 490350
rect 3374 490294 3430 490350
rect 3498 490294 3554 490350
rect 3622 490294 3678 490350
rect 3250 490170 3306 490226
rect 3374 490170 3430 490226
rect 3498 490170 3554 490226
rect 3622 490170 3678 490226
rect 3250 490046 3306 490102
rect 3374 490046 3430 490102
rect 3498 490046 3554 490102
rect 3622 490046 3678 490102
rect 3250 489922 3306 489978
rect 3374 489922 3430 489978
rect 3498 489922 3554 489978
rect 3622 489922 3678 489978
rect 3250 472294 3306 472350
rect 3374 472294 3430 472350
rect 3498 472294 3554 472350
rect 3622 472294 3678 472350
rect 3250 472170 3306 472226
rect 3374 472170 3430 472226
rect 3498 472170 3554 472226
rect 3622 472170 3678 472226
rect 3250 472046 3306 472102
rect 3374 472046 3430 472102
rect 3498 472046 3554 472102
rect 3622 472046 3678 472102
rect 3250 471922 3306 471978
rect 3374 471922 3430 471978
rect 3498 471922 3554 471978
rect 3622 471922 3678 471978
rect 3250 454294 3306 454350
rect 3374 454294 3430 454350
rect 3498 454294 3554 454350
rect 3622 454294 3678 454350
rect 3250 454170 3306 454226
rect 3374 454170 3430 454226
rect 3498 454170 3554 454226
rect 3622 454170 3678 454226
rect 3250 454046 3306 454102
rect 3374 454046 3430 454102
rect 3498 454046 3554 454102
rect 3622 454046 3678 454102
rect 3250 453922 3306 453978
rect 3374 453922 3430 453978
rect 3498 453922 3554 453978
rect 3622 453922 3678 453978
rect 3250 436294 3306 436350
rect 3374 436294 3430 436350
rect 3498 436294 3554 436350
rect 3622 436294 3678 436350
rect 3250 436170 3306 436226
rect 3374 436170 3430 436226
rect 3498 436170 3554 436226
rect 3622 436170 3678 436226
rect 3250 436046 3306 436102
rect 3374 436046 3430 436102
rect 3498 436046 3554 436102
rect 3622 436046 3678 436102
rect 3250 435922 3306 435978
rect 3374 435922 3430 435978
rect 3498 435922 3554 435978
rect 3622 435922 3678 435978
rect 3250 418294 3306 418350
rect 3374 418294 3430 418350
rect 3498 418294 3554 418350
rect 3622 418294 3678 418350
rect 3250 418170 3306 418226
rect 3374 418170 3430 418226
rect 3498 418170 3554 418226
rect 3622 418170 3678 418226
rect 3250 418046 3306 418102
rect 3374 418046 3430 418102
rect 3498 418046 3554 418102
rect 3622 418046 3678 418102
rect 3250 417922 3306 417978
rect 3374 417922 3430 417978
rect 3498 417922 3554 417978
rect 3622 417922 3678 417978
rect 3250 400294 3306 400350
rect 3374 400294 3430 400350
rect 3498 400294 3554 400350
rect 3622 400294 3678 400350
rect 3250 400170 3306 400226
rect 3374 400170 3430 400226
rect 3498 400170 3554 400226
rect 3622 400170 3678 400226
rect 3250 400046 3306 400102
rect 3374 400046 3430 400102
rect 3498 400046 3554 400102
rect 3622 400046 3678 400102
rect 3250 399922 3306 399978
rect 3374 399922 3430 399978
rect 3498 399922 3554 399978
rect 3622 399922 3678 399978
rect 3250 382294 3306 382350
rect 3374 382294 3430 382350
rect 3498 382294 3554 382350
rect 3622 382294 3678 382350
rect 3250 382170 3306 382226
rect 3374 382170 3430 382226
rect 3498 382170 3554 382226
rect 3622 382170 3678 382226
rect 3250 382046 3306 382102
rect 3374 382046 3430 382102
rect 3498 382046 3554 382102
rect 3622 382046 3678 382102
rect 3250 381922 3306 381978
rect 3374 381922 3430 381978
rect 3498 381922 3554 381978
rect 3622 381922 3678 381978
rect 3250 364294 3306 364350
rect 3374 364294 3430 364350
rect 3498 364294 3554 364350
rect 3622 364294 3678 364350
rect 3250 364170 3306 364226
rect 3374 364170 3430 364226
rect 3498 364170 3554 364226
rect 3622 364170 3678 364226
rect 3250 364046 3306 364102
rect 3374 364046 3430 364102
rect 3498 364046 3554 364102
rect 3622 364046 3678 364102
rect 3250 363922 3306 363978
rect 3374 363922 3430 363978
rect 3498 363922 3554 363978
rect 3622 363922 3678 363978
rect 3250 346294 3306 346350
rect 3374 346294 3430 346350
rect 3498 346294 3554 346350
rect 3622 346294 3678 346350
rect 3250 346170 3306 346226
rect 3374 346170 3430 346226
rect 3498 346170 3554 346226
rect 3622 346170 3678 346226
rect 3250 346046 3306 346102
rect 3374 346046 3430 346102
rect 3498 346046 3554 346102
rect 3622 346046 3678 346102
rect 3250 345922 3306 345978
rect 3374 345922 3430 345978
rect 3498 345922 3554 345978
rect 3622 345922 3678 345978
rect 3250 328294 3306 328350
rect 3374 328294 3430 328350
rect 3498 328294 3554 328350
rect 3622 328294 3678 328350
rect 3250 328170 3306 328226
rect 3374 328170 3430 328226
rect 3498 328170 3554 328226
rect 3622 328170 3678 328226
rect 3250 328046 3306 328102
rect 3374 328046 3430 328102
rect 3498 328046 3554 328102
rect 3622 328046 3678 328102
rect 3250 327922 3306 327978
rect 3374 327922 3430 327978
rect 3498 327922 3554 327978
rect 3622 327922 3678 327978
rect 3250 310294 3306 310350
rect 3374 310294 3430 310350
rect 3498 310294 3554 310350
rect 3622 310294 3678 310350
rect 3250 310170 3306 310226
rect 3374 310170 3430 310226
rect 3498 310170 3554 310226
rect 3622 310170 3678 310226
rect 3250 310046 3306 310102
rect 3374 310046 3430 310102
rect 3498 310046 3554 310102
rect 3622 310046 3678 310102
rect 3250 309922 3306 309978
rect 3374 309922 3430 309978
rect 3498 309922 3554 309978
rect 3622 309922 3678 309978
rect 3250 292294 3306 292350
rect 3374 292294 3430 292350
rect 3498 292294 3554 292350
rect 3622 292294 3678 292350
rect 3250 292170 3306 292226
rect 3374 292170 3430 292226
rect 3498 292170 3554 292226
rect 3622 292170 3678 292226
rect 3250 292046 3306 292102
rect 3374 292046 3430 292102
rect 3498 292046 3554 292102
rect 3622 292046 3678 292102
rect 3250 291922 3306 291978
rect 3374 291922 3430 291978
rect 3498 291922 3554 291978
rect 3622 291922 3678 291978
rect 3250 274294 3306 274350
rect 3374 274294 3430 274350
rect 3498 274294 3554 274350
rect 3622 274294 3678 274350
rect 3250 274170 3306 274226
rect 3374 274170 3430 274226
rect 3498 274170 3554 274226
rect 3622 274170 3678 274226
rect 3250 274046 3306 274102
rect 3374 274046 3430 274102
rect 3498 274046 3554 274102
rect 3622 274046 3678 274102
rect 3250 273922 3306 273978
rect 3374 273922 3430 273978
rect 3498 273922 3554 273978
rect 3622 273922 3678 273978
rect 3250 256294 3306 256350
rect 3374 256294 3430 256350
rect 3498 256294 3554 256350
rect 3622 256294 3678 256350
rect 3250 256170 3306 256226
rect 3374 256170 3430 256226
rect 3498 256170 3554 256226
rect 3622 256170 3678 256226
rect 3250 256046 3306 256102
rect 3374 256046 3430 256102
rect 3498 256046 3554 256102
rect 3622 256046 3678 256102
rect 3250 255922 3306 255978
rect 3374 255922 3430 255978
rect 3498 255922 3554 255978
rect 3622 255922 3678 255978
rect 3250 238294 3306 238350
rect 3374 238294 3430 238350
rect 3498 238294 3554 238350
rect 3622 238294 3678 238350
rect 3250 238170 3306 238226
rect 3374 238170 3430 238226
rect 3498 238170 3554 238226
rect 3622 238170 3678 238226
rect 3250 238046 3306 238102
rect 3374 238046 3430 238102
rect 3498 238046 3554 238102
rect 3622 238046 3678 238102
rect 3250 237922 3306 237978
rect 3374 237922 3430 237978
rect 3498 237922 3554 237978
rect 3622 237922 3678 237978
rect 3250 220294 3306 220350
rect 3374 220294 3430 220350
rect 3498 220294 3554 220350
rect 3622 220294 3678 220350
rect 3250 220170 3306 220226
rect 3374 220170 3430 220226
rect 3498 220170 3554 220226
rect 3622 220170 3678 220226
rect 3250 220046 3306 220102
rect 3374 220046 3430 220102
rect 3498 220046 3554 220102
rect 3622 220046 3678 220102
rect 3250 219922 3306 219978
rect 3374 219922 3430 219978
rect 3498 219922 3554 219978
rect 3622 219922 3678 219978
rect 3250 202294 3306 202350
rect 3374 202294 3430 202350
rect 3498 202294 3554 202350
rect 3622 202294 3678 202350
rect 3250 202170 3306 202226
rect 3374 202170 3430 202226
rect 3498 202170 3554 202226
rect 3622 202170 3678 202226
rect 3250 202046 3306 202102
rect 3374 202046 3430 202102
rect 3498 202046 3554 202102
rect 3622 202046 3678 202102
rect 3250 201922 3306 201978
rect 3374 201922 3430 201978
rect 3498 201922 3554 201978
rect 3622 201922 3678 201978
rect 3250 184294 3306 184350
rect 3374 184294 3430 184350
rect 3498 184294 3554 184350
rect 3622 184294 3678 184350
rect 3250 184170 3306 184226
rect 3374 184170 3430 184226
rect 3498 184170 3554 184226
rect 3622 184170 3678 184226
rect 3250 184046 3306 184102
rect 3374 184046 3430 184102
rect 3498 184046 3554 184102
rect 3622 184046 3678 184102
rect 3250 183922 3306 183978
rect 3374 183922 3430 183978
rect 3498 183922 3554 183978
rect 3622 183922 3678 183978
rect 3250 166294 3306 166350
rect 3374 166294 3430 166350
rect 3498 166294 3554 166350
rect 3622 166294 3678 166350
rect 3250 166170 3306 166226
rect 3374 166170 3430 166226
rect 3498 166170 3554 166226
rect 3622 166170 3678 166226
rect 3250 166046 3306 166102
rect 3374 166046 3430 166102
rect 3498 166046 3554 166102
rect 3622 166046 3678 166102
rect 3250 165922 3306 165978
rect 3374 165922 3430 165978
rect 3498 165922 3554 165978
rect 3622 165922 3678 165978
rect 3250 148294 3306 148350
rect 3374 148294 3430 148350
rect 3498 148294 3554 148350
rect 3622 148294 3678 148350
rect 3250 148170 3306 148226
rect 3374 148170 3430 148226
rect 3498 148170 3554 148226
rect 3622 148170 3678 148226
rect 3250 148046 3306 148102
rect 3374 148046 3430 148102
rect 3498 148046 3554 148102
rect 3622 148046 3678 148102
rect 3250 147922 3306 147978
rect 3374 147922 3430 147978
rect 3498 147922 3554 147978
rect 3622 147922 3678 147978
rect 3250 130294 3306 130350
rect 3374 130294 3430 130350
rect 3498 130294 3554 130350
rect 3622 130294 3678 130350
rect 3250 130170 3306 130226
rect 3374 130170 3430 130226
rect 3498 130170 3554 130226
rect 3622 130170 3678 130226
rect 3250 130046 3306 130102
rect 3374 130046 3430 130102
rect 3498 130046 3554 130102
rect 3622 130046 3678 130102
rect 3250 129922 3306 129978
rect 3374 129922 3430 129978
rect 3498 129922 3554 129978
rect 3622 129922 3678 129978
rect 3250 112294 3306 112350
rect 3374 112294 3430 112350
rect 3498 112294 3554 112350
rect 3622 112294 3678 112350
rect 3250 112170 3306 112226
rect 3374 112170 3430 112226
rect 3498 112170 3554 112226
rect 3622 112170 3678 112226
rect 3250 112046 3306 112102
rect 3374 112046 3430 112102
rect 3498 112046 3554 112102
rect 3622 112046 3678 112102
rect 3250 111922 3306 111978
rect 3374 111922 3430 111978
rect 3498 111922 3554 111978
rect 3622 111922 3678 111978
rect 3250 94294 3306 94350
rect 3374 94294 3430 94350
rect 3498 94294 3554 94350
rect 3622 94294 3678 94350
rect 3250 94170 3306 94226
rect 3374 94170 3430 94226
rect 3498 94170 3554 94226
rect 3622 94170 3678 94226
rect 3250 94046 3306 94102
rect 3374 94046 3430 94102
rect 3498 94046 3554 94102
rect 3622 94046 3678 94102
rect 3250 93922 3306 93978
rect 3374 93922 3430 93978
rect 3498 93922 3554 93978
rect 3622 93922 3678 93978
rect 3250 76294 3306 76350
rect 3374 76294 3430 76350
rect 3498 76294 3554 76350
rect 3622 76294 3678 76350
rect 3250 76170 3306 76226
rect 3374 76170 3430 76226
rect 3498 76170 3554 76226
rect 3622 76170 3678 76226
rect 3250 76046 3306 76102
rect 3374 76046 3430 76102
rect 3498 76046 3554 76102
rect 3622 76046 3678 76102
rect 3250 75922 3306 75978
rect 3374 75922 3430 75978
rect 3498 75922 3554 75978
rect 3622 75922 3678 75978
rect 3250 58294 3306 58350
rect 3374 58294 3430 58350
rect 3498 58294 3554 58350
rect 3622 58294 3678 58350
rect 3250 58170 3306 58226
rect 3374 58170 3430 58226
rect 3498 58170 3554 58226
rect 3622 58170 3678 58226
rect 3250 58046 3306 58102
rect 3374 58046 3430 58102
rect 3498 58046 3554 58102
rect 3622 58046 3678 58102
rect 3250 57922 3306 57978
rect 3374 57922 3430 57978
rect 3498 57922 3554 57978
rect 3622 57922 3678 57978
rect 3250 40294 3306 40350
rect 3374 40294 3430 40350
rect 3498 40294 3554 40350
rect 3622 40294 3678 40350
rect 3250 40170 3306 40226
rect 3374 40170 3430 40226
rect 3498 40170 3554 40226
rect 3622 40170 3678 40226
rect 3250 40046 3306 40102
rect 3374 40046 3430 40102
rect 3498 40046 3554 40102
rect 3622 40046 3678 40102
rect 3250 39922 3306 39978
rect 3374 39922 3430 39978
rect 3498 39922 3554 39978
rect 3622 39922 3678 39978
rect 3250 22294 3306 22350
rect 3374 22294 3430 22350
rect 3498 22294 3554 22350
rect 3622 22294 3678 22350
rect 3250 22170 3306 22226
rect 3374 22170 3430 22226
rect 3498 22170 3554 22226
rect 3622 22170 3678 22226
rect 3250 22046 3306 22102
rect 3374 22046 3430 22102
rect 3498 22046 3554 22102
rect 3622 22046 3678 22102
rect 3250 21922 3306 21978
rect 3374 21922 3430 21978
rect 3498 21922 3554 21978
rect 3622 21922 3678 21978
rect 3250 4294 3306 4350
rect 3374 4294 3430 4350
rect 3498 4294 3554 4350
rect 3622 4294 3678 4350
rect 3250 4170 3306 4226
rect 3374 4170 3430 4226
rect 3498 4170 3554 4226
rect 3622 4170 3678 4226
rect 3250 4046 3306 4102
rect 3374 4046 3430 4102
rect 3498 4046 3554 4102
rect 3622 4046 3678 4102
rect 3250 3922 3306 3978
rect 3374 3922 3430 3978
rect 3498 3922 3554 3978
rect 3622 3922 3678 3978
rect 3250 -216 3306 -160
rect 3374 -216 3430 -160
rect 3498 -216 3554 -160
rect 3622 -216 3678 -160
rect 3250 -340 3306 -284
rect 3374 -340 3430 -284
rect 3498 -340 3554 -284
rect 3622 -340 3678 -284
rect 3250 -464 3306 -408
rect 3374 -464 3430 -408
rect 3498 -464 3554 -408
rect 3622 -464 3678 -408
rect 3250 -588 3306 -532
rect 3374 -588 3430 -532
rect 3498 -588 3554 -532
rect 3622 -588 3678 -532
rect -1820 -1176 -1764 -1120
rect -1696 -1176 -1640 -1120
rect -1572 -1176 -1516 -1120
rect -1448 -1176 -1392 -1120
rect -1820 -1300 -1764 -1244
rect -1696 -1300 -1640 -1244
rect -1572 -1300 -1516 -1244
rect -1448 -1300 -1392 -1244
rect -1820 -1424 -1764 -1368
rect -1696 -1424 -1640 -1368
rect -1572 -1424 -1516 -1368
rect -1448 -1424 -1392 -1368
rect -1820 -1548 -1764 -1492
rect -1696 -1548 -1640 -1492
rect -1572 -1548 -1516 -1492
rect -1448 -1548 -1392 -1492
rect 6970 598116 7026 598172
rect 7094 598116 7150 598172
rect 7218 598116 7274 598172
rect 7342 598116 7398 598172
rect 6970 597992 7026 598048
rect 7094 597992 7150 598048
rect 7218 597992 7274 598048
rect 7342 597992 7398 598048
rect 6970 597868 7026 597924
rect 7094 597868 7150 597924
rect 7218 597868 7274 597924
rect 7342 597868 7398 597924
rect 6970 597744 7026 597800
rect 7094 597744 7150 597800
rect 7218 597744 7274 597800
rect 7342 597744 7398 597800
rect 21250 597156 21306 597212
rect 21374 597156 21430 597212
rect 21498 597156 21554 597212
rect 21622 597156 21678 597212
rect 21250 597032 21306 597088
rect 21374 597032 21430 597088
rect 21498 597032 21554 597088
rect 21622 597032 21678 597088
rect 21250 596908 21306 596964
rect 21374 596908 21430 596964
rect 21498 596908 21554 596964
rect 21622 596908 21678 596964
rect 21250 596784 21306 596840
rect 21374 596784 21430 596840
rect 21498 596784 21554 596840
rect 21622 596784 21678 596840
rect 6970 586294 7026 586350
rect 7094 586294 7150 586350
rect 7218 586294 7274 586350
rect 7342 586294 7398 586350
rect 6970 586170 7026 586226
rect 7094 586170 7150 586226
rect 7218 586170 7274 586226
rect 7342 586170 7398 586226
rect 6970 586046 7026 586102
rect 7094 586046 7150 586102
rect 7218 586046 7274 586102
rect 7342 586046 7398 586102
rect 6970 585922 7026 585978
rect 7094 585922 7150 585978
rect 7218 585922 7274 585978
rect 7342 585922 7398 585978
rect 6970 568294 7026 568350
rect 7094 568294 7150 568350
rect 7218 568294 7274 568350
rect 7342 568294 7398 568350
rect 6970 568170 7026 568226
rect 7094 568170 7150 568226
rect 7218 568170 7274 568226
rect 7342 568170 7398 568226
rect 6970 568046 7026 568102
rect 7094 568046 7150 568102
rect 7218 568046 7274 568102
rect 7342 568046 7398 568102
rect 6970 567922 7026 567978
rect 7094 567922 7150 567978
rect 7218 567922 7274 567978
rect 7342 567922 7398 567978
rect 6970 550294 7026 550350
rect 7094 550294 7150 550350
rect 7218 550294 7274 550350
rect 7342 550294 7398 550350
rect 6970 550170 7026 550226
rect 7094 550170 7150 550226
rect 7218 550170 7274 550226
rect 7342 550170 7398 550226
rect 6970 550046 7026 550102
rect 7094 550046 7150 550102
rect 7218 550046 7274 550102
rect 7342 550046 7398 550102
rect 6970 549922 7026 549978
rect 7094 549922 7150 549978
rect 7218 549922 7274 549978
rect 7342 549922 7398 549978
rect 6970 532294 7026 532350
rect 7094 532294 7150 532350
rect 7218 532294 7274 532350
rect 7342 532294 7398 532350
rect 6970 532170 7026 532226
rect 7094 532170 7150 532226
rect 7218 532170 7274 532226
rect 7342 532170 7398 532226
rect 6970 532046 7026 532102
rect 7094 532046 7150 532102
rect 7218 532046 7274 532102
rect 7342 532046 7398 532102
rect 6970 531922 7026 531978
rect 7094 531922 7150 531978
rect 7218 531922 7274 531978
rect 7342 531922 7398 531978
rect 6970 514294 7026 514350
rect 7094 514294 7150 514350
rect 7218 514294 7274 514350
rect 7342 514294 7398 514350
rect 6970 514170 7026 514226
rect 7094 514170 7150 514226
rect 7218 514170 7274 514226
rect 7342 514170 7398 514226
rect 6970 514046 7026 514102
rect 7094 514046 7150 514102
rect 7218 514046 7274 514102
rect 7342 514046 7398 514102
rect 6970 513922 7026 513978
rect 7094 513922 7150 513978
rect 7218 513922 7274 513978
rect 7342 513922 7398 513978
rect 6970 496294 7026 496350
rect 7094 496294 7150 496350
rect 7218 496294 7274 496350
rect 7342 496294 7398 496350
rect 6970 496170 7026 496226
rect 7094 496170 7150 496226
rect 7218 496170 7274 496226
rect 7342 496170 7398 496226
rect 6970 496046 7026 496102
rect 7094 496046 7150 496102
rect 7218 496046 7274 496102
rect 7342 496046 7398 496102
rect 6970 495922 7026 495978
rect 7094 495922 7150 495978
rect 7218 495922 7274 495978
rect 7342 495922 7398 495978
rect 6970 478294 7026 478350
rect 7094 478294 7150 478350
rect 7218 478294 7274 478350
rect 7342 478294 7398 478350
rect 6970 478170 7026 478226
rect 7094 478170 7150 478226
rect 7218 478170 7274 478226
rect 7342 478170 7398 478226
rect 6970 478046 7026 478102
rect 7094 478046 7150 478102
rect 7218 478046 7274 478102
rect 7342 478046 7398 478102
rect 6970 477922 7026 477978
rect 7094 477922 7150 477978
rect 7218 477922 7274 477978
rect 7342 477922 7398 477978
rect 6970 460294 7026 460350
rect 7094 460294 7150 460350
rect 7218 460294 7274 460350
rect 7342 460294 7398 460350
rect 6970 460170 7026 460226
rect 7094 460170 7150 460226
rect 7218 460170 7274 460226
rect 7342 460170 7398 460226
rect 6970 460046 7026 460102
rect 7094 460046 7150 460102
rect 7218 460046 7274 460102
rect 7342 460046 7398 460102
rect 6970 459922 7026 459978
rect 7094 459922 7150 459978
rect 7218 459922 7274 459978
rect 7342 459922 7398 459978
rect 6970 442294 7026 442350
rect 7094 442294 7150 442350
rect 7218 442294 7274 442350
rect 7342 442294 7398 442350
rect 6970 442170 7026 442226
rect 7094 442170 7150 442226
rect 7218 442170 7274 442226
rect 7342 442170 7398 442226
rect 6970 442046 7026 442102
rect 7094 442046 7150 442102
rect 7218 442046 7274 442102
rect 7342 442046 7398 442102
rect 6970 441922 7026 441978
rect 7094 441922 7150 441978
rect 7218 441922 7274 441978
rect 7342 441922 7398 441978
rect 6970 424294 7026 424350
rect 7094 424294 7150 424350
rect 7218 424294 7274 424350
rect 7342 424294 7398 424350
rect 6970 424170 7026 424226
rect 7094 424170 7150 424226
rect 7218 424170 7274 424226
rect 7342 424170 7398 424226
rect 6970 424046 7026 424102
rect 7094 424046 7150 424102
rect 7218 424046 7274 424102
rect 7342 424046 7398 424102
rect 6970 423922 7026 423978
rect 7094 423922 7150 423978
rect 7218 423922 7274 423978
rect 7342 423922 7398 423978
rect 6970 406294 7026 406350
rect 7094 406294 7150 406350
rect 7218 406294 7274 406350
rect 7342 406294 7398 406350
rect 6970 406170 7026 406226
rect 7094 406170 7150 406226
rect 7218 406170 7274 406226
rect 7342 406170 7398 406226
rect 6970 406046 7026 406102
rect 7094 406046 7150 406102
rect 7218 406046 7274 406102
rect 7342 406046 7398 406102
rect 6970 405922 7026 405978
rect 7094 405922 7150 405978
rect 7218 405922 7274 405978
rect 7342 405922 7398 405978
rect 6970 388294 7026 388350
rect 7094 388294 7150 388350
rect 7218 388294 7274 388350
rect 7342 388294 7398 388350
rect 6970 388170 7026 388226
rect 7094 388170 7150 388226
rect 7218 388170 7274 388226
rect 7342 388170 7398 388226
rect 6970 388046 7026 388102
rect 7094 388046 7150 388102
rect 7218 388046 7274 388102
rect 7342 388046 7398 388102
rect 6970 387922 7026 387978
rect 7094 387922 7150 387978
rect 7218 387922 7274 387978
rect 7342 387922 7398 387978
rect 6970 370294 7026 370350
rect 7094 370294 7150 370350
rect 7218 370294 7274 370350
rect 7342 370294 7398 370350
rect 6970 370170 7026 370226
rect 7094 370170 7150 370226
rect 7218 370170 7274 370226
rect 7342 370170 7398 370226
rect 6970 370046 7026 370102
rect 7094 370046 7150 370102
rect 7218 370046 7274 370102
rect 7342 370046 7398 370102
rect 6970 369922 7026 369978
rect 7094 369922 7150 369978
rect 7218 369922 7274 369978
rect 7342 369922 7398 369978
rect 6970 352294 7026 352350
rect 7094 352294 7150 352350
rect 7218 352294 7274 352350
rect 7342 352294 7398 352350
rect 6970 352170 7026 352226
rect 7094 352170 7150 352226
rect 7218 352170 7274 352226
rect 7342 352170 7398 352226
rect 6970 352046 7026 352102
rect 7094 352046 7150 352102
rect 7218 352046 7274 352102
rect 7342 352046 7398 352102
rect 6970 351922 7026 351978
rect 7094 351922 7150 351978
rect 7218 351922 7274 351978
rect 7342 351922 7398 351978
rect 6970 334294 7026 334350
rect 7094 334294 7150 334350
rect 7218 334294 7274 334350
rect 7342 334294 7398 334350
rect 6970 334170 7026 334226
rect 7094 334170 7150 334226
rect 7218 334170 7274 334226
rect 7342 334170 7398 334226
rect 6970 334046 7026 334102
rect 7094 334046 7150 334102
rect 7218 334046 7274 334102
rect 7342 334046 7398 334102
rect 6970 333922 7026 333978
rect 7094 333922 7150 333978
rect 7218 333922 7274 333978
rect 7342 333922 7398 333978
rect 6970 316294 7026 316350
rect 7094 316294 7150 316350
rect 7218 316294 7274 316350
rect 7342 316294 7398 316350
rect 6970 316170 7026 316226
rect 7094 316170 7150 316226
rect 7218 316170 7274 316226
rect 7342 316170 7398 316226
rect 6970 316046 7026 316102
rect 7094 316046 7150 316102
rect 7218 316046 7274 316102
rect 7342 316046 7398 316102
rect 6970 315922 7026 315978
rect 7094 315922 7150 315978
rect 7218 315922 7274 315978
rect 7342 315922 7398 315978
rect 6970 298294 7026 298350
rect 7094 298294 7150 298350
rect 7218 298294 7274 298350
rect 7342 298294 7398 298350
rect 6970 298170 7026 298226
rect 7094 298170 7150 298226
rect 7218 298170 7274 298226
rect 7342 298170 7398 298226
rect 6970 298046 7026 298102
rect 7094 298046 7150 298102
rect 7218 298046 7274 298102
rect 7342 298046 7398 298102
rect 6970 297922 7026 297978
rect 7094 297922 7150 297978
rect 7218 297922 7274 297978
rect 7342 297922 7398 297978
rect 6970 280294 7026 280350
rect 7094 280294 7150 280350
rect 7218 280294 7274 280350
rect 7342 280294 7398 280350
rect 6970 280170 7026 280226
rect 7094 280170 7150 280226
rect 7218 280170 7274 280226
rect 7342 280170 7398 280226
rect 6970 280046 7026 280102
rect 7094 280046 7150 280102
rect 7218 280046 7274 280102
rect 7342 280046 7398 280102
rect 6970 279922 7026 279978
rect 7094 279922 7150 279978
rect 7218 279922 7274 279978
rect 7342 279922 7398 279978
rect 6970 262294 7026 262350
rect 7094 262294 7150 262350
rect 7218 262294 7274 262350
rect 7342 262294 7398 262350
rect 6970 262170 7026 262226
rect 7094 262170 7150 262226
rect 7218 262170 7274 262226
rect 7342 262170 7398 262226
rect 6970 262046 7026 262102
rect 7094 262046 7150 262102
rect 7218 262046 7274 262102
rect 7342 262046 7398 262102
rect 6970 261922 7026 261978
rect 7094 261922 7150 261978
rect 7218 261922 7274 261978
rect 7342 261922 7398 261978
rect 6970 244294 7026 244350
rect 7094 244294 7150 244350
rect 7218 244294 7274 244350
rect 7342 244294 7398 244350
rect 6970 244170 7026 244226
rect 7094 244170 7150 244226
rect 7218 244170 7274 244226
rect 7342 244170 7398 244226
rect 6970 244046 7026 244102
rect 7094 244046 7150 244102
rect 7218 244046 7274 244102
rect 7342 244046 7398 244102
rect 6970 243922 7026 243978
rect 7094 243922 7150 243978
rect 7218 243922 7274 243978
rect 7342 243922 7398 243978
rect 6970 226294 7026 226350
rect 7094 226294 7150 226350
rect 7218 226294 7274 226350
rect 7342 226294 7398 226350
rect 6970 226170 7026 226226
rect 7094 226170 7150 226226
rect 7218 226170 7274 226226
rect 7342 226170 7398 226226
rect 6970 226046 7026 226102
rect 7094 226046 7150 226102
rect 7218 226046 7274 226102
rect 7342 226046 7398 226102
rect 6970 225922 7026 225978
rect 7094 225922 7150 225978
rect 7218 225922 7274 225978
rect 7342 225922 7398 225978
rect 6970 208294 7026 208350
rect 7094 208294 7150 208350
rect 7218 208294 7274 208350
rect 7342 208294 7398 208350
rect 6970 208170 7026 208226
rect 7094 208170 7150 208226
rect 7218 208170 7274 208226
rect 7342 208170 7398 208226
rect 6970 208046 7026 208102
rect 7094 208046 7150 208102
rect 7218 208046 7274 208102
rect 7342 208046 7398 208102
rect 6970 207922 7026 207978
rect 7094 207922 7150 207978
rect 7218 207922 7274 207978
rect 7342 207922 7398 207978
rect 6970 190294 7026 190350
rect 7094 190294 7150 190350
rect 7218 190294 7274 190350
rect 7342 190294 7398 190350
rect 6970 190170 7026 190226
rect 7094 190170 7150 190226
rect 7218 190170 7274 190226
rect 7342 190170 7398 190226
rect 6970 190046 7026 190102
rect 7094 190046 7150 190102
rect 7218 190046 7274 190102
rect 7342 190046 7398 190102
rect 6970 189922 7026 189978
rect 7094 189922 7150 189978
rect 7218 189922 7274 189978
rect 7342 189922 7398 189978
rect 6970 172294 7026 172350
rect 7094 172294 7150 172350
rect 7218 172294 7274 172350
rect 7342 172294 7398 172350
rect 6970 172170 7026 172226
rect 7094 172170 7150 172226
rect 7218 172170 7274 172226
rect 7342 172170 7398 172226
rect 6970 172046 7026 172102
rect 7094 172046 7150 172102
rect 7218 172046 7274 172102
rect 7342 172046 7398 172102
rect 6970 171922 7026 171978
rect 7094 171922 7150 171978
rect 7218 171922 7274 171978
rect 7342 171922 7398 171978
rect 6970 154294 7026 154350
rect 7094 154294 7150 154350
rect 7218 154294 7274 154350
rect 7342 154294 7398 154350
rect 6970 154170 7026 154226
rect 7094 154170 7150 154226
rect 7218 154170 7274 154226
rect 7342 154170 7398 154226
rect 6970 154046 7026 154102
rect 7094 154046 7150 154102
rect 7218 154046 7274 154102
rect 7342 154046 7398 154102
rect 6970 153922 7026 153978
rect 7094 153922 7150 153978
rect 7218 153922 7274 153978
rect 7342 153922 7398 153978
rect 6970 136294 7026 136350
rect 7094 136294 7150 136350
rect 7218 136294 7274 136350
rect 7342 136294 7398 136350
rect 6970 136170 7026 136226
rect 7094 136170 7150 136226
rect 7218 136170 7274 136226
rect 7342 136170 7398 136226
rect 6970 136046 7026 136102
rect 7094 136046 7150 136102
rect 7218 136046 7274 136102
rect 7342 136046 7398 136102
rect 6970 135922 7026 135978
rect 7094 135922 7150 135978
rect 7218 135922 7274 135978
rect 7342 135922 7398 135978
rect 6970 118294 7026 118350
rect 7094 118294 7150 118350
rect 7218 118294 7274 118350
rect 7342 118294 7398 118350
rect 6970 118170 7026 118226
rect 7094 118170 7150 118226
rect 7218 118170 7274 118226
rect 7342 118170 7398 118226
rect 6970 118046 7026 118102
rect 7094 118046 7150 118102
rect 7218 118046 7274 118102
rect 7342 118046 7398 118102
rect 6970 117922 7026 117978
rect 7094 117922 7150 117978
rect 7218 117922 7274 117978
rect 7342 117922 7398 117978
rect 6970 100294 7026 100350
rect 7094 100294 7150 100350
rect 7218 100294 7274 100350
rect 7342 100294 7398 100350
rect 6970 100170 7026 100226
rect 7094 100170 7150 100226
rect 7218 100170 7274 100226
rect 7342 100170 7398 100226
rect 6970 100046 7026 100102
rect 7094 100046 7150 100102
rect 7218 100046 7274 100102
rect 7342 100046 7398 100102
rect 6970 99922 7026 99978
rect 7094 99922 7150 99978
rect 7218 99922 7274 99978
rect 7342 99922 7398 99978
rect 6970 82294 7026 82350
rect 7094 82294 7150 82350
rect 7218 82294 7274 82350
rect 7342 82294 7398 82350
rect 6970 82170 7026 82226
rect 7094 82170 7150 82226
rect 7218 82170 7274 82226
rect 7342 82170 7398 82226
rect 6970 82046 7026 82102
rect 7094 82046 7150 82102
rect 7218 82046 7274 82102
rect 7342 82046 7398 82102
rect 6970 81922 7026 81978
rect 7094 81922 7150 81978
rect 7218 81922 7274 81978
rect 7342 81922 7398 81978
rect 6970 64294 7026 64350
rect 7094 64294 7150 64350
rect 7218 64294 7274 64350
rect 7342 64294 7398 64350
rect 6970 64170 7026 64226
rect 7094 64170 7150 64226
rect 7218 64170 7274 64226
rect 7342 64170 7398 64226
rect 6970 64046 7026 64102
rect 7094 64046 7150 64102
rect 7218 64046 7274 64102
rect 7342 64046 7398 64102
rect 6970 63922 7026 63978
rect 7094 63922 7150 63978
rect 7218 63922 7274 63978
rect 7342 63922 7398 63978
rect 6970 46294 7026 46350
rect 7094 46294 7150 46350
rect 7218 46294 7274 46350
rect 7342 46294 7398 46350
rect 6970 46170 7026 46226
rect 7094 46170 7150 46226
rect 7218 46170 7274 46226
rect 7342 46170 7398 46226
rect 6970 46046 7026 46102
rect 7094 46046 7150 46102
rect 7218 46046 7274 46102
rect 7342 46046 7398 46102
rect 6970 45922 7026 45978
rect 7094 45922 7150 45978
rect 7218 45922 7274 45978
rect 7342 45922 7398 45978
rect 6970 28294 7026 28350
rect 7094 28294 7150 28350
rect 7218 28294 7274 28350
rect 7342 28294 7398 28350
rect 6970 28170 7026 28226
rect 7094 28170 7150 28226
rect 7218 28170 7274 28226
rect 7342 28170 7398 28226
rect 6970 28046 7026 28102
rect 7094 28046 7150 28102
rect 7218 28046 7274 28102
rect 7342 28046 7398 28102
rect 6970 27922 7026 27978
rect 7094 27922 7150 27978
rect 7218 27922 7274 27978
rect 7342 27922 7398 27978
rect 21250 580294 21306 580350
rect 21374 580294 21430 580350
rect 21498 580294 21554 580350
rect 21622 580294 21678 580350
rect 21250 580170 21306 580226
rect 21374 580170 21430 580226
rect 21498 580170 21554 580226
rect 21622 580170 21678 580226
rect 21250 580046 21306 580102
rect 21374 580046 21430 580102
rect 21498 580046 21554 580102
rect 21622 580046 21678 580102
rect 21250 579922 21306 579978
rect 21374 579922 21430 579978
rect 21498 579922 21554 579978
rect 21622 579922 21678 579978
rect 21250 562294 21306 562350
rect 21374 562294 21430 562350
rect 21498 562294 21554 562350
rect 21622 562294 21678 562350
rect 21250 562170 21306 562226
rect 21374 562170 21430 562226
rect 21498 562170 21554 562226
rect 21622 562170 21678 562226
rect 21250 562046 21306 562102
rect 21374 562046 21430 562102
rect 21498 562046 21554 562102
rect 21622 562046 21678 562102
rect 21250 561922 21306 561978
rect 21374 561922 21430 561978
rect 21498 561922 21554 561978
rect 21622 561922 21678 561978
rect 21250 544294 21306 544350
rect 21374 544294 21430 544350
rect 21498 544294 21554 544350
rect 21622 544294 21678 544350
rect 21250 544170 21306 544226
rect 21374 544170 21430 544226
rect 21498 544170 21554 544226
rect 21622 544170 21678 544226
rect 21250 544046 21306 544102
rect 21374 544046 21430 544102
rect 21498 544046 21554 544102
rect 21622 544046 21678 544102
rect 21250 543922 21306 543978
rect 21374 543922 21430 543978
rect 21498 543922 21554 543978
rect 21622 543922 21678 543978
rect 21250 526294 21306 526350
rect 21374 526294 21430 526350
rect 21498 526294 21554 526350
rect 21622 526294 21678 526350
rect 21250 526170 21306 526226
rect 21374 526170 21430 526226
rect 21498 526170 21554 526226
rect 21622 526170 21678 526226
rect 21250 526046 21306 526102
rect 21374 526046 21430 526102
rect 21498 526046 21554 526102
rect 21622 526046 21678 526102
rect 21250 525922 21306 525978
rect 21374 525922 21430 525978
rect 21498 525922 21554 525978
rect 21622 525922 21678 525978
rect 21250 508294 21306 508350
rect 21374 508294 21430 508350
rect 21498 508294 21554 508350
rect 21622 508294 21678 508350
rect 21250 508170 21306 508226
rect 21374 508170 21430 508226
rect 21498 508170 21554 508226
rect 21622 508170 21678 508226
rect 21250 508046 21306 508102
rect 21374 508046 21430 508102
rect 21498 508046 21554 508102
rect 21622 508046 21678 508102
rect 21250 507922 21306 507978
rect 21374 507922 21430 507978
rect 21498 507922 21554 507978
rect 21622 507922 21678 507978
rect 21250 490294 21306 490350
rect 21374 490294 21430 490350
rect 21498 490294 21554 490350
rect 21622 490294 21678 490350
rect 21250 490170 21306 490226
rect 21374 490170 21430 490226
rect 21498 490170 21554 490226
rect 21622 490170 21678 490226
rect 21250 490046 21306 490102
rect 21374 490046 21430 490102
rect 21498 490046 21554 490102
rect 21622 490046 21678 490102
rect 21250 489922 21306 489978
rect 21374 489922 21430 489978
rect 21498 489922 21554 489978
rect 21622 489922 21678 489978
rect 21250 472294 21306 472350
rect 21374 472294 21430 472350
rect 21498 472294 21554 472350
rect 21622 472294 21678 472350
rect 21250 472170 21306 472226
rect 21374 472170 21430 472226
rect 21498 472170 21554 472226
rect 21622 472170 21678 472226
rect 21250 472046 21306 472102
rect 21374 472046 21430 472102
rect 21498 472046 21554 472102
rect 21622 472046 21678 472102
rect 21250 471922 21306 471978
rect 21374 471922 21430 471978
rect 21498 471922 21554 471978
rect 21622 471922 21678 471978
rect 24970 598116 25026 598172
rect 25094 598116 25150 598172
rect 25218 598116 25274 598172
rect 25342 598116 25398 598172
rect 24970 597992 25026 598048
rect 25094 597992 25150 598048
rect 25218 597992 25274 598048
rect 25342 597992 25398 598048
rect 24970 597868 25026 597924
rect 25094 597868 25150 597924
rect 25218 597868 25274 597924
rect 25342 597868 25398 597924
rect 24970 597744 25026 597800
rect 25094 597744 25150 597800
rect 25218 597744 25274 597800
rect 25342 597744 25398 597800
rect 24970 586294 25026 586350
rect 25094 586294 25150 586350
rect 25218 586294 25274 586350
rect 25342 586294 25398 586350
rect 24970 586170 25026 586226
rect 25094 586170 25150 586226
rect 25218 586170 25274 586226
rect 25342 586170 25398 586226
rect 24970 586046 25026 586102
rect 25094 586046 25150 586102
rect 25218 586046 25274 586102
rect 25342 586046 25398 586102
rect 24970 585922 25026 585978
rect 25094 585922 25150 585978
rect 25218 585922 25274 585978
rect 25342 585922 25398 585978
rect 24970 568294 25026 568350
rect 25094 568294 25150 568350
rect 25218 568294 25274 568350
rect 25342 568294 25398 568350
rect 24970 568170 25026 568226
rect 25094 568170 25150 568226
rect 25218 568170 25274 568226
rect 25342 568170 25398 568226
rect 24970 568046 25026 568102
rect 25094 568046 25150 568102
rect 25218 568046 25274 568102
rect 25342 568046 25398 568102
rect 24970 567922 25026 567978
rect 25094 567922 25150 567978
rect 25218 567922 25274 567978
rect 25342 567922 25398 567978
rect 24970 550294 25026 550350
rect 25094 550294 25150 550350
rect 25218 550294 25274 550350
rect 25342 550294 25398 550350
rect 24970 550170 25026 550226
rect 25094 550170 25150 550226
rect 25218 550170 25274 550226
rect 25342 550170 25398 550226
rect 24970 550046 25026 550102
rect 25094 550046 25150 550102
rect 25218 550046 25274 550102
rect 25342 550046 25398 550102
rect 24970 549922 25026 549978
rect 25094 549922 25150 549978
rect 25218 549922 25274 549978
rect 25342 549922 25398 549978
rect 24970 532294 25026 532350
rect 25094 532294 25150 532350
rect 25218 532294 25274 532350
rect 25342 532294 25398 532350
rect 24970 532170 25026 532226
rect 25094 532170 25150 532226
rect 25218 532170 25274 532226
rect 25342 532170 25398 532226
rect 24970 532046 25026 532102
rect 25094 532046 25150 532102
rect 25218 532046 25274 532102
rect 25342 532046 25398 532102
rect 24970 531922 25026 531978
rect 25094 531922 25150 531978
rect 25218 531922 25274 531978
rect 25342 531922 25398 531978
rect 24970 514294 25026 514350
rect 25094 514294 25150 514350
rect 25218 514294 25274 514350
rect 25342 514294 25398 514350
rect 24970 514170 25026 514226
rect 25094 514170 25150 514226
rect 25218 514170 25274 514226
rect 25342 514170 25398 514226
rect 24970 514046 25026 514102
rect 25094 514046 25150 514102
rect 25218 514046 25274 514102
rect 25342 514046 25398 514102
rect 24970 513922 25026 513978
rect 25094 513922 25150 513978
rect 25218 513922 25274 513978
rect 25342 513922 25398 513978
rect 24970 496294 25026 496350
rect 25094 496294 25150 496350
rect 25218 496294 25274 496350
rect 25342 496294 25398 496350
rect 24970 496170 25026 496226
rect 25094 496170 25150 496226
rect 25218 496170 25274 496226
rect 25342 496170 25398 496226
rect 24970 496046 25026 496102
rect 25094 496046 25150 496102
rect 25218 496046 25274 496102
rect 25342 496046 25398 496102
rect 24970 495922 25026 495978
rect 25094 495922 25150 495978
rect 25218 495922 25274 495978
rect 25342 495922 25398 495978
rect 24970 478294 25026 478350
rect 25094 478294 25150 478350
rect 25218 478294 25274 478350
rect 25342 478294 25398 478350
rect 24970 478170 25026 478226
rect 25094 478170 25150 478226
rect 25218 478170 25274 478226
rect 25342 478170 25398 478226
rect 24970 478046 25026 478102
rect 25094 478046 25150 478102
rect 25218 478046 25274 478102
rect 25342 478046 25398 478102
rect 24970 477922 25026 477978
rect 25094 477922 25150 477978
rect 25218 477922 25274 477978
rect 25342 477922 25398 477978
rect 24970 460294 25026 460350
rect 25094 460294 25150 460350
rect 25218 460294 25274 460350
rect 25342 460294 25398 460350
rect 24970 460170 25026 460226
rect 25094 460170 25150 460226
rect 25218 460170 25274 460226
rect 25342 460170 25398 460226
rect 24970 460046 25026 460102
rect 25094 460046 25150 460102
rect 25218 460046 25274 460102
rect 25342 460046 25398 460102
rect 24970 459922 25026 459978
rect 25094 459922 25150 459978
rect 25218 459922 25274 459978
rect 25342 459922 25398 459978
rect 39250 597156 39306 597212
rect 39374 597156 39430 597212
rect 39498 597156 39554 597212
rect 39622 597156 39678 597212
rect 39250 597032 39306 597088
rect 39374 597032 39430 597088
rect 39498 597032 39554 597088
rect 39622 597032 39678 597088
rect 39250 596908 39306 596964
rect 39374 596908 39430 596964
rect 39498 596908 39554 596964
rect 39622 596908 39678 596964
rect 39250 596784 39306 596840
rect 39374 596784 39430 596840
rect 39498 596784 39554 596840
rect 39622 596784 39678 596840
rect 39250 580294 39306 580350
rect 39374 580294 39430 580350
rect 39498 580294 39554 580350
rect 39622 580294 39678 580350
rect 39250 580170 39306 580226
rect 39374 580170 39430 580226
rect 39498 580170 39554 580226
rect 39622 580170 39678 580226
rect 39250 580046 39306 580102
rect 39374 580046 39430 580102
rect 39498 580046 39554 580102
rect 39622 580046 39678 580102
rect 39250 579922 39306 579978
rect 39374 579922 39430 579978
rect 39498 579922 39554 579978
rect 39622 579922 39678 579978
rect 39250 562294 39306 562350
rect 39374 562294 39430 562350
rect 39498 562294 39554 562350
rect 39622 562294 39678 562350
rect 39250 562170 39306 562226
rect 39374 562170 39430 562226
rect 39498 562170 39554 562226
rect 39622 562170 39678 562226
rect 39250 562046 39306 562102
rect 39374 562046 39430 562102
rect 39498 562046 39554 562102
rect 39622 562046 39678 562102
rect 39250 561922 39306 561978
rect 39374 561922 39430 561978
rect 39498 561922 39554 561978
rect 39622 561922 39678 561978
rect 39250 544294 39306 544350
rect 39374 544294 39430 544350
rect 39498 544294 39554 544350
rect 39622 544294 39678 544350
rect 39250 544170 39306 544226
rect 39374 544170 39430 544226
rect 39498 544170 39554 544226
rect 39622 544170 39678 544226
rect 39250 544046 39306 544102
rect 39374 544046 39430 544102
rect 39498 544046 39554 544102
rect 39622 544046 39678 544102
rect 39250 543922 39306 543978
rect 39374 543922 39430 543978
rect 39498 543922 39554 543978
rect 39622 543922 39678 543978
rect 39250 526294 39306 526350
rect 39374 526294 39430 526350
rect 39498 526294 39554 526350
rect 39622 526294 39678 526350
rect 39250 526170 39306 526226
rect 39374 526170 39430 526226
rect 39498 526170 39554 526226
rect 39622 526170 39678 526226
rect 39250 526046 39306 526102
rect 39374 526046 39430 526102
rect 39498 526046 39554 526102
rect 39622 526046 39678 526102
rect 39250 525922 39306 525978
rect 39374 525922 39430 525978
rect 39498 525922 39554 525978
rect 39622 525922 39678 525978
rect 39250 508294 39306 508350
rect 39374 508294 39430 508350
rect 39498 508294 39554 508350
rect 39622 508294 39678 508350
rect 39250 508170 39306 508226
rect 39374 508170 39430 508226
rect 39498 508170 39554 508226
rect 39622 508170 39678 508226
rect 39250 508046 39306 508102
rect 39374 508046 39430 508102
rect 39498 508046 39554 508102
rect 39622 508046 39678 508102
rect 39250 507922 39306 507978
rect 39374 507922 39430 507978
rect 39498 507922 39554 507978
rect 39622 507922 39678 507978
rect 39250 490294 39306 490350
rect 39374 490294 39430 490350
rect 39498 490294 39554 490350
rect 39622 490294 39678 490350
rect 39250 490170 39306 490226
rect 39374 490170 39430 490226
rect 39498 490170 39554 490226
rect 39622 490170 39678 490226
rect 39250 490046 39306 490102
rect 39374 490046 39430 490102
rect 39498 490046 39554 490102
rect 39622 490046 39678 490102
rect 39250 489922 39306 489978
rect 39374 489922 39430 489978
rect 39498 489922 39554 489978
rect 39622 489922 39678 489978
rect 39250 472294 39306 472350
rect 39374 472294 39430 472350
rect 39498 472294 39554 472350
rect 39622 472294 39678 472350
rect 39250 472170 39306 472226
rect 39374 472170 39430 472226
rect 39498 472170 39554 472226
rect 39622 472170 39678 472226
rect 39250 472046 39306 472102
rect 39374 472046 39430 472102
rect 39498 472046 39554 472102
rect 39622 472046 39678 472102
rect 39250 471922 39306 471978
rect 39374 471922 39430 471978
rect 39498 471922 39554 471978
rect 39622 471922 39678 471978
rect 42970 598116 43026 598172
rect 43094 598116 43150 598172
rect 43218 598116 43274 598172
rect 43342 598116 43398 598172
rect 42970 597992 43026 598048
rect 43094 597992 43150 598048
rect 43218 597992 43274 598048
rect 43342 597992 43398 598048
rect 42970 597868 43026 597924
rect 43094 597868 43150 597924
rect 43218 597868 43274 597924
rect 43342 597868 43398 597924
rect 42970 597744 43026 597800
rect 43094 597744 43150 597800
rect 43218 597744 43274 597800
rect 43342 597744 43398 597800
rect 42970 586294 43026 586350
rect 43094 586294 43150 586350
rect 43218 586294 43274 586350
rect 43342 586294 43398 586350
rect 42970 586170 43026 586226
rect 43094 586170 43150 586226
rect 43218 586170 43274 586226
rect 43342 586170 43398 586226
rect 42970 586046 43026 586102
rect 43094 586046 43150 586102
rect 43218 586046 43274 586102
rect 43342 586046 43398 586102
rect 42970 585922 43026 585978
rect 43094 585922 43150 585978
rect 43218 585922 43274 585978
rect 43342 585922 43398 585978
rect 42970 568294 43026 568350
rect 43094 568294 43150 568350
rect 43218 568294 43274 568350
rect 43342 568294 43398 568350
rect 42970 568170 43026 568226
rect 43094 568170 43150 568226
rect 43218 568170 43274 568226
rect 43342 568170 43398 568226
rect 42970 568046 43026 568102
rect 43094 568046 43150 568102
rect 43218 568046 43274 568102
rect 43342 568046 43398 568102
rect 42970 567922 43026 567978
rect 43094 567922 43150 567978
rect 43218 567922 43274 567978
rect 43342 567922 43398 567978
rect 42970 550294 43026 550350
rect 43094 550294 43150 550350
rect 43218 550294 43274 550350
rect 43342 550294 43398 550350
rect 42970 550170 43026 550226
rect 43094 550170 43150 550226
rect 43218 550170 43274 550226
rect 43342 550170 43398 550226
rect 42970 550046 43026 550102
rect 43094 550046 43150 550102
rect 43218 550046 43274 550102
rect 43342 550046 43398 550102
rect 42970 549922 43026 549978
rect 43094 549922 43150 549978
rect 43218 549922 43274 549978
rect 43342 549922 43398 549978
rect 42970 532294 43026 532350
rect 43094 532294 43150 532350
rect 43218 532294 43274 532350
rect 43342 532294 43398 532350
rect 42970 532170 43026 532226
rect 43094 532170 43150 532226
rect 43218 532170 43274 532226
rect 43342 532170 43398 532226
rect 42970 532046 43026 532102
rect 43094 532046 43150 532102
rect 43218 532046 43274 532102
rect 43342 532046 43398 532102
rect 42970 531922 43026 531978
rect 43094 531922 43150 531978
rect 43218 531922 43274 531978
rect 43342 531922 43398 531978
rect 42970 514294 43026 514350
rect 43094 514294 43150 514350
rect 43218 514294 43274 514350
rect 43342 514294 43398 514350
rect 42970 514170 43026 514226
rect 43094 514170 43150 514226
rect 43218 514170 43274 514226
rect 43342 514170 43398 514226
rect 42970 514046 43026 514102
rect 43094 514046 43150 514102
rect 43218 514046 43274 514102
rect 43342 514046 43398 514102
rect 42970 513922 43026 513978
rect 43094 513922 43150 513978
rect 43218 513922 43274 513978
rect 43342 513922 43398 513978
rect 42970 496294 43026 496350
rect 43094 496294 43150 496350
rect 43218 496294 43274 496350
rect 43342 496294 43398 496350
rect 42970 496170 43026 496226
rect 43094 496170 43150 496226
rect 43218 496170 43274 496226
rect 43342 496170 43398 496226
rect 42970 496046 43026 496102
rect 43094 496046 43150 496102
rect 43218 496046 43274 496102
rect 43342 496046 43398 496102
rect 42970 495922 43026 495978
rect 43094 495922 43150 495978
rect 43218 495922 43274 495978
rect 43342 495922 43398 495978
rect 42970 478294 43026 478350
rect 43094 478294 43150 478350
rect 43218 478294 43274 478350
rect 43342 478294 43398 478350
rect 42970 478170 43026 478226
rect 43094 478170 43150 478226
rect 43218 478170 43274 478226
rect 43342 478170 43398 478226
rect 42970 478046 43026 478102
rect 43094 478046 43150 478102
rect 43218 478046 43274 478102
rect 43342 478046 43398 478102
rect 42970 477922 43026 477978
rect 43094 477922 43150 477978
rect 43218 477922 43274 477978
rect 43342 477922 43398 477978
rect 42970 460294 43026 460350
rect 43094 460294 43150 460350
rect 43218 460294 43274 460350
rect 43342 460294 43398 460350
rect 42970 460170 43026 460226
rect 43094 460170 43150 460226
rect 43218 460170 43274 460226
rect 43342 460170 43398 460226
rect 42970 460046 43026 460102
rect 43094 460046 43150 460102
rect 43218 460046 43274 460102
rect 43342 460046 43398 460102
rect 42970 459922 43026 459978
rect 43094 459922 43150 459978
rect 43218 459922 43274 459978
rect 43342 459922 43398 459978
rect 57250 597156 57306 597212
rect 57374 597156 57430 597212
rect 57498 597156 57554 597212
rect 57622 597156 57678 597212
rect 57250 597032 57306 597088
rect 57374 597032 57430 597088
rect 57498 597032 57554 597088
rect 57622 597032 57678 597088
rect 57250 596908 57306 596964
rect 57374 596908 57430 596964
rect 57498 596908 57554 596964
rect 57622 596908 57678 596964
rect 57250 596784 57306 596840
rect 57374 596784 57430 596840
rect 57498 596784 57554 596840
rect 57622 596784 57678 596840
rect 57250 580294 57306 580350
rect 57374 580294 57430 580350
rect 57498 580294 57554 580350
rect 57622 580294 57678 580350
rect 57250 580170 57306 580226
rect 57374 580170 57430 580226
rect 57498 580170 57554 580226
rect 57622 580170 57678 580226
rect 57250 580046 57306 580102
rect 57374 580046 57430 580102
rect 57498 580046 57554 580102
rect 57622 580046 57678 580102
rect 57250 579922 57306 579978
rect 57374 579922 57430 579978
rect 57498 579922 57554 579978
rect 57622 579922 57678 579978
rect 57250 562294 57306 562350
rect 57374 562294 57430 562350
rect 57498 562294 57554 562350
rect 57622 562294 57678 562350
rect 57250 562170 57306 562226
rect 57374 562170 57430 562226
rect 57498 562170 57554 562226
rect 57622 562170 57678 562226
rect 57250 562046 57306 562102
rect 57374 562046 57430 562102
rect 57498 562046 57554 562102
rect 57622 562046 57678 562102
rect 57250 561922 57306 561978
rect 57374 561922 57430 561978
rect 57498 561922 57554 561978
rect 57622 561922 57678 561978
rect 57250 544294 57306 544350
rect 57374 544294 57430 544350
rect 57498 544294 57554 544350
rect 57622 544294 57678 544350
rect 57250 544170 57306 544226
rect 57374 544170 57430 544226
rect 57498 544170 57554 544226
rect 57622 544170 57678 544226
rect 57250 544046 57306 544102
rect 57374 544046 57430 544102
rect 57498 544046 57554 544102
rect 57622 544046 57678 544102
rect 57250 543922 57306 543978
rect 57374 543922 57430 543978
rect 57498 543922 57554 543978
rect 57622 543922 57678 543978
rect 57250 526294 57306 526350
rect 57374 526294 57430 526350
rect 57498 526294 57554 526350
rect 57622 526294 57678 526350
rect 57250 526170 57306 526226
rect 57374 526170 57430 526226
rect 57498 526170 57554 526226
rect 57622 526170 57678 526226
rect 57250 526046 57306 526102
rect 57374 526046 57430 526102
rect 57498 526046 57554 526102
rect 57622 526046 57678 526102
rect 57250 525922 57306 525978
rect 57374 525922 57430 525978
rect 57498 525922 57554 525978
rect 57622 525922 57678 525978
rect 57250 508294 57306 508350
rect 57374 508294 57430 508350
rect 57498 508294 57554 508350
rect 57622 508294 57678 508350
rect 57250 508170 57306 508226
rect 57374 508170 57430 508226
rect 57498 508170 57554 508226
rect 57622 508170 57678 508226
rect 57250 508046 57306 508102
rect 57374 508046 57430 508102
rect 57498 508046 57554 508102
rect 57622 508046 57678 508102
rect 57250 507922 57306 507978
rect 57374 507922 57430 507978
rect 57498 507922 57554 507978
rect 57622 507922 57678 507978
rect 57250 490294 57306 490350
rect 57374 490294 57430 490350
rect 57498 490294 57554 490350
rect 57622 490294 57678 490350
rect 57250 490170 57306 490226
rect 57374 490170 57430 490226
rect 57498 490170 57554 490226
rect 57622 490170 57678 490226
rect 57250 490046 57306 490102
rect 57374 490046 57430 490102
rect 57498 490046 57554 490102
rect 57622 490046 57678 490102
rect 57250 489922 57306 489978
rect 57374 489922 57430 489978
rect 57498 489922 57554 489978
rect 57622 489922 57678 489978
rect 57250 472294 57306 472350
rect 57374 472294 57430 472350
rect 57498 472294 57554 472350
rect 57622 472294 57678 472350
rect 57250 472170 57306 472226
rect 57374 472170 57430 472226
rect 57498 472170 57554 472226
rect 57622 472170 57678 472226
rect 57250 472046 57306 472102
rect 57374 472046 57430 472102
rect 57498 472046 57554 472102
rect 57622 472046 57678 472102
rect 57250 471922 57306 471978
rect 57374 471922 57430 471978
rect 57498 471922 57554 471978
rect 57622 471922 57678 471978
rect 60970 598116 61026 598172
rect 61094 598116 61150 598172
rect 61218 598116 61274 598172
rect 61342 598116 61398 598172
rect 60970 597992 61026 598048
rect 61094 597992 61150 598048
rect 61218 597992 61274 598048
rect 61342 597992 61398 598048
rect 60970 597868 61026 597924
rect 61094 597868 61150 597924
rect 61218 597868 61274 597924
rect 61342 597868 61398 597924
rect 60970 597744 61026 597800
rect 61094 597744 61150 597800
rect 61218 597744 61274 597800
rect 61342 597744 61398 597800
rect 60970 586294 61026 586350
rect 61094 586294 61150 586350
rect 61218 586294 61274 586350
rect 61342 586294 61398 586350
rect 60970 586170 61026 586226
rect 61094 586170 61150 586226
rect 61218 586170 61274 586226
rect 61342 586170 61398 586226
rect 60970 586046 61026 586102
rect 61094 586046 61150 586102
rect 61218 586046 61274 586102
rect 61342 586046 61398 586102
rect 60970 585922 61026 585978
rect 61094 585922 61150 585978
rect 61218 585922 61274 585978
rect 61342 585922 61398 585978
rect 60970 568294 61026 568350
rect 61094 568294 61150 568350
rect 61218 568294 61274 568350
rect 61342 568294 61398 568350
rect 60970 568170 61026 568226
rect 61094 568170 61150 568226
rect 61218 568170 61274 568226
rect 61342 568170 61398 568226
rect 60970 568046 61026 568102
rect 61094 568046 61150 568102
rect 61218 568046 61274 568102
rect 61342 568046 61398 568102
rect 60970 567922 61026 567978
rect 61094 567922 61150 567978
rect 61218 567922 61274 567978
rect 61342 567922 61398 567978
rect 60970 550294 61026 550350
rect 61094 550294 61150 550350
rect 61218 550294 61274 550350
rect 61342 550294 61398 550350
rect 60970 550170 61026 550226
rect 61094 550170 61150 550226
rect 61218 550170 61274 550226
rect 61342 550170 61398 550226
rect 60970 550046 61026 550102
rect 61094 550046 61150 550102
rect 61218 550046 61274 550102
rect 61342 550046 61398 550102
rect 60970 549922 61026 549978
rect 61094 549922 61150 549978
rect 61218 549922 61274 549978
rect 61342 549922 61398 549978
rect 60970 532294 61026 532350
rect 61094 532294 61150 532350
rect 61218 532294 61274 532350
rect 61342 532294 61398 532350
rect 60970 532170 61026 532226
rect 61094 532170 61150 532226
rect 61218 532170 61274 532226
rect 61342 532170 61398 532226
rect 60970 532046 61026 532102
rect 61094 532046 61150 532102
rect 61218 532046 61274 532102
rect 61342 532046 61398 532102
rect 60970 531922 61026 531978
rect 61094 531922 61150 531978
rect 61218 531922 61274 531978
rect 61342 531922 61398 531978
rect 60970 514294 61026 514350
rect 61094 514294 61150 514350
rect 61218 514294 61274 514350
rect 61342 514294 61398 514350
rect 60970 514170 61026 514226
rect 61094 514170 61150 514226
rect 61218 514170 61274 514226
rect 61342 514170 61398 514226
rect 60970 514046 61026 514102
rect 61094 514046 61150 514102
rect 61218 514046 61274 514102
rect 61342 514046 61398 514102
rect 60970 513922 61026 513978
rect 61094 513922 61150 513978
rect 61218 513922 61274 513978
rect 61342 513922 61398 513978
rect 60970 496294 61026 496350
rect 61094 496294 61150 496350
rect 61218 496294 61274 496350
rect 61342 496294 61398 496350
rect 60970 496170 61026 496226
rect 61094 496170 61150 496226
rect 61218 496170 61274 496226
rect 61342 496170 61398 496226
rect 60970 496046 61026 496102
rect 61094 496046 61150 496102
rect 61218 496046 61274 496102
rect 61342 496046 61398 496102
rect 60970 495922 61026 495978
rect 61094 495922 61150 495978
rect 61218 495922 61274 495978
rect 61342 495922 61398 495978
rect 60970 478294 61026 478350
rect 61094 478294 61150 478350
rect 61218 478294 61274 478350
rect 61342 478294 61398 478350
rect 60970 478170 61026 478226
rect 61094 478170 61150 478226
rect 61218 478170 61274 478226
rect 61342 478170 61398 478226
rect 60970 478046 61026 478102
rect 61094 478046 61150 478102
rect 61218 478046 61274 478102
rect 61342 478046 61398 478102
rect 60970 477922 61026 477978
rect 61094 477922 61150 477978
rect 61218 477922 61274 477978
rect 61342 477922 61398 477978
rect 60970 460294 61026 460350
rect 61094 460294 61150 460350
rect 61218 460294 61274 460350
rect 61342 460294 61398 460350
rect 60970 460170 61026 460226
rect 61094 460170 61150 460226
rect 61218 460170 61274 460226
rect 61342 460170 61398 460226
rect 60970 460046 61026 460102
rect 61094 460046 61150 460102
rect 61218 460046 61274 460102
rect 61342 460046 61398 460102
rect 60970 459922 61026 459978
rect 61094 459922 61150 459978
rect 61218 459922 61274 459978
rect 61342 459922 61398 459978
rect 75250 597156 75306 597212
rect 75374 597156 75430 597212
rect 75498 597156 75554 597212
rect 75622 597156 75678 597212
rect 75250 597032 75306 597088
rect 75374 597032 75430 597088
rect 75498 597032 75554 597088
rect 75622 597032 75678 597088
rect 75250 596908 75306 596964
rect 75374 596908 75430 596964
rect 75498 596908 75554 596964
rect 75622 596908 75678 596964
rect 75250 596784 75306 596840
rect 75374 596784 75430 596840
rect 75498 596784 75554 596840
rect 75622 596784 75678 596840
rect 75250 580294 75306 580350
rect 75374 580294 75430 580350
rect 75498 580294 75554 580350
rect 75622 580294 75678 580350
rect 75250 580170 75306 580226
rect 75374 580170 75430 580226
rect 75498 580170 75554 580226
rect 75622 580170 75678 580226
rect 75250 580046 75306 580102
rect 75374 580046 75430 580102
rect 75498 580046 75554 580102
rect 75622 580046 75678 580102
rect 75250 579922 75306 579978
rect 75374 579922 75430 579978
rect 75498 579922 75554 579978
rect 75622 579922 75678 579978
rect 75250 562294 75306 562350
rect 75374 562294 75430 562350
rect 75498 562294 75554 562350
rect 75622 562294 75678 562350
rect 75250 562170 75306 562226
rect 75374 562170 75430 562226
rect 75498 562170 75554 562226
rect 75622 562170 75678 562226
rect 75250 562046 75306 562102
rect 75374 562046 75430 562102
rect 75498 562046 75554 562102
rect 75622 562046 75678 562102
rect 75250 561922 75306 561978
rect 75374 561922 75430 561978
rect 75498 561922 75554 561978
rect 75622 561922 75678 561978
rect 75250 544294 75306 544350
rect 75374 544294 75430 544350
rect 75498 544294 75554 544350
rect 75622 544294 75678 544350
rect 75250 544170 75306 544226
rect 75374 544170 75430 544226
rect 75498 544170 75554 544226
rect 75622 544170 75678 544226
rect 75250 544046 75306 544102
rect 75374 544046 75430 544102
rect 75498 544046 75554 544102
rect 75622 544046 75678 544102
rect 75250 543922 75306 543978
rect 75374 543922 75430 543978
rect 75498 543922 75554 543978
rect 75622 543922 75678 543978
rect 75250 526294 75306 526350
rect 75374 526294 75430 526350
rect 75498 526294 75554 526350
rect 75622 526294 75678 526350
rect 75250 526170 75306 526226
rect 75374 526170 75430 526226
rect 75498 526170 75554 526226
rect 75622 526170 75678 526226
rect 75250 526046 75306 526102
rect 75374 526046 75430 526102
rect 75498 526046 75554 526102
rect 75622 526046 75678 526102
rect 75250 525922 75306 525978
rect 75374 525922 75430 525978
rect 75498 525922 75554 525978
rect 75622 525922 75678 525978
rect 75250 508294 75306 508350
rect 75374 508294 75430 508350
rect 75498 508294 75554 508350
rect 75622 508294 75678 508350
rect 75250 508170 75306 508226
rect 75374 508170 75430 508226
rect 75498 508170 75554 508226
rect 75622 508170 75678 508226
rect 75250 508046 75306 508102
rect 75374 508046 75430 508102
rect 75498 508046 75554 508102
rect 75622 508046 75678 508102
rect 75250 507922 75306 507978
rect 75374 507922 75430 507978
rect 75498 507922 75554 507978
rect 75622 507922 75678 507978
rect 75250 490294 75306 490350
rect 75374 490294 75430 490350
rect 75498 490294 75554 490350
rect 75622 490294 75678 490350
rect 75250 490170 75306 490226
rect 75374 490170 75430 490226
rect 75498 490170 75554 490226
rect 75622 490170 75678 490226
rect 75250 490046 75306 490102
rect 75374 490046 75430 490102
rect 75498 490046 75554 490102
rect 75622 490046 75678 490102
rect 75250 489922 75306 489978
rect 75374 489922 75430 489978
rect 75498 489922 75554 489978
rect 75622 489922 75678 489978
rect 75250 472294 75306 472350
rect 75374 472294 75430 472350
rect 75498 472294 75554 472350
rect 75622 472294 75678 472350
rect 75250 472170 75306 472226
rect 75374 472170 75430 472226
rect 75498 472170 75554 472226
rect 75622 472170 75678 472226
rect 75250 472046 75306 472102
rect 75374 472046 75430 472102
rect 75498 472046 75554 472102
rect 75622 472046 75678 472102
rect 75250 471922 75306 471978
rect 75374 471922 75430 471978
rect 75498 471922 75554 471978
rect 75622 471922 75678 471978
rect 78970 598116 79026 598172
rect 79094 598116 79150 598172
rect 79218 598116 79274 598172
rect 79342 598116 79398 598172
rect 78970 597992 79026 598048
rect 79094 597992 79150 598048
rect 79218 597992 79274 598048
rect 79342 597992 79398 598048
rect 78970 597868 79026 597924
rect 79094 597868 79150 597924
rect 79218 597868 79274 597924
rect 79342 597868 79398 597924
rect 78970 597744 79026 597800
rect 79094 597744 79150 597800
rect 79218 597744 79274 597800
rect 79342 597744 79398 597800
rect 78970 586294 79026 586350
rect 79094 586294 79150 586350
rect 79218 586294 79274 586350
rect 79342 586294 79398 586350
rect 78970 586170 79026 586226
rect 79094 586170 79150 586226
rect 79218 586170 79274 586226
rect 79342 586170 79398 586226
rect 78970 586046 79026 586102
rect 79094 586046 79150 586102
rect 79218 586046 79274 586102
rect 79342 586046 79398 586102
rect 78970 585922 79026 585978
rect 79094 585922 79150 585978
rect 79218 585922 79274 585978
rect 79342 585922 79398 585978
rect 78970 568294 79026 568350
rect 79094 568294 79150 568350
rect 79218 568294 79274 568350
rect 79342 568294 79398 568350
rect 78970 568170 79026 568226
rect 79094 568170 79150 568226
rect 79218 568170 79274 568226
rect 79342 568170 79398 568226
rect 78970 568046 79026 568102
rect 79094 568046 79150 568102
rect 79218 568046 79274 568102
rect 79342 568046 79398 568102
rect 78970 567922 79026 567978
rect 79094 567922 79150 567978
rect 79218 567922 79274 567978
rect 79342 567922 79398 567978
rect 78970 550294 79026 550350
rect 79094 550294 79150 550350
rect 79218 550294 79274 550350
rect 79342 550294 79398 550350
rect 78970 550170 79026 550226
rect 79094 550170 79150 550226
rect 79218 550170 79274 550226
rect 79342 550170 79398 550226
rect 78970 550046 79026 550102
rect 79094 550046 79150 550102
rect 79218 550046 79274 550102
rect 79342 550046 79398 550102
rect 78970 549922 79026 549978
rect 79094 549922 79150 549978
rect 79218 549922 79274 549978
rect 79342 549922 79398 549978
rect 78970 532294 79026 532350
rect 79094 532294 79150 532350
rect 79218 532294 79274 532350
rect 79342 532294 79398 532350
rect 78970 532170 79026 532226
rect 79094 532170 79150 532226
rect 79218 532170 79274 532226
rect 79342 532170 79398 532226
rect 78970 532046 79026 532102
rect 79094 532046 79150 532102
rect 79218 532046 79274 532102
rect 79342 532046 79398 532102
rect 78970 531922 79026 531978
rect 79094 531922 79150 531978
rect 79218 531922 79274 531978
rect 79342 531922 79398 531978
rect 78970 514294 79026 514350
rect 79094 514294 79150 514350
rect 79218 514294 79274 514350
rect 79342 514294 79398 514350
rect 78970 514170 79026 514226
rect 79094 514170 79150 514226
rect 79218 514170 79274 514226
rect 79342 514170 79398 514226
rect 78970 514046 79026 514102
rect 79094 514046 79150 514102
rect 79218 514046 79274 514102
rect 79342 514046 79398 514102
rect 78970 513922 79026 513978
rect 79094 513922 79150 513978
rect 79218 513922 79274 513978
rect 79342 513922 79398 513978
rect 78970 496294 79026 496350
rect 79094 496294 79150 496350
rect 79218 496294 79274 496350
rect 79342 496294 79398 496350
rect 78970 496170 79026 496226
rect 79094 496170 79150 496226
rect 79218 496170 79274 496226
rect 79342 496170 79398 496226
rect 78970 496046 79026 496102
rect 79094 496046 79150 496102
rect 79218 496046 79274 496102
rect 79342 496046 79398 496102
rect 78970 495922 79026 495978
rect 79094 495922 79150 495978
rect 79218 495922 79274 495978
rect 79342 495922 79398 495978
rect 78970 478294 79026 478350
rect 79094 478294 79150 478350
rect 79218 478294 79274 478350
rect 79342 478294 79398 478350
rect 78970 478170 79026 478226
rect 79094 478170 79150 478226
rect 79218 478170 79274 478226
rect 79342 478170 79398 478226
rect 78970 478046 79026 478102
rect 79094 478046 79150 478102
rect 79218 478046 79274 478102
rect 79342 478046 79398 478102
rect 78970 477922 79026 477978
rect 79094 477922 79150 477978
rect 79218 477922 79274 477978
rect 79342 477922 79398 477978
rect 78970 460294 79026 460350
rect 79094 460294 79150 460350
rect 79218 460294 79274 460350
rect 79342 460294 79398 460350
rect 78970 460170 79026 460226
rect 79094 460170 79150 460226
rect 79218 460170 79274 460226
rect 79342 460170 79398 460226
rect 78970 460046 79026 460102
rect 79094 460046 79150 460102
rect 79218 460046 79274 460102
rect 79342 460046 79398 460102
rect 78970 459922 79026 459978
rect 79094 459922 79150 459978
rect 79218 459922 79274 459978
rect 79342 459922 79398 459978
rect 93250 597156 93306 597212
rect 93374 597156 93430 597212
rect 93498 597156 93554 597212
rect 93622 597156 93678 597212
rect 93250 597032 93306 597088
rect 93374 597032 93430 597088
rect 93498 597032 93554 597088
rect 93622 597032 93678 597088
rect 93250 596908 93306 596964
rect 93374 596908 93430 596964
rect 93498 596908 93554 596964
rect 93622 596908 93678 596964
rect 93250 596784 93306 596840
rect 93374 596784 93430 596840
rect 93498 596784 93554 596840
rect 93622 596784 93678 596840
rect 93250 580294 93306 580350
rect 93374 580294 93430 580350
rect 93498 580294 93554 580350
rect 93622 580294 93678 580350
rect 93250 580170 93306 580226
rect 93374 580170 93430 580226
rect 93498 580170 93554 580226
rect 93622 580170 93678 580226
rect 93250 580046 93306 580102
rect 93374 580046 93430 580102
rect 93498 580046 93554 580102
rect 93622 580046 93678 580102
rect 93250 579922 93306 579978
rect 93374 579922 93430 579978
rect 93498 579922 93554 579978
rect 93622 579922 93678 579978
rect 93250 562294 93306 562350
rect 93374 562294 93430 562350
rect 93498 562294 93554 562350
rect 93622 562294 93678 562350
rect 93250 562170 93306 562226
rect 93374 562170 93430 562226
rect 93498 562170 93554 562226
rect 93622 562170 93678 562226
rect 93250 562046 93306 562102
rect 93374 562046 93430 562102
rect 93498 562046 93554 562102
rect 93622 562046 93678 562102
rect 93250 561922 93306 561978
rect 93374 561922 93430 561978
rect 93498 561922 93554 561978
rect 93622 561922 93678 561978
rect 93250 544294 93306 544350
rect 93374 544294 93430 544350
rect 93498 544294 93554 544350
rect 93622 544294 93678 544350
rect 93250 544170 93306 544226
rect 93374 544170 93430 544226
rect 93498 544170 93554 544226
rect 93622 544170 93678 544226
rect 93250 544046 93306 544102
rect 93374 544046 93430 544102
rect 93498 544046 93554 544102
rect 93622 544046 93678 544102
rect 93250 543922 93306 543978
rect 93374 543922 93430 543978
rect 93498 543922 93554 543978
rect 93622 543922 93678 543978
rect 93250 526294 93306 526350
rect 93374 526294 93430 526350
rect 93498 526294 93554 526350
rect 93622 526294 93678 526350
rect 93250 526170 93306 526226
rect 93374 526170 93430 526226
rect 93498 526170 93554 526226
rect 93622 526170 93678 526226
rect 93250 526046 93306 526102
rect 93374 526046 93430 526102
rect 93498 526046 93554 526102
rect 93622 526046 93678 526102
rect 93250 525922 93306 525978
rect 93374 525922 93430 525978
rect 93498 525922 93554 525978
rect 93622 525922 93678 525978
rect 93250 508294 93306 508350
rect 93374 508294 93430 508350
rect 93498 508294 93554 508350
rect 93622 508294 93678 508350
rect 93250 508170 93306 508226
rect 93374 508170 93430 508226
rect 93498 508170 93554 508226
rect 93622 508170 93678 508226
rect 93250 508046 93306 508102
rect 93374 508046 93430 508102
rect 93498 508046 93554 508102
rect 93622 508046 93678 508102
rect 93250 507922 93306 507978
rect 93374 507922 93430 507978
rect 93498 507922 93554 507978
rect 93622 507922 93678 507978
rect 93250 490294 93306 490350
rect 93374 490294 93430 490350
rect 93498 490294 93554 490350
rect 93622 490294 93678 490350
rect 93250 490170 93306 490226
rect 93374 490170 93430 490226
rect 93498 490170 93554 490226
rect 93622 490170 93678 490226
rect 93250 490046 93306 490102
rect 93374 490046 93430 490102
rect 93498 490046 93554 490102
rect 93622 490046 93678 490102
rect 93250 489922 93306 489978
rect 93374 489922 93430 489978
rect 93498 489922 93554 489978
rect 93622 489922 93678 489978
rect 93250 472294 93306 472350
rect 93374 472294 93430 472350
rect 93498 472294 93554 472350
rect 93622 472294 93678 472350
rect 93250 472170 93306 472226
rect 93374 472170 93430 472226
rect 93498 472170 93554 472226
rect 93622 472170 93678 472226
rect 93250 472046 93306 472102
rect 93374 472046 93430 472102
rect 93498 472046 93554 472102
rect 93622 472046 93678 472102
rect 93250 471922 93306 471978
rect 93374 471922 93430 471978
rect 93498 471922 93554 471978
rect 93622 471922 93678 471978
rect 96970 598116 97026 598172
rect 97094 598116 97150 598172
rect 97218 598116 97274 598172
rect 97342 598116 97398 598172
rect 96970 597992 97026 598048
rect 97094 597992 97150 598048
rect 97218 597992 97274 598048
rect 97342 597992 97398 598048
rect 96970 597868 97026 597924
rect 97094 597868 97150 597924
rect 97218 597868 97274 597924
rect 97342 597868 97398 597924
rect 96970 597744 97026 597800
rect 97094 597744 97150 597800
rect 97218 597744 97274 597800
rect 97342 597744 97398 597800
rect 96970 586294 97026 586350
rect 97094 586294 97150 586350
rect 97218 586294 97274 586350
rect 97342 586294 97398 586350
rect 96970 586170 97026 586226
rect 97094 586170 97150 586226
rect 97218 586170 97274 586226
rect 97342 586170 97398 586226
rect 96970 586046 97026 586102
rect 97094 586046 97150 586102
rect 97218 586046 97274 586102
rect 97342 586046 97398 586102
rect 96970 585922 97026 585978
rect 97094 585922 97150 585978
rect 97218 585922 97274 585978
rect 97342 585922 97398 585978
rect 96970 568294 97026 568350
rect 97094 568294 97150 568350
rect 97218 568294 97274 568350
rect 97342 568294 97398 568350
rect 96970 568170 97026 568226
rect 97094 568170 97150 568226
rect 97218 568170 97274 568226
rect 97342 568170 97398 568226
rect 96970 568046 97026 568102
rect 97094 568046 97150 568102
rect 97218 568046 97274 568102
rect 97342 568046 97398 568102
rect 96970 567922 97026 567978
rect 97094 567922 97150 567978
rect 97218 567922 97274 567978
rect 97342 567922 97398 567978
rect 96970 550294 97026 550350
rect 97094 550294 97150 550350
rect 97218 550294 97274 550350
rect 97342 550294 97398 550350
rect 96970 550170 97026 550226
rect 97094 550170 97150 550226
rect 97218 550170 97274 550226
rect 97342 550170 97398 550226
rect 96970 550046 97026 550102
rect 97094 550046 97150 550102
rect 97218 550046 97274 550102
rect 97342 550046 97398 550102
rect 96970 549922 97026 549978
rect 97094 549922 97150 549978
rect 97218 549922 97274 549978
rect 97342 549922 97398 549978
rect 96970 532294 97026 532350
rect 97094 532294 97150 532350
rect 97218 532294 97274 532350
rect 97342 532294 97398 532350
rect 96970 532170 97026 532226
rect 97094 532170 97150 532226
rect 97218 532170 97274 532226
rect 97342 532170 97398 532226
rect 96970 532046 97026 532102
rect 97094 532046 97150 532102
rect 97218 532046 97274 532102
rect 97342 532046 97398 532102
rect 96970 531922 97026 531978
rect 97094 531922 97150 531978
rect 97218 531922 97274 531978
rect 97342 531922 97398 531978
rect 96970 514294 97026 514350
rect 97094 514294 97150 514350
rect 97218 514294 97274 514350
rect 97342 514294 97398 514350
rect 96970 514170 97026 514226
rect 97094 514170 97150 514226
rect 97218 514170 97274 514226
rect 97342 514170 97398 514226
rect 96970 514046 97026 514102
rect 97094 514046 97150 514102
rect 97218 514046 97274 514102
rect 97342 514046 97398 514102
rect 96970 513922 97026 513978
rect 97094 513922 97150 513978
rect 97218 513922 97274 513978
rect 97342 513922 97398 513978
rect 96970 496294 97026 496350
rect 97094 496294 97150 496350
rect 97218 496294 97274 496350
rect 97342 496294 97398 496350
rect 96970 496170 97026 496226
rect 97094 496170 97150 496226
rect 97218 496170 97274 496226
rect 97342 496170 97398 496226
rect 96970 496046 97026 496102
rect 97094 496046 97150 496102
rect 97218 496046 97274 496102
rect 97342 496046 97398 496102
rect 96970 495922 97026 495978
rect 97094 495922 97150 495978
rect 97218 495922 97274 495978
rect 97342 495922 97398 495978
rect 96970 478294 97026 478350
rect 97094 478294 97150 478350
rect 97218 478294 97274 478350
rect 97342 478294 97398 478350
rect 96970 478170 97026 478226
rect 97094 478170 97150 478226
rect 97218 478170 97274 478226
rect 97342 478170 97398 478226
rect 96970 478046 97026 478102
rect 97094 478046 97150 478102
rect 97218 478046 97274 478102
rect 97342 478046 97398 478102
rect 96970 477922 97026 477978
rect 97094 477922 97150 477978
rect 97218 477922 97274 477978
rect 97342 477922 97398 477978
rect 96970 460294 97026 460350
rect 97094 460294 97150 460350
rect 97218 460294 97274 460350
rect 97342 460294 97398 460350
rect 96970 460170 97026 460226
rect 97094 460170 97150 460226
rect 97218 460170 97274 460226
rect 97342 460170 97398 460226
rect 96970 460046 97026 460102
rect 97094 460046 97150 460102
rect 97218 460046 97274 460102
rect 97342 460046 97398 460102
rect 96970 459922 97026 459978
rect 97094 459922 97150 459978
rect 97218 459922 97274 459978
rect 97342 459922 97398 459978
rect 111250 597156 111306 597212
rect 111374 597156 111430 597212
rect 111498 597156 111554 597212
rect 111622 597156 111678 597212
rect 111250 597032 111306 597088
rect 111374 597032 111430 597088
rect 111498 597032 111554 597088
rect 111622 597032 111678 597088
rect 111250 596908 111306 596964
rect 111374 596908 111430 596964
rect 111498 596908 111554 596964
rect 111622 596908 111678 596964
rect 111250 596784 111306 596840
rect 111374 596784 111430 596840
rect 111498 596784 111554 596840
rect 111622 596784 111678 596840
rect 111250 580294 111306 580350
rect 111374 580294 111430 580350
rect 111498 580294 111554 580350
rect 111622 580294 111678 580350
rect 111250 580170 111306 580226
rect 111374 580170 111430 580226
rect 111498 580170 111554 580226
rect 111622 580170 111678 580226
rect 111250 580046 111306 580102
rect 111374 580046 111430 580102
rect 111498 580046 111554 580102
rect 111622 580046 111678 580102
rect 111250 579922 111306 579978
rect 111374 579922 111430 579978
rect 111498 579922 111554 579978
rect 111622 579922 111678 579978
rect 111250 562294 111306 562350
rect 111374 562294 111430 562350
rect 111498 562294 111554 562350
rect 111622 562294 111678 562350
rect 111250 562170 111306 562226
rect 111374 562170 111430 562226
rect 111498 562170 111554 562226
rect 111622 562170 111678 562226
rect 111250 562046 111306 562102
rect 111374 562046 111430 562102
rect 111498 562046 111554 562102
rect 111622 562046 111678 562102
rect 111250 561922 111306 561978
rect 111374 561922 111430 561978
rect 111498 561922 111554 561978
rect 111622 561922 111678 561978
rect 111250 544294 111306 544350
rect 111374 544294 111430 544350
rect 111498 544294 111554 544350
rect 111622 544294 111678 544350
rect 111250 544170 111306 544226
rect 111374 544170 111430 544226
rect 111498 544170 111554 544226
rect 111622 544170 111678 544226
rect 111250 544046 111306 544102
rect 111374 544046 111430 544102
rect 111498 544046 111554 544102
rect 111622 544046 111678 544102
rect 111250 543922 111306 543978
rect 111374 543922 111430 543978
rect 111498 543922 111554 543978
rect 111622 543922 111678 543978
rect 111250 526294 111306 526350
rect 111374 526294 111430 526350
rect 111498 526294 111554 526350
rect 111622 526294 111678 526350
rect 111250 526170 111306 526226
rect 111374 526170 111430 526226
rect 111498 526170 111554 526226
rect 111622 526170 111678 526226
rect 111250 526046 111306 526102
rect 111374 526046 111430 526102
rect 111498 526046 111554 526102
rect 111622 526046 111678 526102
rect 111250 525922 111306 525978
rect 111374 525922 111430 525978
rect 111498 525922 111554 525978
rect 111622 525922 111678 525978
rect 111250 508294 111306 508350
rect 111374 508294 111430 508350
rect 111498 508294 111554 508350
rect 111622 508294 111678 508350
rect 111250 508170 111306 508226
rect 111374 508170 111430 508226
rect 111498 508170 111554 508226
rect 111622 508170 111678 508226
rect 111250 508046 111306 508102
rect 111374 508046 111430 508102
rect 111498 508046 111554 508102
rect 111622 508046 111678 508102
rect 111250 507922 111306 507978
rect 111374 507922 111430 507978
rect 111498 507922 111554 507978
rect 111622 507922 111678 507978
rect 111250 490294 111306 490350
rect 111374 490294 111430 490350
rect 111498 490294 111554 490350
rect 111622 490294 111678 490350
rect 111250 490170 111306 490226
rect 111374 490170 111430 490226
rect 111498 490170 111554 490226
rect 111622 490170 111678 490226
rect 111250 490046 111306 490102
rect 111374 490046 111430 490102
rect 111498 490046 111554 490102
rect 111622 490046 111678 490102
rect 111250 489922 111306 489978
rect 111374 489922 111430 489978
rect 111498 489922 111554 489978
rect 111622 489922 111678 489978
rect 111250 472294 111306 472350
rect 111374 472294 111430 472350
rect 111498 472294 111554 472350
rect 111622 472294 111678 472350
rect 111250 472170 111306 472226
rect 111374 472170 111430 472226
rect 111498 472170 111554 472226
rect 111622 472170 111678 472226
rect 111250 472046 111306 472102
rect 111374 472046 111430 472102
rect 111498 472046 111554 472102
rect 111622 472046 111678 472102
rect 111250 471922 111306 471978
rect 111374 471922 111430 471978
rect 111498 471922 111554 471978
rect 111622 471922 111678 471978
rect 114970 598116 115026 598172
rect 115094 598116 115150 598172
rect 115218 598116 115274 598172
rect 115342 598116 115398 598172
rect 114970 597992 115026 598048
rect 115094 597992 115150 598048
rect 115218 597992 115274 598048
rect 115342 597992 115398 598048
rect 114970 597868 115026 597924
rect 115094 597868 115150 597924
rect 115218 597868 115274 597924
rect 115342 597868 115398 597924
rect 114970 597744 115026 597800
rect 115094 597744 115150 597800
rect 115218 597744 115274 597800
rect 115342 597744 115398 597800
rect 114970 586294 115026 586350
rect 115094 586294 115150 586350
rect 115218 586294 115274 586350
rect 115342 586294 115398 586350
rect 114970 586170 115026 586226
rect 115094 586170 115150 586226
rect 115218 586170 115274 586226
rect 115342 586170 115398 586226
rect 114970 586046 115026 586102
rect 115094 586046 115150 586102
rect 115218 586046 115274 586102
rect 115342 586046 115398 586102
rect 114970 585922 115026 585978
rect 115094 585922 115150 585978
rect 115218 585922 115274 585978
rect 115342 585922 115398 585978
rect 114970 568294 115026 568350
rect 115094 568294 115150 568350
rect 115218 568294 115274 568350
rect 115342 568294 115398 568350
rect 114970 568170 115026 568226
rect 115094 568170 115150 568226
rect 115218 568170 115274 568226
rect 115342 568170 115398 568226
rect 114970 568046 115026 568102
rect 115094 568046 115150 568102
rect 115218 568046 115274 568102
rect 115342 568046 115398 568102
rect 114970 567922 115026 567978
rect 115094 567922 115150 567978
rect 115218 567922 115274 567978
rect 115342 567922 115398 567978
rect 114970 550294 115026 550350
rect 115094 550294 115150 550350
rect 115218 550294 115274 550350
rect 115342 550294 115398 550350
rect 114970 550170 115026 550226
rect 115094 550170 115150 550226
rect 115218 550170 115274 550226
rect 115342 550170 115398 550226
rect 114970 550046 115026 550102
rect 115094 550046 115150 550102
rect 115218 550046 115274 550102
rect 115342 550046 115398 550102
rect 114970 549922 115026 549978
rect 115094 549922 115150 549978
rect 115218 549922 115274 549978
rect 115342 549922 115398 549978
rect 114970 532294 115026 532350
rect 115094 532294 115150 532350
rect 115218 532294 115274 532350
rect 115342 532294 115398 532350
rect 114970 532170 115026 532226
rect 115094 532170 115150 532226
rect 115218 532170 115274 532226
rect 115342 532170 115398 532226
rect 114970 532046 115026 532102
rect 115094 532046 115150 532102
rect 115218 532046 115274 532102
rect 115342 532046 115398 532102
rect 114970 531922 115026 531978
rect 115094 531922 115150 531978
rect 115218 531922 115274 531978
rect 115342 531922 115398 531978
rect 114970 514294 115026 514350
rect 115094 514294 115150 514350
rect 115218 514294 115274 514350
rect 115342 514294 115398 514350
rect 114970 514170 115026 514226
rect 115094 514170 115150 514226
rect 115218 514170 115274 514226
rect 115342 514170 115398 514226
rect 114970 514046 115026 514102
rect 115094 514046 115150 514102
rect 115218 514046 115274 514102
rect 115342 514046 115398 514102
rect 114970 513922 115026 513978
rect 115094 513922 115150 513978
rect 115218 513922 115274 513978
rect 115342 513922 115398 513978
rect 114970 496294 115026 496350
rect 115094 496294 115150 496350
rect 115218 496294 115274 496350
rect 115342 496294 115398 496350
rect 114970 496170 115026 496226
rect 115094 496170 115150 496226
rect 115218 496170 115274 496226
rect 115342 496170 115398 496226
rect 114970 496046 115026 496102
rect 115094 496046 115150 496102
rect 115218 496046 115274 496102
rect 115342 496046 115398 496102
rect 114970 495922 115026 495978
rect 115094 495922 115150 495978
rect 115218 495922 115274 495978
rect 115342 495922 115398 495978
rect 114970 478294 115026 478350
rect 115094 478294 115150 478350
rect 115218 478294 115274 478350
rect 115342 478294 115398 478350
rect 114970 478170 115026 478226
rect 115094 478170 115150 478226
rect 115218 478170 115274 478226
rect 115342 478170 115398 478226
rect 114970 478046 115026 478102
rect 115094 478046 115150 478102
rect 115218 478046 115274 478102
rect 115342 478046 115398 478102
rect 114970 477922 115026 477978
rect 115094 477922 115150 477978
rect 115218 477922 115274 477978
rect 115342 477922 115398 477978
rect 114970 460294 115026 460350
rect 115094 460294 115150 460350
rect 115218 460294 115274 460350
rect 115342 460294 115398 460350
rect 114970 460170 115026 460226
rect 115094 460170 115150 460226
rect 115218 460170 115274 460226
rect 115342 460170 115398 460226
rect 114970 460046 115026 460102
rect 115094 460046 115150 460102
rect 115218 460046 115274 460102
rect 115342 460046 115398 460102
rect 114970 459922 115026 459978
rect 115094 459922 115150 459978
rect 115218 459922 115274 459978
rect 115342 459922 115398 459978
rect 129250 597156 129306 597212
rect 129374 597156 129430 597212
rect 129498 597156 129554 597212
rect 129622 597156 129678 597212
rect 129250 597032 129306 597088
rect 129374 597032 129430 597088
rect 129498 597032 129554 597088
rect 129622 597032 129678 597088
rect 129250 596908 129306 596964
rect 129374 596908 129430 596964
rect 129498 596908 129554 596964
rect 129622 596908 129678 596964
rect 129250 596784 129306 596840
rect 129374 596784 129430 596840
rect 129498 596784 129554 596840
rect 129622 596784 129678 596840
rect 129250 580294 129306 580350
rect 129374 580294 129430 580350
rect 129498 580294 129554 580350
rect 129622 580294 129678 580350
rect 129250 580170 129306 580226
rect 129374 580170 129430 580226
rect 129498 580170 129554 580226
rect 129622 580170 129678 580226
rect 129250 580046 129306 580102
rect 129374 580046 129430 580102
rect 129498 580046 129554 580102
rect 129622 580046 129678 580102
rect 129250 579922 129306 579978
rect 129374 579922 129430 579978
rect 129498 579922 129554 579978
rect 129622 579922 129678 579978
rect 129250 562294 129306 562350
rect 129374 562294 129430 562350
rect 129498 562294 129554 562350
rect 129622 562294 129678 562350
rect 129250 562170 129306 562226
rect 129374 562170 129430 562226
rect 129498 562170 129554 562226
rect 129622 562170 129678 562226
rect 129250 562046 129306 562102
rect 129374 562046 129430 562102
rect 129498 562046 129554 562102
rect 129622 562046 129678 562102
rect 129250 561922 129306 561978
rect 129374 561922 129430 561978
rect 129498 561922 129554 561978
rect 129622 561922 129678 561978
rect 129250 544294 129306 544350
rect 129374 544294 129430 544350
rect 129498 544294 129554 544350
rect 129622 544294 129678 544350
rect 129250 544170 129306 544226
rect 129374 544170 129430 544226
rect 129498 544170 129554 544226
rect 129622 544170 129678 544226
rect 129250 544046 129306 544102
rect 129374 544046 129430 544102
rect 129498 544046 129554 544102
rect 129622 544046 129678 544102
rect 129250 543922 129306 543978
rect 129374 543922 129430 543978
rect 129498 543922 129554 543978
rect 129622 543922 129678 543978
rect 129250 526294 129306 526350
rect 129374 526294 129430 526350
rect 129498 526294 129554 526350
rect 129622 526294 129678 526350
rect 129250 526170 129306 526226
rect 129374 526170 129430 526226
rect 129498 526170 129554 526226
rect 129622 526170 129678 526226
rect 129250 526046 129306 526102
rect 129374 526046 129430 526102
rect 129498 526046 129554 526102
rect 129622 526046 129678 526102
rect 129250 525922 129306 525978
rect 129374 525922 129430 525978
rect 129498 525922 129554 525978
rect 129622 525922 129678 525978
rect 129250 508294 129306 508350
rect 129374 508294 129430 508350
rect 129498 508294 129554 508350
rect 129622 508294 129678 508350
rect 129250 508170 129306 508226
rect 129374 508170 129430 508226
rect 129498 508170 129554 508226
rect 129622 508170 129678 508226
rect 129250 508046 129306 508102
rect 129374 508046 129430 508102
rect 129498 508046 129554 508102
rect 129622 508046 129678 508102
rect 129250 507922 129306 507978
rect 129374 507922 129430 507978
rect 129498 507922 129554 507978
rect 129622 507922 129678 507978
rect 129250 490294 129306 490350
rect 129374 490294 129430 490350
rect 129498 490294 129554 490350
rect 129622 490294 129678 490350
rect 129250 490170 129306 490226
rect 129374 490170 129430 490226
rect 129498 490170 129554 490226
rect 129622 490170 129678 490226
rect 129250 490046 129306 490102
rect 129374 490046 129430 490102
rect 129498 490046 129554 490102
rect 129622 490046 129678 490102
rect 129250 489922 129306 489978
rect 129374 489922 129430 489978
rect 129498 489922 129554 489978
rect 129622 489922 129678 489978
rect 129250 472294 129306 472350
rect 129374 472294 129430 472350
rect 129498 472294 129554 472350
rect 129622 472294 129678 472350
rect 129250 472170 129306 472226
rect 129374 472170 129430 472226
rect 129498 472170 129554 472226
rect 129622 472170 129678 472226
rect 129250 472046 129306 472102
rect 129374 472046 129430 472102
rect 129498 472046 129554 472102
rect 129622 472046 129678 472102
rect 129250 471922 129306 471978
rect 129374 471922 129430 471978
rect 129498 471922 129554 471978
rect 129622 471922 129678 471978
rect 132970 598116 133026 598172
rect 133094 598116 133150 598172
rect 133218 598116 133274 598172
rect 133342 598116 133398 598172
rect 132970 597992 133026 598048
rect 133094 597992 133150 598048
rect 133218 597992 133274 598048
rect 133342 597992 133398 598048
rect 132970 597868 133026 597924
rect 133094 597868 133150 597924
rect 133218 597868 133274 597924
rect 133342 597868 133398 597924
rect 132970 597744 133026 597800
rect 133094 597744 133150 597800
rect 133218 597744 133274 597800
rect 133342 597744 133398 597800
rect 132970 586294 133026 586350
rect 133094 586294 133150 586350
rect 133218 586294 133274 586350
rect 133342 586294 133398 586350
rect 132970 586170 133026 586226
rect 133094 586170 133150 586226
rect 133218 586170 133274 586226
rect 133342 586170 133398 586226
rect 132970 586046 133026 586102
rect 133094 586046 133150 586102
rect 133218 586046 133274 586102
rect 133342 586046 133398 586102
rect 132970 585922 133026 585978
rect 133094 585922 133150 585978
rect 133218 585922 133274 585978
rect 133342 585922 133398 585978
rect 132970 568294 133026 568350
rect 133094 568294 133150 568350
rect 133218 568294 133274 568350
rect 133342 568294 133398 568350
rect 132970 568170 133026 568226
rect 133094 568170 133150 568226
rect 133218 568170 133274 568226
rect 133342 568170 133398 568226
rect 132970 568046 133026 568102
rect 133094 568046 133150 568102
rect 133218 568046 133274 568102
rect 133342 568046 133398 568102
rect 132970 567922 133026 567978
rect 133094 567922 133150 567978
rect 133218 567922 133274 567978
rect 133342 567922 133398 567978
rect 132970 550294 133026 550350
rect 133094 550294 133150 550350
rect 133218 550294 133274 550350
rect 133342 550294 133398 550350
rect 132970 550170 133026 550226
rect 133094 550170 133150 550226
rect 133218 550170 133274 550226
rect 133342 550170 133398 550226
rect 132970 550046 133026 550102
rect 133094 550046 133150 550102
rect 133218 550046 133274 550102
rect 133342 550046 133398 550102
rect 132970 549922 133026 549978
rect 133094 549922 133150 549978
rect 133218 549922 133274 549978
rect 133342 549922 133398 549978
rect 132970 532294 133026 532350
rect 133094 532294 133150 532350
rect 133218 532294 133274 532350
rect 133342 532294 133398 532350
rect 132970 532170 133026 532226
rect 133094 532170 133150 532226
rect 133218 532170 133274 532226
rect 133342 532170 133398 532226
rect 132970 532046 133026 532102
rect 133094 532046 133150 532102
rect 133218 532046 133274 532102
rect 133342 532046 133398 532102
rect 132970 531922 133026 531978
rect 133094 531922 133150 531978
rect 133218 531922 133274 531978
rect 133342 531922 133398 531978
rect 132970 514294 133026 514350
rect 133094 514294 133150 514350
rect 133218 514294 133274 514350
rect 133342 514294 133398 514350
rect 132970 514170 133026 514226
rect 133094 514170 133150 514226
rect 133218 514170 133274 514226
rect 133342 514170 133398 514226
rect 132970 514046 133026 514102
rect 133094 514046 133150 514102
rect 133218 514046 133274 514102
rect 133342 514046 133398 514102
rect 132970 513922 133026 513978
rect 133094 513922 133150 513978
rect 133218 513922 133274 513978
rect 133342 513922 133398 513978
rect 132970 496294 133026 496350
rect 133094 496294 133150 496350
rect 133218 496294 133274 496350
rect 133342 496294 133398 496350
rect 132970 496170 133026 496226
rect 133094 496170 133150 496226
rect 133218 496170 133274 496226
rect 133342 496170 133398 496226
rect 132970 496046 133026 496102
rect 133094 496046 133150 496102
rect 133218 496046 133274 496102
rect 133342 496046 133398 496102
rect 132970 495922 133026 495978
rect 133094 495922 133150 495978
rect 133218 495922 133274 495978
rect 133342 495922 133398 495978
rect 132970 478294 133026 478350
rect 133094 478294 133150 478350
rect 133218 478294 133274 478350
rect 133342 478294 133398 478350
rect 132970 478170 133026 478226
rect 133094 478170 133150 478226
rect 133218 478170 133274 478226
rect 133342 478170 133398 478226
rect 132970 478046 133026 478102
rect 133094 478046 133150 478102
rect 133218 478046 133274 478102
rect 133342 478046 133398 478102
rect 132970 477922 133026 477978
rect 133094 477922 133150 477978
rect 133218 477922 133274 477978
rect 133342 477922 133398 477978
rect 132970 460294 133026 460350
rect 133094 460294 133150 460350
rect 133218 460294 133274 460350
rect 133342 460294 133398 460350
rect 132970 460170 133026 460226
rect 133094 460170 133150 460226
rect 133218 460170 133274 460226
rect 133342 460170 133398 460226
rect 132970 460046 133026 460102
rect 133094 460046 133150 460102
rect 133218 460046 133274 460102
rect 133342 460046 133398 460102
rect 132970 459922 133026 459978
rect 133094 459922 133150 459978
rect 133218 459922 133274 459978
rect 133342 459922 133398 459978
rect 147250 597156 147306 597212
rect 147374 597156 147430 597212
rect 147498 597156 147554 597212
rect 147622 597156 147678 597212
rect 147250 597032 147306 597088
rect 147374 597032 147430 597088
rect 147498 597032 147554 597088
rect 147622 597032 147678 597088
rect 147250 596908 147306 596964
rect 147374 596908 147430 596964
rect 147498 596908 147554 596964
rect 147622 596908 147678 596964
rect 147250 596784 147306 596840
rect 147374 596784 147430 596840
rect 147498 596784 147554 596840
rect 147622 596784 147678 596840
rect 147250 580294 147306 580350
rect 147374 580294 147430 580350
rect 147498 580294 147554 580350
rect 147622 580294 147678 580350
rect 147250 580170 147306 580226
rect 147374 580170 147430 580226
rect 147498 580170 147554 580226
rect 147622 580170 147678 580226
rect 147250 580046 147306 580102
rect 147374 580046 147430 580102
rect 147498 580046 147554 580102
rect 147622 580046 147678 580102
rect 147250 579922 147306 579978
rect 147374 579922 147430 579978
rect 147498 579922 147554 579978
rect 147622 579922 147678 579978
rect 147250 562294 147306 562350
rect 147374 562294 147430 562350
rect 147498 562294 147554 562350
rect 147622 562294 147678 562350
rect 147250 562170 147306 562226
rect 147374 562170 147430 562226
rect 147498 562170 147554 562226
rect 147622 562170 147678 562226
rect 147250 562046 147306 562102
rect 147374 562046 147430 562102
rect 147498 562046 147554 562102
rect 147622 562046 147678 562102
rect 147250 561922 147306 561978
rect 147374 561922 147430 561978
rect 147498 561922 147554 561978
rect 147622 561922 147678 561978
rect 147250 544294 147306 544350
rect 147374 544294 147430 544350
rect 147498 544294 147554 544350
rect 147622 544294 147678 544350
rect 147250 544170 147306 544226
rect 147374 544170 147430 544226
rect 147498 544170 147554 544226
rect 147622 544170 147678 544226
rect 147250 544046 147306 544102
rect 147374 544046 147430 544102
rect 147498 544046 147554 544102
rect 147622 544046 147678 544102
rect 147250 543922 147306 543978
rect 147374 543922 147430 543978
rect 147498 543922 147554 543978
rect 147622 543922 147678 543978
rect 147250 526294 147306 526350
rect 147374 526294 147430 526350
rect 147498 526294 147554 526350
rect 147622 526294 147678 526350
rect 147250 526170 147306 526226
rect 147374 526170 147430 526226
rect 147498 526170 147554 526226
rect 147622 526170 147678 526226
rect 147250 526046 147306 526102
rect 147374 526046 147430 526102
rect 147498 526046 147554 526102
rect 147622 526046 147678 526102
rect 147250 525922 147306 525978
rect 147374 525922 147430 525978
rect 147498 525922 147554 525978
rect 147622 525922 147678 525978
rect 147250 508294 147306 508350
rect 147374 508294 147430 508350
rect 147498 508294 147554 508350
rect 147622 508294 147678 508350
rect 147250 508170 147306 508226
rect 147374 508170 147430 508226
rect 147498 508170 147554 508226
rect 147622 508170 147678 508226
rect 147250 508046 147306 508102
rect 147374 508046 147430 508102
rect 147498 508046 147554 508102
rect 147622 508046 147678 508102
rect 147250 507922 147306 507978
rect 147374 507922 147430 507978
rect 147498 507922 147554 507978
rect 147622 507922 147678 507978
rect 147250 490294 147306 490350
rect 147374 490294 147430 490350
rect 147498 490294 147554 490350
rect 147622 490294 147678 490350
rect 147250 490170 147306 490226
rect 147374 490170 147430 490226
rect 147498 490170 147554 490226
rect 147622 490170 147678 490226
rect 147250 490046 147306 490102
rect 147374 490046 147430 490102
rect 147498 490046 147554 490102
rect 147622 490046 147678 490102
rect 147250 489922 147306 489978
rect 147374 489922 147430 489978
rect 147498 489922 147554 489978
rect 147622 489922 147678 489978
rect 147250 472294 147306 472350
rect 147374 472294 147430 472350
rect 147498 472294 147554 472350
rect 147622 472294 147678 472350
rect 147250 472170 147306 472226
rect 147374 472170 147430 472226
rect 147498 472170 147554 472226
rect 147622 472170 147678 472226
rect 147250 472046 147306 472102
rect 147374 472046 147430 472102
rect 147498 472046 147554 472102
rect 147622 472046 147678 472102
rect 147250 471922 147306 471978
rect 147374 471922 147430 471978
rect 147498 471922 147554 471978
rect 147622 471922 147678 471978
rect 150970 598116 151026 598172
rect 151094 598116 151150 598172
rect 151218 598116 151274 598172
rect 151342 598116 151398 598172
rect 150970 597992 151026 598048
rect 151094 597992 151150 598048
rect 151218 597992 151274 598048
rect 151342 597992 151398 598048
rect 150970 597868 151026 597924
rect 151094 597868 151150 597924
rect 151218 597868 151274 597924
rect 151342 597868 151398 597924
rect 150970 597744 151026 597800
rect 151094 597744 151150 597800
rect 151218 597744 151274 597800
rect 151342 597744 151398 597800
rect 150970 586294 151026 586350
rect 151094 586294 151150 586350
rect 151218 586294 151274 586350
rect 151342 586294 151398 586350
rect 150970 586170 151026 586226
rect 151094 586170 151150 586226
rect 151218 586170 151274 586226
rect 151342 586170 151398 586226
rect 150970 586046 151026 586102
rect 151094 586046 151150 586102
rect 151218 586046 151274 586102
rect 151342 586046 151398 586102
rect 150970 585922 151026 585978
rect 151094 585922 151150 585978
rect 151218 585922 151274 585978
rect 151342 585922 151398 585978
rect 150970 568294 151026 568350
rect 151094 568294 151150 568350
rect 151218 568294 151274 568350
rect 151342 568294 151398 568350
rect 150970 568170 151026 568226
rect 151094 568170 151150 568226
rect 151218 568170 151274 568226
rect 151342 568170 151398 568226
rect 150970 568046 151026 568102
rect 151094 568046 151150 568102
rect 151218 568046 151274 568102
rect 151342 568046 151398 568102
rect 150970 567922 151026 567978
rect 151094 567922 151150 567978
rect 151218 567922 151274 567978
rect 151342 567922 151398 567978
rect 150970 550294 151026 550350
rect 151094 550294 151150 550350
rect 151218 550294 151274 550350
rect 151342 550294 151398 550350
rect 150970 550170 151026 550226
rect 151094 550170 151150 550226
rect 151218 550170 151274 550226
rect 151342 550170 151398 550226
rect 150970 550046 151026 550102
rect 151094 550046 151150 550102
rect 151218 550046 151274 550102
rect 151342 550046 151398 550102
rect 150970 549922 151026 549978
rect 151094 549922 151150 549978
rect 151218 549922 151274 549978
rect 151342 549922 151398 549978
rect 150970 532294 151026 532350
rect 151094 532294 151150 532350
rect 151218 532294 151274 532350
rect 151342 532294 151398 532350
rect 150970 532170 151026 532226
rect 151094 532170 151150 532226
rect 151218 532170 151274 532226
rect 151342 532170 151398 532226
rect 150970 532046 151026 532102
rect 151094 532046 151150 532102
rect 151218 532046 151274 532102
rect 151342 532046 151398 532102
rect 150970 531922 151026 531978
rect 151094 531922 151150 531978
rect 151218 531922 151274 531978
rect 151342 531922 151398 531978
rect 150970 514294 151026 514350
rect 151094 514294 151150 514350
rect 151218 514294 151274 514350
rect 151342 514294 151398 514350
rect 150970 514170 151026 514226
rect 151094 514170 151150 514226
rect 151218 514170 151274 514226
rect 151342 514170 151398 514226
rect 150970 514046 151026 514102
rect 151094 514046 151150 514102
rect 151218 514046 151274 514102
rect 151342 514046 151398 514102
rect 150970 513922 151026 513978
rect 151094 513922 151150 513978
rect 151218 513922 151274 513978
rect 151342 513922 151398 513978
rect 150970 496294 151026 496350
rect 151094 496294 151150 496350
rect 151218 496294 151274 496350
rect 151342 496294 151398 496350
rect 150970 496170 151026 496226
rect 151094 496170 151150 496226
rect 151218 496170 151274 496226
rect 151342 496170 151398 496226
rect 150970 496046 151026 496102
rect 151094 496046 151150 496102
rect 151218 496046 151274 496102
rect 151342 496046 151398 496102
rect 150970 495922 151026 495978
rect 151094 495922 151150 495978
rect 151218 495922 151274 495978
rect 151342 495922 151398 495978
rect 150970 478294 151026 478350
rect 151094 478294 151150 478350
rect 151218 478294 151274 478350
rect 151342 478294 151398 478350
rect 150970 478170 151026 478226
rect 151094 478170 151150 478226
rect 151218 478170 151274 478226
rect 151342 478170 151398 478226
rect 150970 478046 151026 478102
rect 151094 478046 151150 478102
rect 151218 478046 151274 478102
rect 151342 478046 151398 478102
rect 150970 477922 151026 477978
rect 151094 477922 151150 477978
rect 151218 477922 151274 477978
rect 151342 477922 151398 477978
rect 150970 460294 151026 460350
rect 151094 460294 151150 460350
rect 151218 460294 151274 460350
rect 151342 460294 151398 460350
rect 150970 460170 151026 460226
rect 151094 460170 151150 460226
rect 151218 460170 151274 460226
rect 151342 460170 151398 460226
rect 150970 460046 151026 460102
rect 151094 460046 151150 460102
rect 151218 460046 151274 460102
rect 151342 460046 151398 460102
rect 150970 459922 151026 459978
rect 151094 459922 151150 459978
rect 151218 459922 151274 459978
rect 151342 459922 151398 459978
rect 165250 597156 165306 597212
rect 165374 597156 165430 597212
rect 165498 597156 165554 597212
rect 165622 597156 165678 597212
rect 165250 597032 165306 597088
rect 165374 597032 165430 597088
rect 165498 597032 165554 597088
rect 165622 597032 165678 597088
rect 165250 596908 165306 596964
rect 165374 596908 165430 596964
rect 165498 596908 165554 596964
rect 165622 596908 165678 596964
rect 165250 596784 165306 596840
rect 165374 596784 165430 596840
rect 165498 596784 165554 596840
rect 165622 596784 165678 596840
rect 165250 580294 165306 580350
rect 165374 580294 165430 580350
rect 165498 580294 165554 580350
rect 165622 580294 165678 580350
rect 165250 580170 165306 580226
rect 165374 580170 165430 580226
rect 165498 580170 165554 580226
rect 165622 580170 165678 580226
rect 165250 580046 165306 580102
rect 165374 580046 165430 580102
rect 165498 580046 165554 580102
rect 165622 580046 165678 580102
rect 165250 579922 165306 579978
rect 165374 579922 165430 579978
rect 165498 579922 165554 579978
rect 165622 579922 165678 579978
rect 165250 562294 165306 562350
rect 165374 562294 165430 562350
rect 165498 562294 165554 562350
rect 165622 562294 165678 562350
rect 165250 562170 165306 562226
rect 165374 562170 165430 562226
rect 165498 562170 165554 562226
rect 165622 562170 165678 562226
rect 165250 562046 165306 562102
rect 165374 562046 165430 562102
rect 165498 562046 165554 562102
rect 165622 562046 165678 562102
rect 165250 561922 165306 561978
rect 165374 561922 165430 561978
rect 165498 561922 165554 561978
rect 165622 561922 165678 561978
rect 165250 544294 165306 544350
rect 165374 544294 165430 544350
rect 165498 544294 165554 544350
rect 165622 544294 165678 544350
rect 165250 544170 165306 544226
rect 165374 544170 165430 544226
rect 165498 544170 165554 544226
rect 165622 544170 165678 544226
rect 165250 544046 165306 544102
rect 165374 544046 165430 544102
rect 165498 544046 165554 544102
rect 165622 544046 165678 544102
rect 165250 543922 165306 543978
rect 165374 543922 165430 543978
rect 165498 543922 165554 543978
rect 165622 543922 165678 543978
rect 165250 526294 165306 526350
rect 165374 526294 165430 526350
rect 165498 526294 165554 526350
rect 165622 526294 165678 526350
rect 165250 526170 165306 526226
rect 165374 526170 165430 526226
rect 165498 526170 165554 526226
rect 165622 526170 165678 526226
rect 165250 526046 165306 526102
rect 165374 526046 165430 526102
rect 165498 526046 165554 526102
rect 165622 526046 165678 526102
rect 165250 525922 165306 525978
rect 165374 525922 165430 525978
rect 165498 525922 165554 525978
rect 165622 525922 165678 525978
rect 165250 508294 165306 508350
rect 165374 508294 165430 508350
rect 165498 508294 165554 508350
rect 165622 508294 165678 508350
rect 165250 508170 165306 508226
rect 165374 508170 165430 508226
rect 165498 508170 165554 508226
rect 165622 508170 165678 508226
rect 165250 508046 165306 508102
rect 165374 508046 165430 508102
rect 165498 508046 165554 508102
rect 165622 508046 165678 508102
rect 165250 507922 165306 507978
rect 165374 507922 165430 507978
rect 165498 507922 165554 507978
rect 165622 507922 165678 507978
rect 165250 490294 165306 490350
rect 165374 490294 165430 490350
rect 165498 490294 165554 490350
rect 165622 490294 165678 490350
rect 165250 490170 165306 490226
rect 165374 490170 165430 490226
rect 165498 490170 165554 490226
rect 165622 490170 165678 490226
rect 165250 490046 165306 490102
rect 165374 490046 165430 490102
rect 165498 490046 165554 490102
rect 165622 490046 165678 490102
rect 165250 489922 165306 489978
rect 165374 489922 165430 489978
rect 165498 489922 165554 489978
rect 165622 489922 165678 489978
rect 165250 472294 165306 472350
rect 165374 472294 165430 472350
rect 165498 472294 165554 472350
rect 165622 472294 165678 472350
rect 165250 472170 165306 472226
rect 165374 472170 165430 472226
rect 165498 472170 165554 472226
rect 165622 472170 165678 472226
rect 165250 472046 165306 472102
rect 165374 472046 165430 472102
rect 165498 472046 165554 472102
rect 165622 472046 165678 472102
rect 165250 471922 165306 471978
rect 165374 471922 165430 471978
rect 165498 471922 165554 471978
rect 165622 471922 165678 471978
rect 168970 598116 169026 598172
rect 169094 598116 169150 598172
rect 169218 598116 169274 598172
rect 169342 598116 169398 598172
rect 168970 597992 169026 598048
rect 169094 597992 169150 598048
rect 169218 597992 169274 598048
rect 169342 597992 169398 598048
rect 168970 597868 169026 597924
rect 169094 597868 169150 597924
rect 169218 597868 169274 597924
rect 169342 597868 169398 597924
rect 168970 597744 169026 597800
rect 169094 597744 169150 597800
rect 169218 597744 169274 597800
rect 169342 597744 169398 597800
rect 168970 586294 169026 586350
rect 169094 586294 169150 586350
rect 169218 586294 169274 586350
rect 169342 586294 169398 586350
rect 168970 586170 169026 586226
rect 169094 586170 169150 586226
rect 169218 586170 169274 586226
rect 169342 586170 169398 586226
rect 168970 586046 169026 586102
rect 169094 586046 169150 586102
rect 169218 586046 169274 586102
rect 169342 586046 169398 586102
rect 168970 585922 169026 585978
rect 169094 585922 169150 585978
rect 169218 585922 169274 585978
rect 169342 585922 169398 585978
rect 168970 568294 169026 568350
rect 169094 568294 169150 568350
rect 169218 568294 169274 568350
rect 169342 568294 169398 568350
rect 168970 568170 169026 568226
rect 169094 568170 169150 568226
rect 169218 568170 169274 568226
rect 169342 568170 169398 568226
rect 168970 568046 169026 568102
rect 169094 568046 169150 568102
rect 169218 568046 169274 568102
rect 169342 568046 169398 568102
rect 168970 567922 169026 567978
rect 169094 567922 169150 567978
rect 169218 567922 169274 567978
rect 169342 567922 169398 567978
rect 168970 550294 169026 550350
rect 169094 550294 169150 550350
rect 169218 550294 169274 550350
rect 169342 550294 169398 550350
rect 168970 550170 169026 550226
rect 169094 550170 169150 550226
rect 169218 550170 169274 550226
rect 169342 550170 169398 550226
rect 168970 550046 169026 550102
rect 169094 550046 169150 550102
rect 169218 550046 169274 550102
rect 169342 550046 169398 550102
rect 168970 549922 169026 549978
rect 169094 549922 169150 549978
rect 169218 549922 169274 549978
rect 169342 549922 169398 549978
rect 168970 532294 169026 532350
rect 169094 532294 169150 532350
rect 169218 532294 169274 532350
rect 169342 532294 169398 532350
rect 168970 532170 169026 532226
rect 169094 532170 169150 532226
rect 169218 532170 169274 532226
rect 169342 532170 169398 532226
rect 168970 532046 169026 532102
rect 169094 532046 169150 532102
rect 169218 532046 169274 532102
rect 169342 532046 169398 532102
rect 168970 531922 169026 531978
rect 169094 531922 169150 531978
rect 169218 531922 169274 531978
rect 169342 531922 169398 531978
rect 168970 514294 169026 514350
rect 169094 514294 169150 514350
rect 169218 514294 169274 514350
rect 169342 514294 169398 514350
rect 168970 514170 169026 514226
rect 169094 514170 169150 514226
rect 169218 514170 169274 514226
rect 169342 514170 169398 514226
rect 168970 514046 169026 514102
rect 169094 514046 169150 514102
rect 169218 514046 169274 514102
rect 169342 514046 169398 514102
rect 168970 513922 169026 513978
rect 169094 513922 169150 513978
rect 169218 513922 169274 513978
rect 169342 513922 169398 513978
rect 168970 496294 169026 496350
rect 169094 496294 169150 496350
rect 169218 496294 169274 496350
rect 169342 496294 169398 496350
rect 168970 496170 169026 496226
rect 169094 496170 169150 496226
rect 169218 496170 169274 496226
rect 169342 496170 169398 496226
rect 168970 496046 169026 496102
rect 169094 496046 169150 496102
rect 169218 496046 169274 496102
rect 169342 496046 169398 496102
rect 168970 495922 169026 495978
rect 169094 495922 169150 495978
rect 169218 495922 169274 495978
rect 169342 495922 169398 495978
rect 168970 478294 169026 478350
rect 169094 478294 169150 478350
rect 169218 478294 169274 478350
rect 169342 478294 169398 478350
rect 168970 478170 169026 478226
rect 169094 478170 169150 478226
rect 169218 478170 169274 478226
rect 169342 478170 169398 478226
rect 168970 478046 169026 478102
rect 169094 478046 169150 478102
rect 169218 478046 169274 478102
rect 169342 478046 169398 478102
rect 168970 477922 169026 477978
rect 169094 477922 169150 477978
rect 169218 477922 169274 477978
rect 169342 477922 169398 477978
rect 168970 460294 169026 460350
rect 169094 460294 169150 460350
rect 169218 460294 169274 460350
rect 169342 460294 169398 460350
rect 168970 460170 169026 460226
rect 169094 460170 169150 460226
rect 169218 460170 169274 460226
rect 169342 460170 169398 460226
rect 168970 460046 169026 460102
rect 169094 460046 169150 460102
rect 169218 460046 169274 460102
rect 169342 460046 169398 460102
rect 168970 459922 169026 459978
rect 169094 459922 169150 459978
rect 169218 459922 169274 459978
rect 169342 459922 169398 459978
rect 183250 597156 183306 597212
rect 183374 597156 183430 597212
rect 183498 597156 183554 597212
rect 183622 597156 183678 597212
rect 183250 597032 183306 597088
rect 183374 597032 183430 597088
rect 183498 597032 183554 597088
rect 183622 597032 183678 597088
rect 183250 596908 183306 596964
rect 183374 596908 183430 596964
rect 183498 596908 183554 596964
rect 183622 596908 183678 596964
rect 183250 596784 183306 596840
rect 183374 596784 183430 596840
rect 183498 596784 183554 596840
rect 183622 596784 183678 596840
rect 183250 580294 183306 580350
rect 183374 580294 183430 580350
rect 183498 580294 183554 580350
rect 183622 580294 183678 580350
rect 183250 580170 183306 580226
rect 183374 580170 183430 580226
rect 183498 580170 183554 580226
rect 183622 580170 183678 580226
rect 183250 580046 183306 580102
rect 183374 580046 183430 580102
rect 183498 580046 183554 580102
rect 183622 580046 183678 580102
rect 183250 579922 183306 579978
rect 183374 579922 183430 579978
rect 183498 579922 183554 579978
rect 183622 579922 183678 579978
rect 183250 562294 183306 562350
rect 183374 562294 183430 562350
rect 183498 562294 183554 562350
rect 183622 562294 183678 562350
rect 183250 562170 183306 562226
rect 183374 562170 183430 562226
rect 183498 562170 183554 562226
rect 183622 562170 183678 562226
rect 183250 562046 183306 562102
rect 183374 562046 183430 562102
rect 183498 562046 183554 562102
rect 183622 562046 183678 562102
rect 183250 561922 183306 561978
rect 183374 561922 183430 561978
rect 183498 561922 183554 561978
rect 183622 561922 183678 561978
rect 183250 544294 183306 544350
rect 183374 544294 183430 544350
rect 183498 544294 183554 544350
rect 183622 544294 183678 544350
rect 183250 544170 183306 544226
rect 183374 544170 183430 544226
rect 183498 544170 183554 544226
rect 183622 544170 183678 544226
rect 183250 544046 183306 544102
rect 183374 544046 183430 544102
rect 183498 544046 183554 544102
rect 183622 544046 183678 544102
rect 183250 543922 183306 543978
rect 183374 543922 183430 543978
rect 183498 543922 183554 543978
rect 183622 543922 183678 543978
rect 183250 526294 183306 526350
rect 183374 526294 183430 526350
rect 183498 526294 183554 526350
rect 183622 526294 183678 526350
rect 183250 526170 183306 526226
rect 183374 526170 183430 526226
rect 183498 526170 183554 526226
rect 183622 526170 183678 526226
rect 183250 526046 183306 526102
rect 183374 526046 183430 526102
rect 183498 526046 183554 526102
rect 183622 526046 183678 526102
rect 183250 525922 183306 525978
rect 183374 525922 183430 525978
rect 183498 525922 183554 525978
rect 183622 525922 183678 525978
rect 183250 508294 183306 508350
rect 183374 508294 183430 508350
rect 183498 508294 183554 508350
rect 183622 508294 183678 508350
rect 183250 508170 183306 508226
rect 183374 508170 183430 508226
rect 183498 508170 183554 508226
rect 183622 508170 183678 508226
rect 183250 508046 183306 508102
rect 183374 508046 183430 508102
rect 183498 508046 183554 508102
rect 183622 508046 183678 508102
rect 183250 507922 183306 507978
rect 183374 507922 183430 507978
rect 183498 507922 183554 507978
rect 183622 507922 183678 507978
rect 183250 490294 183306 490350
rect 183374 490294 183430 490350
rect 183498 490294 183554 490350
rect 183622 490294 183678 490350
rect 183250 490170 183306 490226
rect 183374 490170 183430 490226
rect 183498 490170 183554 490226
rect 183622 490170 183678 490226
rect 183250 490046 183306 490102
rect 183374 490046 183430 490102
rect 183498 490046 183554 490102
rect 183622 490046 183678 490102
rect 183250 489922 183306 489978
rect 183374 489922 183430 489978
rect 183498 489922 183554 489978
rect 183622 489922 183678 489978
rect 183250 472294 183306 472350
rect 183374 472294 183430 472350
rect 183498 472294 183554 472350
rect 183622 472294 183678 472350
rect 183250 472170 183306 472226
rect 183374 472170 183430 472226
rect 183498 472170 183554 472226
rect 183622 472170 183678 472226
rect 183250 472046 183306 472102
rect 183374 472046 183430 472102
rect 183498 472046 183554 472102
rect 183622 472046 183678 472102
rect 183250 471922 183306 471978
rect 183374 471922 183430 471978
rect 183498 471922 183554 471978
rect 183622 471922 183678 471978
rect 186970 598116 187026 598172
rect 187094 598116 187150 598172
rect 187218 598116 187274 598172
rect 187342 598116 187398 598172
rect 186970 597992 187026 598048
rect 187094 597992 187150 598048
rect 187218 597992 187274 598048
rect 187342 597992 187398 598048
rect 186970 597868 187026 597924
rect 187094 597868 187150 597924
rect 187218 597868 187274 597924
rect 187342 597868 187398 597924
rect 186970 597744 187026 597800
rect 187094 597744 187150 597800
rect 187218 597744 187274 597800
rect 187342 597744 187398 597800
rect 201250 597156 201306 597212
rect 201374 597156 201430 597212
rect 201498 597156 201554 597212
rect 201622 597156 201678 597212
rect 201250 597032 201306 597088
rect 201374 597032 201430 597088
rect 201498 597032 201554 597088
rect 201622 597032 201678 597088
rect 201250 596908 201306 596964
rect 201374 596908 201430 596964
rect 201498 596908 201554 596964
rect 201622 596908 201678 596964
rect 201250 596784 201306 596840
rect 201374 596784 201430 596840
rect 201498 596784 201554 596840
rect 201622 596784 201678 596840
rect 186970 586294 187026 586350
rect 187094 586294 187150 586350
rect 187218 586294 187274 586350
rect 187342 586294 187398 586350
rect 186970 586170 187026 586226
rect 187094 586170 187150 586226
rect 187218 586170 187274 586226
rect 187342 586170 187398 586226
rect 186970 586046 187026 586102
rect 187094 586046 187150 586102
rect 187218 586046 187274 586102
rect 187342 586046 187398 586102
rect 186970 585922 187026 585978
rect 187094 585922 187150 585978
rect 187218 585922 187274 585978
rect 187342 585922 187398 585978
rect 186970 568294 187026 568350
rect 187094 568294 187150 568350
rect 187218 568294 187274 568350
rect 187342 568294 187398 568350
rect 186970 568170 187026 568226
rect 187094 568170 187150 568226
rect 187218 568170 187274 568226
rect 187342 568170 187398 568226
rect 186970 568046 187026 568102
rect 187094 568046 187150 568102
rect 187218 568046 187274 568102
rect 187342 568046 187398 568102
rect 186970 567922 187026 567978
rect 187094 567922 187150 567978
rect 187218 567922 187274 567978
rect 187342 567922 187398 567978
rect 186970 550294 187026 550350
rect 187094 550294 187150 550350
rect 187218 550294 187274 550350
rect 187342 550294 187398 550350
rect 186970 550170 187026 550226
rect 187094 550170 187150 550226
rect 187218 550170 187274 550226
rect 187342 550170 187398 550226
rect 186970 550046 187026 550102
rect 187094 550046 187150 550102
rect 187218 550046 187274 550102
rect 187342 550046 187398 550102
rect 186970 549922 187026 549978
rect 187094 549922 187150 549978
rect 187218 549922 187274 549978
rect 187342 549922 187398 549978
rect 186970 532294 187026 532350
rect 187094 532294 187150 532350
rect 187218 532294 187274 532350
rect 187342 532294 187398 532350
rect 186970 532170 187026 532226
rect 187094 532170 187150 532226
rect 187218 532170 187274 532226
rect 187342 532170 187398 532226
rect 186970 532046 187026 532102
rect 187094 532046 187150 532102
rect 187218 532046 187274 532102
rect 187342 532046 187398 532102
rect 186970 531922 187026 531978
rect 187094 531922 187150 531978
rect 187218 531922 187274 531978
rect 187342 531922 187398 531978
rect 186970 514294 187026 514350
rect 187094 514294 187150 514350
rect 187218 514294 187274 514350
rect 187342 514294 187398 514350
rect 186970 514170 187026 514226
rect 187094 514170 187150 514226
rect 187218 514170 187274 514226
rect 187342 514170 187398 514226
rect 186970 514046 187026 514102
rect 187094 514046 187150 514102
rect 187218 514046 187274 514102
rect 187342 514046 187398 514102
rect 186970 513922 187026 513978
rect 187094 513922 187150 513978
rect 187218 513922 187274 513978
rect 187342 513922 187398 513978
rect 186970 496294 187026 496350
rect 187094 496294 187150 496350
rect 187218 496294 187274 496350
rect 187342 496294 187398 496350
rect 186970 496170 187026 496226
rect 187094 496170 187150 496226
rect 187218 496170 187274 496226
rect 187342 496170 187398 496226
rect 186970 496046 187026 496102
rect 187094 496046 187150 496102
rect 187218 496046 187274 496102
rect 187342 496046 187398 496102
rect 186970 495922 187026 495978
rect 187094 495922 187150 495978
rect 187218 495922 187274 495978
rect 187342 495922 187398 495978
rect 186970 478294 187026 478350
rect 187094 478294 187150 478350
rect 187218 478294 187274 478350
rect 187342 478294 187398 478350
rect 186970 478170 187026 478226
rect 187094 478170 187150 478226
rect 187218 478170 187274 478226
rect 187342 478170 187398 478226
rect 186970 478046 187026 478102
rect 187094 478046 187150 478102
rect 187218 478046 187274 478102
rect 187342 478046 187398 478102
rect 186970 477922 187026 477978
rect 187094 477922 187150 477978
rect 187218 477922 187274 477978
rect 187342 477922 187398 477978
rect 186970 460294 187026 460350
rect 187094 460294 187150 460350
rect 187218 460294 187274 460350
rect 187342 460294 187398 460350
rect 186970 460170 187026 460226
rect 187094 460170 187150 460226
rect 187218 460170 187274 460226
rect 187342 460170 187398 460226
rect 186970 460046 187026 460102
rect 187094 460046 187150 460102
rect 187218 460046 187274 460102
rect 187342 460046 187398 460102
rect 186970 459922 187026 459978
rect 187094 459922 187150 459978
rect 187218 459922 187274 459978
rect 187342 459922 187398 459978
rect 24970 316294 25026 316350
rect 25094 316294 25150 316350
rect 25218 316294 25274 316350
rect 25342 316294 25398 316350
rect 24970 316170 25026 316226
rect 25094 316170 25150 316226
rect 25218 316170 25274 316226
rect 25342 316170 25398 316226
rect 24970 316046 25026 316102
rect 25094 316046 25150 316102
rect 25218 316046 25274 316102
rect 25342 316046 25398 316102
rect 24970 315922 25026 315978
rect 25094 315922 25150 315978
rect 25218 315922 25274 315978
rect 25342 315922 25398 315978
rect 24970 298366 25026 298422
rect 25094 298366 25150 298422
rect 25218 298366 25274 298422
rect 25342 298366 25398 298422
rect 42970 316294 43026 316350
rect 43094 316294 43150 316350
rect 43218 316294 43274 316350
rect 43342 316294 43398 316350
rect 42970 316170 43026 316226
rect 43094 316170 43150 316226
rect 43218 316170 43274 316226
rect 43342 316170 43398 316226
rect 42970 316046 43026 316102
rect 43094 316046 43150 316102
rect 43218 316046 43274 316102
rect 43342 316046 43398 316102
rect 42970 315922 43026 315978
rect 43094 315922 43150 315978
rect 43218 315922 43274 315978
rect 43342 315922 43398 315978
rect 42970 298366 43026 298422
rect 43094 298366 43150 298422
rect 43218 298366 43274 298422
rect 43342 298366 43398 298422
rect 60970 316294 61026 316350
rect 61094 316294 61150 316350
rect 61218 316294 61274 316350
rect 61342 316294 61398 316350
rect 60970 316170 61026 316226
rect 61094 316170 61150 316226
rect 61218 316170 61274 316226
rect 61342 316170 61398 316226
rect 60970 316046 61026 316102
rect 61094 316046 61150 316102
rect 61218 316046 61274 316102
rect 61342 316046 61398 316102
rect 60970 315922 61026 315978
rect 61094 315922 61150 315978
rect 61218 315922 61274 315978
rect 61342 315922 61398 315978
rect 60970 298366 61026 298422
rect 61094 298366 61150 298422
rect 61218 298366 61274 298422
rect 61342 298366 61398 298422
rect 78970 316294 79026 316350
rect 79094 316294 79150 316350
rect 79218 316294 79274 316350
rect 79342 316294 79398 316350
rect 78970 316170 79026 316226
rect 79094 316170 79150 316226
rect 79218 316170 79274 316226
rect 79342 316170 79398 316226
rect 78970 316046 79026 316102
rect 79094 316046 79150 316102
rect 79218 316046 79274 316102
rect 79342 316046 79398 316102
rect 78970 315922 79026 315978
rect 79094 315922 79150 315978
rect 79218 315922 79274 315978
rect 79342 315922 79398 315978
rect 78970 298366 79026 298422
rect 79094 298366 79150 298422
rect 79218 298366 79274 298422
rect 79342 298366 79398 298422
rect 96970 316294 97026 316350
rect 97094 316294 97150 316350
rect 97218 316294 97274 316350
rect 97342 316294 97398 316350
rect 96970 316170 97026 316226
rect 97094 316170 97150 316226
rect 97218 316170 97274 316226
rect 97342 316170 97398 316226
rect 96970 316046 97026 316102
rect 97094 316046 97150 316102
rect 97218 316046 97274 316102
rect 97342 316046 97398 316102
rect 96970 315922 97026 315978
rect 97094 315922 97150 315978
rect 97218 315922 97274 315978
rect 97342 315922 97398 315978
rect 96970 298366 97026 298422
rect 97094 298366 97150 298422
rect 97218 298366 97274 298422
rect 97342 298366 97398 298422
rect 114970 316294 115026 316350
rect 115094 316294 115150 316350
rect 115218 316294 115274 316350
rect 115342 316294 115398 316350
rect 114970 316170 115026 316226
rect 115094 316170 115150 316226
rect 115218 316170 115274 316226
rect 115342 316170 115398 316226
rect 114970 316046 115026 316102
rect 115094 316046 115150 316102
rect 115218 316046 115274 316102
rect 115342 316046 115398 316102
rect 114970 315922 115026 315978
rect 115094 315922 115150 315978
rect 115218 315922 115274 315978
rect 115342 315922 115398 315978
rect 114970 298366 115026 298422
rect 115094 298366 115150 298422
rect 115218 298366 115274 298422
rect 115342 298366 115398 298422
rect 132970 316294 133026 316350
rect 133094 316294 133150 316350
rect 133218 316294 133274 316350
rect 133342 316294 133398 316350
rect 132970 316170 133026 316226
rect 133094 316170 133150 316226
rect 133218 316170 133274 316226
rect 133342 316170 133398 316226
rect 132970 316046 133026 316102
rect 133094 316046 133150 316102
rect 133218 316046 133274 316102
rect 133342 316046 133398 316102
rect 132970 315922 133026 315978
rect 133094 315922 133150 315978
rect 133218 315922 133274 315978
rect 133342 315922 133398 315978
rect 132970 298366 133026 298422
rect 133094 298366 133150 298422
rect 133218 298366 133274 298422
rect 133342 298366 133398 298422
rect 150970 316294 151026 316350
rect 151094 316294 151150 316350
rect 151218 316294 151274 316350
rect 151342 316294 151398 316350
rect 150970 316170 151026 316226
rect 151094 316170 151150 316226
rect 151218 316170 151274 316226
rect 151342 316170 151398 316226
rect 150970 316046 151026 316102
rect 151094 316046 151150 316102
rect 151218 316046 151274 316102
rect 151342 316046 151398 316102
rect 150970 315922 151026 315978
rect 151094 315922 151150 315978
rect 151218 315922 151274 315978
rect 151342 315922 151398 315978
rect 150970 298366 151026 298422
rect 151094 298366 151150 298422
rect 151218 298366 151274 298422
rect 151342 298366 151398 298422
rect 168970 316294 169026 316350
rect 169094 316294 169150 316350
rect 169218 316294 169274 316350
rect 169342 316294 169398 316350
rect 168970 316170 169026 316226
rect 169094 316170 169150 316226
rect 169218 316170 169274 316226
rect 169342 316170 169398 316226
rect 168970 316046 169026 316102
rect 169094 316046 169150 316102
rect 169218 316046 169274 316102
rect 169342 316046 169398 316102
rect 168970 315922 169026 315978
rect 169094 315922 169150 315978
rect 169218 315922 169274 315978
rect 169342 315922 169398 315978
rect 168970 298366 169026 298422
rect 169094 298366 169150 298422
rect 169218 298366 169274 298422
rect 169342 298366 169398 298422
rect 186970 316294 187026 316350
rect 187094 316294 187150 316350
rect 187218 316294 187274 316350
rect 187342 316294 187398 316350
rect 186970 316170 187026 316226
rect 187094 316170 187150 316226
rect 187218 316170 187274 316226
rect 187342 316170 187398 316226
rect 186970 316046 187026 316102
rect 187094 316046 187150 316102
rect 187218 316046 187274 316102
rect 187342 316046 187398 316102
rect 186970 315922 187026 315978
rect 187094 315922 187150 315978
rect 187218 315922 187274 315978
rect 187342 315922 187398 315978
rect 186970 298366 187026 298422
rect 187094 298366 187150 298422
rect 187218 298366 187274 298422
rect 187342 298366 187398 298422
rect 21250 148294 21306 148350
rect 21374 148294 21430 148350
rect 21498 148294 21554 148350
rect 21622 148294 21678 148350
rect 21250 148170 21306 148226
rect 21374 148170 21430 148226
rect 21498 148170 21554 148226
rect 21622 148170 21678 148226
rect 21250 148046 21306 148102
rect 21374 148046 21430 148102
rect 21498 148046 21554 148102
rect 21622 148046 21678 148102
rect 21250 147922 21306 147978
rect 21374 147922 21430 147978
rect 21498 147922 21554 147978
rect 21622 147922 21678 147978
rect 21250 130294 21306 130350
rect 21374 130294 21430 130350
rect 21498 130294 21554 130350
rect 21622 130294 21678 130350
rect 21250 130170 21306 130226
rect 21374 130170 21430 130226
rect 21498 130170 21554 130226
rect 21622 130170 21678 130226
rect 21250 130046 21306 130102
rect 21374 130046 21430 130102
rect 21498 130046 21554 130102
rect 21622 130046 21678 130102
rect 21250 129922 21306 129978
rect 21374 129922 21430 129978
rect 21498 129922 21554 129978
rect 21622 129922 21678 129978
rect 6970 10294 7026 10350
rect 7094 10294 7150 10350
rect 7218 10294 7274 10350
rect 7342 10294 7398 10350
rect 6970 10170 7026 10226
rect 7094 10170 7150 10226
rect 7218 10170 7274 10226
rect 7342 10170 7398 10226
rect 6970 10046 7026 10102
rect 7094 10046 7150 10102
rect 7218 10046 7274 10102
rect 7342 10046 7398 10102
rect 21250 112294 21306 112350
rect 21374 112294 21430 112350
rect 21498 112294 21554 112350
rect 21622 112294 21678 112350
rect 21250 112170 21306 112226
rect 21374 112170 21430 112226
rect 21498 112170 21554 112226
rect 21622 112170 21678 112226
rect 21250 112046 21306 112102
rect 21374 112046 21430 112102
rect 21498 112046 21554 112102
rect 21622 112046 21678 112102
rect 21250 111922 21306 111978
rect 21374 111922 21430 111978
rect 21498 111922 21554 111978
rect 21622 111922 21678 111978
rect 21250 94294 21306 94350
rect 21374 94294 21430 94350
rect 21498 94294 21554 94350
rect 21622 94294 21678 94350
rect 21250 94170 21306 94226
rect 21374 94170 21430 94226
rect 21498 94170 21554 94226
rect 21622 94170 21678 94226
rect 21250 94046 21306 94102
rect 21374 94046 21430 94102
rect 21498 94046 21554 94102
rect 21622 94046 21678 94102
rect 21250 93922 21306 93978
rect 21374 93922 21430 93978
rect 21498 93922 21554 93978
rect 21622 93922 21678 93978
rect 24970 154294 25026 154350
rect 25094 154294 25150 154350
rect 25218 154294 25274 154350
rect 25342 154294 25398 154350
rect 24970 154170 25026 154226
rect 25094 154170 25150 154226
rect 25218 154170 25274 154226
rect 25342 154170 25398 154226
rect 24970 154046 25026 154102
rect 25094 154046 25150 154102
rect 25218 154046 25274 154102
rect 25342 154046 25398 154102
rect 24970 153922 25026 153978
rect 25094 153922 25150 153978
rect 25218 153922 25274 153978
rect 25342 153922 25398 153978
rect 24970 136294 25026 136350
rect 25094 136294 25150 136350
rect 25218 136294 25274 136350
rect 25342 136294 25398 136350
rect 24970 136170 25026 136226
rect 25094 136170 25150 136226
rect 25218 136170 25274 136226
rect 25342 136170 25398 136226
rect 24970 136046 25026 136102
rect 25094 136046 25150 136102
rect 25218 136046 25274 136102
rect 25342 136046 25398 136102
rect 24970 135922 25026 135978
rect 25094 135922 25150 135978
rect 25218 135922 25274 135978
rect 25342 135922 25398 135978
rect 24970 118294 25026 118350
rect 25094 118294 25150 118350
rect 25218 118294 25274 118350
rect 25342 118294 25398 118350
rect 24970 118170 25026 118226
rect 25094 118170 25150 118226
rect 25218 118170 25274 118226
rect 25342 118170 25398 118226
rect 24970 118046 25026 118102
rect 25094 118046 25150 118102
rect 25218 118046 25274 118102
rect 25342 118046 25398 118102
rect 24970 117922 25026 117978
rect 25094 117922 25150 117978
rect 25218 117922 25274 117978
rect 25342 117922 25398 117978
rect 24970 100294 25026 100350
rect 25094 100294 25150 100350
rect 25218 100294 25274 100350
rect 25342 100294 25398 100350
rect 24970 100170 25026 100226
rect 25094 100170 25150 100226
rect 25218 100170 25274 100226
rect 25342 100170 25398 100226
rect 24970 100046 25026 100102
rect 25094 100046 25150 100102
rect 25218 100046 25274 100102
rect 25342 100046 25398 100102
rect 24970 99922 25026 99978
rect 25094 99922 25150 99978
rect 25218 99922 25274 99978
rect 25342 99922 25398 99978
rect 24970 82294 25026 82350
rect 25094 82294 25150 82350
rect 25218 82294 25274 82350
rect 25342 82294 25398 82350
rect 21250 76294 21306 76350
rect 21374 76294 21430 76350
rect 21498 76294 21554 76350
rect 21622 76294 21678 76350
rect 21250 76170 21306 76226
rect 21374 76170 21430 76226
rect 21498 76170 21554 76226
rect 21622 76170 21678 76226
rect 21250 76046 21306 76102
rect 21374 76046 21430 76102
rect 21498 76046 21554 76102
rect 21622 76046 21678 76102
rect 21250 75922 21306 75978
rect 21374 75922 21430 75978
rect 21498 75922 21554 75978
rect 21622 75922 21678 75978
rect 21250 58294 21306 58350
rect 21374 58294 21430 58350
rect 21498 58294 21554 58350
rect 21622 58294 21678 58350
rect 21250 58170 21306 58226
rect 21374 58170 21430 58226
rect 21498 58170 21554 58226
rect 21622 58170 21678 58226
rect 21250 58046 21306 58102
rect 21374 58046 21430 58102
rect 21498 58046 21554 58102
rect 21622 58046 21678 58102
rect 21250 57922 21306 57978
rect 21374 57922 21430 57978
rect 21498 57922 21554 57978
rect 21622 57922 21678 57978
rect 21250 40294 21306 40350
rect 21374 40294 21430 40350
rect 21498 40294 21554 40350
rect 21622 40294 21678 40350
rect 21250 40170 21306 40226
rect 21374 40170 21430 40226
rect 21498 40170 21554 40226
rect 21622 40170 21678 40226
rect 21250 40046 21306 40102
rect 21374 40046 21430 40102
rect 21498 40046 21554 40102
rect 21622 40046 21678 40102
rect 21250 39922 21306 39978
rect 21374 39922 21430 39978
rect 21498 39922 21554 39978
rect 21622 39922 21678 39978
rect 21250 22294 21306 22350
rect 21374 22294 21430 22350
rect 21498 22294 21554 22350
rect 21622 22294 21678 22350
rect 21250 22170 21306 22226
rect 21374 22170 21430 22226
rect 21498 22170 21554 22226
rect 21622 22170 21678 22226
rect 21250 22046 21306 22102
rect 21374 22046 21430 22102
rect 21498 22046 21554 22102
rect 21622 22046 21678 22102
rect 21250 21922 21306 21978
rect 21374 21922 21430 21978
rect 21498 21922 21554 21978
rect 21622 21922 21678 21978
rect 6970 9922 7026 9978
rect 7094 9922 7150 9978
rect 7218 9922 7274 9978
rect 7342 9922 7398 9978
rect 6970 -1176 7026 -1120
rect 7094 -1176 7150 -1120
rect 7218 -1176 7274 -1120
rect 7342 -1176 7398 -1120
rect 6970 -1300 7026 -1244
rect 7094 -1300 7150 -1244
rect 7218 -1300 7274 -1244
rect 7342 -1300 7398 -1244
rect 6970 -1424 7026 -1368
rect 7094 -1424 7150 -1368
rect 7218 -1424 7274 -1368
rect 7342 -1424 7398 -1368
rect 6970 -1548 7026 -1492
rect 7094 -1548 7150 -1492
rect 7218 -1548 7274 -1492
rect 7342 -1548 7398 -1492
rect 24970 82170 25026 82226
rect 25094 82170 25150 82226
rect 25218 82170 25274 82226
rect 25342 82170 25398 82226
rect 24970 82046 25026 82102
rect 25094 82046 25150 82102
rect 25218 82046 25274 82102
rect 25342 82046 25398 82102
rect 24970 81922 25026 81978
rect 25094 81922 25150 81978
rect 25218 81922 25274 81978
rect 25342 81922 25398 81978
rect 39250 148294 39306 148350
rect 39374 148294 39430 148350
rect 39498 148294 39554 148350
rect 39622 148294 39678 148350
rect 39250 148170 39306 148226
rect 39374 148170 39430 148226
rect 39498 148170 39554 148226
rect 39622 148170 39678 148226
rect 39250 148046 39306 148102
rect 39374 148046 39430 148102
rect 39498 148046 39554 148102
rect 39622 148046 39678 148102
rect 39250 147922 39306 147978
rect 39374 147922 39430 147978
rect 39498 147922 39554 147978
rect 39622 147922 39678 147978
rect 39250 130294 39306 130350
rect 39374 130294 39430 130350
rect 39498 130294 39554 130350
rect 39622 130294 39678 130350
rect 39250 130170 39306 130226
rect 39374 130170 39430 130226
rect 39498 130170 39554 130226
rect 39622 130170 39678 130226
rect 39250 130046 39306 130102
rect 39374 130046 39430 130102
rect 39498 130046 39554 130102
rect 39622 130046 39678 130102
rect 39250 129922 39306 129978
rect 39374 129922 39430 129978
rect 39498 129922 39554 129978
rect 39622 129922 39678 129978
rect 39250 112294 39306 112350
rect 39374 112294 39430 112350
rect 39498 112294 39554 112350
rect 39622 112294 39678 112350
rect 39250 112170 39306 112226
rect 39374 112170 39430 112226
rect 39498 112170 39554 112226
rect 39622 112170 39678 112226
rect 39250 112046 39306 112102
rect 39374 112046 39430 112102
rect 39498 112046 39554 112102
rect 39622 112046 39678 112102
rect 39250 111922 39306 111978
rect 39374 111922 39430 111978
rect 39498 111922 39554 111978
rect 39622 111922 39678 111978
rect 39250 94294 39306 94350
rect 39374 94294 39430 94350
rect 39498 94294 39554 94350
rect 39622 94294 39678 94350
rect 39250 94170 39306 94226
rect 39374 94170 39430 94226
rect 39498 94170 39554 94226
rect 39622 94170 39678 94226
rect 39250 94046 39306 94102
rect 39374 94046 39430 94102
rect 39498 94046 39554 94102
rect 39622 94046 39678 94102
rect 39250 93922 39306 93978
rect 39374 93922 39430 93978
rect 39498 93922 39554 93978
rect 39622 93922 39678 93978
rect 39250 76294 39306 76350
rect 39374 76294 39430 76350
rect 39498 76294 39554 76350
rect 39622 76294 39678 76350
rect 39250 76170 39306 76226
rect 39374 76170 39430 76226
rect 39498 76170 39554 76226
rect 39622 76170 39678 76226
rect 39250 76046 39306 76102
rect 39374 76046 39430 76102
rect 39498 76046 39554 76102
rect 39622 76046 39678 76102
rect 39250 75922 39306 75978
rect 39374 75922 39430 75978
rect 39498 75922 39554 75978
rect 39622 75922 39678 75978
rect 24970 64294 25026 64350
rect 25094 64294 25150 64350
rect 25218 64294 25274 64350
rect 25342 64294 25398 64350
rect 24970 64170 25026 64226
rect 25094 64170 25150 64226
rect 25218 64170 25274 64226
rect 25342 64170 25398 64226
rect 24970 64046 25026 64102
rect 25094 64046 25150 64102
rect 25218 64046 25274 64102
rect 25342 64046 25398 64102
rect 24970 63922 25026 63978
rect 25094 63922 25150 63978
rect 25218 63922 25274 63978
rect 25342 63922 25398 63978
rect 24970 46294 25026 46350
rect 25094 46294 25150 46350
rect 25218 46294 25274 46350
rect 25342 46294 25398 46350
rect 24970 46170 25026 46226
rect 25094 46170 25150 46226
rect 25218 46170 25274 46226
rect 25342 46170 25398 46226
rect 24970 46046 25026 46102
rect 25094 46046 25150 46102
rect 25218 46046 25274 46102
rect 25342 46046 25398 46102
rect 24970 45922 25026 45978
rect 25094 45922 25150 45978
rect 25218 45922 25274 45978
rect 25342 45922 25398 45978
rect 24970 28294 25026 28350
rect 25094 28294 25150 28350
rect 25218 28294 25274 28350
rect 25342 28294 25398 28350
rect 24970 28170 25026 28226
rect 25094 28170 25150 28226
rect 25218 28170 25274 28226
rect 25342 28170 25398 28226
rect 24970 28046 25026 28102
rect 25094 28046 25150 28102
rect 25218 28046 25274 28102
rect 25342 28046 25398 28102
rect 24970 27922 25026 27978
rect 25094 27922 25150 27978
rect 25218 27922 25274 27978
rect 25342 27922 25398 27978
rect 21250 4294 21306 4350
rect 21374 4294 21430 4350
rect 21498 4294 21554 4350
rect 21622 4294 21678 4350
rect 21250 4170 21306 4226
rect 21374 4170 21430 4226
rect 21498 4170 21554 4226
rect 21622 4170 21678 4226
rect 21250 4046 21306 4102
rect 21374 4046 21430 4102
rect 21498 4046 21554 4102
rect 21622 4046 21678 4102
rect 21250 3922 21306 3978
rect 21374 3922 21430 3978
rect 21498 3922 21554 3978
rect 21622 3922 21678 3978
rect 21250 -216 21306 -160
rect 21374 -216 21430 -160
rect 21498 -216 21554 -160
rect 21622 -216 21678 -160
rect 21250 -340 21306 -284
rect 21374 -340 21430 -284
rect 21498 -340 21554 -284
rect 21622 -340 21678 -284
rect 21250 -464 21306 -408
rect 21374 -464 21430 -408
rect 21498 -464 21554 -408
rect 21622 -464 21678 -408
rect 21250 -588 21306 -532
rect 21374 -588 21430 -532
rect 21498 -588 21554 -532
rect 21622 -588 21678 -532
rect 24970 10294 25026 10350
rect 25094 10294 25150 10350
rect 25218 10294 25274 10350
rect 25342 10294 25398 10350
rect 24970 10170 25026 10226
rect 25094 10170 25150 10226
rect 25218 10170 25274 10226
rect 25342 10170 25398 10226
rect 24970 10046 25026 10102
rect 25094 10046 25150 10102
rect 25218 10046 25274 10102
rect 25342 10046 25398 10102
rect 24970 9922 25026 9978
rect 25094 9922 25150 9978
rect 25218 9922 25274 9978
rect 25342 9922 25398 9978
rect 42970 154294 43026 154350
rect 43094 154294 43150 154350
rect 43218 154294 43274 154350
rect 43342 154294 43398 154350
rect 42970 154170 43026 154226
rect 43094 154170 43150 154226
rect 43218 154170 43274 154226
rect 43342 154170 43398 154226
rect 42970 154046 43026 154102
rect 43094 154046 43150 154102
rect 43218 154046 43274 154102
rect 43342 154046 43398 154102
rect 42970 153922 43026 153978
rect 43094 153922 43150 153978
rect 43218 153922 43274 153978
rect 43342 153922 43398 153978
rect 42970 136294 43026 136350
rect 43094 136294 43150 136350
rect 43218 136294 43274 136350
rect 43342 136294 43398 136350
rect 42970 136170 43026 136226
rect 43094 136170 43150 136226
rect 43218 136170 43274 136226
rect 43342 136170 43398 136226
rect 42970 136046 43026 136102
rect 43094 136046 43150 136102
rect 43218 136046 43274 136102
rect 43342 136046 43398 136102
rect 42970 135922 43026 135978
rect 43094 135922 43150 135978
rect 43218 135922 43274 135978
rect 43342 135922 43398 135978
rect 42970 118294 43026 118350
rect 43094 118294 43150 118350
rect 43218 118294 43274 118350
rect 43342 118294 43398 118350
rect 42970 118170 43026 118226
rect 43094 118170 43150 118226
rect 43218 118170 43274 118226
rect 43342 118170 43398 118226
rect 42970 118046 43026 118102
rect 43094 118046 43150 118102
rect 43218 118046 43274 118102
rect 43342 118046 43398 118102
rect 42970 117922 43026 117978
rect 43094 117922 43150 117978
rect 43218 117922 43274 117978
rect 43342 117922 43398 117978
rect 57250 148294 57306 148350
rect 57374 148294 57430 148350
rect 57498 148294 57554 148350
rect 57622 148294 57678 148350
rect 57250 148170 57306 148226
rect 57374 148170 57430 148226
rect 57498 148170 57554 148226
rect 57622 148170 57678 148226
rect 57250 148046 57306 148102
rect 57374 148046 57430 148102
rect 57498 148046 57554 148102
rect 57622 148046 57678 148102
rect 57250 147922 57306 147978
rect 57374 147922 57430 147978
rect 57498 147922 57554 147978
rect 57622 147922 57678 147978
rect 57250 130294 57306 130350
rect 57374 130294 57430 130350
rect 57498 130294 57554 130350
rect 57622 130294 57678 130350
rect 57250 130170 57306 130226
rect 57374 130170 57430 130226
rect 57498 130170 57554 130226
rect 57622 130170 57678 130226
rect 57250 130046 57306 130102
rect 57374 130046 57430 130102
rect 57498 130046 57554 130102
rect 57622 130046 57678 130102
rect 57250 129922 57306 129978
rect 57374 129922 57430 129978
rect 57498 129922 57554 129978
rect 57622 129922 57678 129978
rect 57250 112294 57306 112350
rect 57374 112294 57430 112350
rect 57498 112294 57554 112350
rect 57622 112294 57678 112350
rect 57250 112170 57306 112226
rect 57374 112170 57430 112226
rect 57498 112170 57554 112226
rect 57622 112170 57678 112226
rect 57250 112046 57306 112102
rect 57374 112046 57430 112102
rect 57498 112046 57554 112102
rect 57622 112046 57678 112102
rect 57250 111922 57306 111978
rect 57374 111922 57430 111978
rect 57498 111922 57554 111978
rect 57622 111922 57678 111978
rect 60970 154294 61026 154350
rect 61094 154294 61150 154350
rect 61218 154294 61274 154350
rect 61342 154294 61398 154350
rect 60970 154170 61026 154226
rect 61094 154170 61150 154226
rect 61218 154170 61274 154226
rect 61342 154170 61398 154226
rect 60970 154046 61026 154102
rect 61094 154046 61150 154102
rect 61218 154046 61274 154102
rect 61342 154046 61398 154102
rect 60970 153922 61026 153978
rect 61094 153922 61150 153978
rect 61218 153922 61274 153978
rect 61342 153922 61398 153978
rect 60970 136294 61026 136350
rect 61094 136294 61150 136350
rect 61218 136294 61274 136350
rect 61342 136294 61398 136350
rect 60970 136170 61026 136226
rect 61094 136170 61150 136226
rect 61218 136170 61274 136226
rect 61342 136170 61398 136226
rect 60970 136046 61026 136102
rect 61094 136046 61150 136102
rect 61218 136046 61274 136102
rect 61342 136046 61398 136102
rect 60970 135922 61026 135978
rect 61094 135922 61150 135978
rect 61218 135922 61274 135978
rect 61342 135922 61398 135978
rect 60970 118294 61026 118350
rect 61094 118294 61150 118350
rect 61218 118294 61274 118350
rect 61342 118294 61398 118350
rect 60970 118170 61026 118226
rect 61094 118170 61150 118226
rect 61218 118170 61274 118226
rect 61342 118170 61398 118226
rect 60970 118046 61026 118102
rect 61094 118046 61150 118102
rect 61218 118046 61274 118102
rect 61342 118046 61398 118102
rect 60970 117922 61026 117978
rect 61094 117922 61150 117978
rect 61218 117922 61274 117978
rect 61342 117922 61398 117978
rect 75250 148294 75306 148350
rect 75374 148294 75430 148350
rect 75498 148294 75554 148350
rect 75622 148294 75678 148350
rect 75250 148170 75306 148226
rect 75374 148170 75430 148226
rect 75498 148170 75554 148226
rect 75622 148170 75678 148226
rect 75250 148046 75306 148102
rect 75374 148046 75430 148102
rect 75498 148046 75554 148102
rect 75622 148046 75678 148102
rect 75250 147922 75306 147978
rect 75374 147922 75430 147978
rect 75498 147922 75554 147978
rect 75622 147922 75678 147978
rect 75250 130294 75306 130350
rect 75374 130294 75430 130350
rect 75498 130294 75554 130350
rect 75622 130294 75678 130350
rect 75250 130170 75306 130226
rect 75374 130170 75430 130226
rect 75498 130170 75554 130226
rect 75622 130170 75678 130226
rect 75250 130046 75306 130102
rect 75374 130046 75430 130102
rect 75498 130046 75554 130102
rect 75622 130046 75678 130102
rect 75250 129922 75306 129978
rect 75374 129922 75430 129978
rect 75498 129922 75554 129978
rect 75622 129922 75678 129978
rect 75250 112294 75306 112350
rect 75374 112294 75430 112350
rect 75498 112294 75554 112350
rect 75622 112294 75678 112350
rect 75250 112170 75306 112226
rect 75374 112170 75430 112226
rect 75498 112170 75554 112226
rect 75622 112170 75678 112226
rect 75250 112046 75306 112102
rect 75374 112046 75430 112102
rect 75498 112046 75554 112102
rect 75622 112046 75678 112102
rect 75250 111922 75306 111978
rect 75374 111922 75430 111978
rect 75498 111922 75554 111978
rect 75622 111922 75678 111978
rect 78970 154294 79026 154350
rect 79094 154294 79150 154350
rect 79218 154294 79274 154350
rect 79342 154294 79398 154350
rect 78970 154170 79026 154226
rect 79094 154170 79150 154226
rect 79218 154170 79274 154226
rect 79342 154170 79398 154226
rect 78970 154046 79026 154102
rect 79094 154046 79150 154102
rect 79218 154046 79274 154102
rect 79342 154046 79398 154102
rect 78970 153922 79026 153978
rect 79094 153922 79150 153978
rect 79218 153922 79274 153978
rect 79342 153922 79398 153978
rect 78970 136294 79026 136350
rect 79094 136294 79150 136350
rect 79218 136294 79274 136350
rect 79342 136294 79398 136350
rect 78970 136170 79026 136226
rect 79094 136170 79150 136226
rect 79218 136170 79274 136226
rect 79342 136170 79398 136226
rect 78970 136046 79026 136102
rect 79094 136046 79150 136102
rect 79218 136046 79274 136102
rect 79342 136046 79398 136102
rect 78970 135922 79026 135978
rect 79094 135922 79150 135978
rect 79218 135922 79274 135978
rect 79342 135922 79398 135978
rect 78970 118294 79026 118350
rect 79094 118294 79150 118350
rect 79218 118294 79274 118350
rect 79342 118294 79398 118350
rect 78970 118170 79026 118226
rect 79094 118170 79150 118226
rect 79218 118170 79274 118226
rect 79342 118170 79398 118226
rect 78970 118046 79026 118102
rect 79094 118046 79150 118102
rect 79218 118046 79274 118102
rect 79342 118046 79398 118102
rect 78970 117922 79026 117978
rect 79094 117922 79150 117978
rect 79218 117922 79274 117978
rect 79342 117922 79398 117978
rect 93250 148294 93306 148350
rect 93374 148294 93430 148350
rect 93498 148294 93554 148350
rect 93622 148294 93678 148350
rect 93250 148170 93306 148226
rect 93374 148170 93430 148226
rect 93498 148170 93554 148226
rect 93622 148170 93678 148226
rect 93250 148046 93306 148102
rect 93374 148046 93430 148102
rect 93498 148046 93554 148102
rect 93622 148046 93678 148102
rect 93250 147922 93306 147978
rect 93374 147922 93430 147978
rect 93498 147922 93554 147978
rect 93622 147922 93678 147978
rect 93250 130294 93306 130350
rect 93374 130294 93430 130350
rect 93498 130294 93554 130350
rect 93622 130294 93678 130350
rect 93250 130170 93306 130226
rect 93374 130170 93430 130226
rect 93498 130170 93554 130226
rect 93622 130170 93678 130226
rect 93250 130046 93306 130102
rect 93374 130046 93430 130102
rect 93498 130046 93554 130102
rect 93622 130046 93678 130102
rect 93250 129922 93306 129978
rect 93374 129922 93430 129978
rect 93498 129922 93554 129978
rect 93622 129922 93678 129978
rect 93250 112294 93306 112350
rect 93374 112294 93430 112350
rect 93498 112294 93554 112350
rect 93622 112294 93678 112350
rect 93250 112170 93306 112226
rect 93374 112170 93430 112226
rect 93498 112170 93554 112226
rect 93622 112170 93678 112226
rect 93250 112046 93306 112102
rect 93374 112046 93430 112102
rect 93498 112046 93554 112102
rect 93622 112046 93678 112102
rect 93250 111922 93306 111978
rect 93374 111922 93430 111978
rect 93498 111922 93554 111978
rect 93622 111922 93678 111978
rect 96970 154294 97026 154350
rect 97094 154294 97150 154350
rect 97218 154294 97274 154350
rect 97342 154294 97398 154350
rect 96970 154170 97026 154226
rect 97094 154170 97150 154226
rect 97218 154170 97274 154226
rect 97342 154170 97398 154226
rect 96970 154046 97026 154102
rect 97094 154046 97150 154102
rect 97218 154046 97274 154102
rect 97342 154046 97398 154102
rect 96970 153922 97026 153978
rect 97094 153922 97150 153978
rect 97218 153922 97274 153978
rect 97342 153922 97398 153978
rect 96970 136294 97026 136350
rect 97094 136294 97150 136350
rect 97218 136294 97274 136350
rect 97342 136294 97398 136350
rect 96970 136170 97026 136226
rect 97094 136170 97150 136226
rect 97218 136170 97274 136226
rect 97342 136170 97398 136226
rect 96970 136046 97026 136102
rect 97094 136046 97150 136102
rect 97218 136046 97274 136102
rect 97342 136046 97398 136102
rect 96970 135922 97026 135978
rect 97094 135922 97150 135978
rect 97218 135922 97274 135978
rect 97342 135922 97398 135978
rect 96970 118294 97026 118350
rect 97094 118294 97150 118350
rect 97218 118294 97274 118350
rect 97342 118294 97398 118350
rect 96970 118170 97026 118226
rect 97094 118170 97150 118226
rect 97218 118170 97274 118226
rect 97342 118170 97398 118226
rect 96970 118046 97026 118102
rect 97094 118046 97150 118102
rect 97218 118046 97274 118102
rect 97342 118046 97398 118102
rect 96970 117922 97026 117978
rect 97094 117922 97150 117978
rect 97218 117922 97274 117978
rect 97342 117922 97398 117978
rect 111250 148294 111306 148350
rect 111374 148294 111430 148350
rect 111498 148294 111554 148350
rect 111622 148294 111678 148350
rect 111250 148170 111306 148226
rect 111374 148170 111430 148226
rect 111498 148170 111554 148226
rect 111622 148170 111678 148226
rect 111250 148046 111306 148102
rect 111374 148046 111430 148102
rect 111498 148046 111554 148102
rect 111622 148046 111678 148102
rect 111250 147922 111306 147978
rect 111374 147922 111430 147978
rect 111498 147922 111554 147978
rect 111622 147922 111678 147978
rect 111250 130294 111306 130350
rect 111374 130294 111430 130350
rect 111498 130294 111554 130350
rect 111622 130294 111678 130350
rect 111250 130170 111306 130226
rect 111374 130170 111430 130226
rect 111498 130170 111554 130226
rect 111622 130170 111678 130226
rect 111250 130046 111306 130102
rect 111374 130046 111430 130102
rect 111498 130046 111554 130102
rect 111622 130046 111678 130102
rect 111250 129922 111306 129978
rect 111374 129922 111430 129978
rect 111498 129922 111554 129978
rect 111622 129922 111678 129978
rect 111250 112294 111306 112350
rect 111374 112294 111430 112350
rect 111498 112294 111554 112350
rect 111622 112294 111678 112350
rect 111250 112170 111306 112226
rect 111374 112170 111430 112226
rect 111498 112170 111554 112226
rect 111622 112170 111678 112226
rect 111250 112046 111306 112102
rect 111374 112046 111430 112102
rect 111498 112046 111554 112102
rect 111622 112046 111678 112102
rect 111250 111922 111306 111978
rect 111374 111922 111430 111978
rect 111498 111922 111554 111978
rect 111622 111922 111678 111978
rect 114970 154294 115026 154350
rect 115094 154294 115150 154350
rect 115218 154294 115274 154350
rect 115342 154294 115398 154350
rect 114970 154170 115026 154226
rect 115094 154170 115150 154226
rect 115218 154170 115274 154226
rect 115342 154170 115398 154226
rect 114970 154046 115026 154102
rect 115094 154046 115150 154102
rect 115218 154046 115274 154102
rect 115342 154046 115398 154102
rect 114970 153922 115026 153978
rect 115094 153922 115150 153978
rect 115218 153922 115274 153978
rect 115342 153922 115398 153978
rect 114970 136294 115026 136350
rect 115094 136294 115150 136350
rect 115218 136294 115274 136350
rect 115342 136294 115398 136350
rect 114970 136170 115026 136226
rect 115094 136170 115150 136226
rect 115218 136170 115274 136226
rect 115342 136170 115398 136226
rect 114970 136046 115026 136102
rect 115094 136046 115150 136102
rect 115218 136046 115274 136102
rect 115342 136046 115398 136102
rect 114970 135922 115026 135978
rect 115094 135922 115150 135978
rect 115218 135922 115274 135978
rect 115342 135922 115398 135978
rect 114970 118294 115026 118350
rect 115094 118294 115150 118350
rect 115218 118294 115274 118350
rect 115342 118294 115398 118350
rect 114970 118170 115026 118226
rect 115094 118170 115150 118226
rect 115218 118170 115274 118226
rect 115342 118170 115398 118226
rect 114970 118046 115026 118102
rect 115094 118046 115150 118102
rect 115218 118046 115274 118102
rect 115342 118046 115398 118102
rect 114970 117922 115026 117978
rect 115094 117922 115150 117978
rect 115218 117922 115274 117978
rect 115342 117922 115398 117978
rect 129250 148294 129306 148350
rect 129374 148294 129430 148350
rect 129498 148294 129554 148350
rect 129622 148294 129678 148350
rect 129250 148170 129306 148226
rect 129374 148170 129430 148226
rect 129498 148170 129554 148226
rect 129622 148170 129678 148226
rect 129250 148046 129306 148102
rect 129374 148046 129430 148102
rect 129498 148046 129554 148102
rect 129622 148046 129678 148102
rect 129250 147922 129306 147978
rect 129374 147922 129430 147978
rect 129498 147922 129554 147978
rect 129622 147922 129678 147978
rect 129250 130294 129306 130350
rect 129374 130294 129430 130350
rect 129498 130294 129554 130350
rect 129622 130294 129678 130350
rect 129250 130170 129306 130226
rect 129374 130170 129430 130226
rect 129498 130170 129554 130226
rect 129622 130170 129678 130226
rect 129250 130046 129306 130102
rect 129374 130046 129430 130102
rect 129498 130046 129554 130102
rect 129622 130046 129678 130102
rect 129250 129922 129306 129978
rect 129374 129922 129430 129978
rect 129498 129922 129554 129978
rect 129622 129922 129678 129978
rect 129250 112294 129306 112350
rect 129374 112294 129430 112350
rect 129498 112294 129554 112350
rect 129622 112294 129678 112350
rect 129250 112170 129306 112226
rect 129374 112170 129430 112226
rect 129498 112170 129554 112226
rect 129622 112170 129678 112226
rect 129250 112046 129306 112102
rect 129374 112046 129430 112102
rect 129498 112046 129554 112102
rect 129622 112046 129678 112102
rect 129250 111922 129306 111978
rect 129374 111922 129430 111978
rect 129498 111922 129554 111978
rect 129622 111922 129678 111978
rect 132970 154294 133026 154350
rect 133094 154294 133150 154350
rect 133218 154294 133274 154350
rect 133342 154294 133398 154350
rect 132970 154170 133026 154226
rect 133094 154170 133150 154226
rect 133218 154170 133274 154226
rect 133342 154170 133398 154226
rect 132970 154046 133026 154102
rect 133094 154046 133150 154102
rect 133218 154046 133274 154102
rect 133342 154046 133398 154102
rect 132970 153922 133026 153978
rect 133094 153922 133150 153978
rect 133218 153922 133274 153978
rect 133342 153922 133398 153978
rect 132970 136294 133026 136350
rect 133094 136294 133150 136350
rect 133218 136294 133274 136350
rect 133342 136294 133398 136350
rect 132970 136170 133026 136226
rect 133094 136170 133150 136226
rect 133218 136170 133274 136226
rect 133342 136170 133398 136226
rect 132970 136046 133026 136102
rect 133094 136046 133150 136102
rect 133218 136046 133274 136102
rect 133342 136046 133398 136102
rect 132970 135922 133026 135978
rect 133094 135922 133150 135978
rect 133218 135922 133274 135978
rect 133342 135922 133398 135978
rect 132970 118294 133026 118350
rect 133094 118294 133150 118350
rect 133218 118294 133274 118350
rect 133342 118294 133398 118350
rect 132970 118170 133026 118226
rect 133094 118170 133150 118226
rect 133218 118170 133274 118226
rect 133342 118170 133398 118226
rect 132970 118046 133026 118102
rect 133094 118046 133150 118102
rect 133218 118046 133274 118102
rect 133342 118046 133398 118102
rect 132970 117922 133026 117978
rect 133094 117922 133150 117978
rect 133218 117922 133274 117978
rect 133342 117922 133398 117978
rect 147250 148294 147306 148350
rect 147374 148294 147430 148350
rect 147498 148294 147554 148350
rect 147622 148294 147678 148350
rect 147250 148170 147306 148226
rect 147374 148170 147430 148226
rect 147498 148170 147554 148226
rect 147622 148170 147678 148226
rect 147250 148046 147306 148102
rect 147374 148046 147430 148102
rect 147498 148046 147554 148102
rect 147622 148046 147678 148102
rect 147250 147922 147306 147978
rect 147374 147922 147430 147978
rect 147498 147922 147554 147978
rect 147622 147922 147678 147978
rect 147250 130294 147306 130350
rect 147374 130294 147430 130350
rect 147498 130294 147554 130350
rect 147622 130294 147678 130350
rect 147250 130170 147306 130226
rect 147374 130170 147430 130226
rect 147498 130170 147554 130226
rect 147622 130170 147678 130226
rect 147250 130046 147306 130102
rect 147374 130046 147430 130102
rect 147498 130046 147554 130102
rect 147622 130046 147678 130102
rect 147250 129922 147306 129978
rect 147374 129922 147430 129978
rect 147498 129922 147554 129978
rect 147622 129922 147678 129978
rect 147250 112294 147306 112350
rect 147374 112294 147430 112350
rect 147498 112294 147554 112350
rect 147622 112294 147678 112350
rect 147250 112170 147306 112226
rect 147374 112170 147430 112226
rect 147498 112170 147554 112226
rect 147622 112170 147678 112226
rect 147250 112046 147306 112102
rect 147374 112046 147430 112102
rect 147498 112046 147554 112102
rect 147622 112046 147678 112102
rect 147250 111922 147306 111978
rect 147374 111922 147430 111978
rect 147498 111922 147554 111978
rect 147622 111922 147678 111978
rect 150970 154294 151026 154350
rect 151094 154294 151150 154350
rect 151218 154294 151274 154350
rect 151342 154294 151398 154350
rect 150970 154170 151026 154226
rect 151094 154170 151150 154226
rect 151218 154170 151274 154226
rect 151342 154170 151398 154226
rect 150970 154046 151026 154102
rect 151094 154046 151150 154102
rect 151218 154046 151274 154102
rect 151342 154046 151398 154102
rect 150970 153922 151026 153978
rect 151094 153922 151150 153978
rect 151218 153922 151274 153978
rect 151342 153922 151398 153978
rect 150970 136294 151026 136350
rect 151094 136294 151150 136350
rect 151218 136294 151274 136350
rect 151342 136294 151398 136350
rect 150970 136170 151026 136226
rect 151094 136170 151150 136226
rect 151218 136170 151274 136226
rect 151342 136170 151398 136226
rect 150970 136046 151026 136102
rect 151094 136046 151150 136102
rect 151218 136046 151274 136102
rect 151342 136046 151398 136102
rect 150970 135922 151026 135978
rect 151094 135922 151150 135978
rect 151218 135922 151274 135978
rect 151342 135922 151398 135978
rect 150970 118294 151026 118350
rect 151094 118294 151150 118350
rect 151218 118294 151274 118350
rect 151342 118294 151398 118350
rect 150970 118170 151026 118226
rect 151094 118170 151150 118226
rect 151218 118170 151274 118226
rect 151342 118170 151398 118226
rect 150970 118046 151026 118102
rect 151094 118046 151150 118102
rect 151218 118046 151274 118102
rect 151342 118046 151398 118102
rect 150970 117922 151026 117978
rect 151094 117922 151150 117978
rect 151218 117922 151274 117978
rect 151342 117922 151398 117978
rect 165250 148294 165306 148350
rect 165374 148294 165430 148350
rect 165498 148294 165554 148350
rect 165622 148294 165678 148350
rect 165250 148170 165306 148226
rect 165374 148170 165430 148226
rect 165498 148170 165554 148226
rect 165622 148170 165678 148226
rect 165250 148046 165306 148102
rect 165374 148046 165430 148102
rect 165498 148046 165554 148102
rect 165622 148046 165678 148102
rect 165250 147922 165306 147978
rect 165374 147922 165430 147978
rect 165498 147922 165554 147978
rect 165622 147922 165678 147978
rect 165250 130294 165306 130350
rect 165374 130294 165430 130350
rect 165498 130294 165554 130350
rect 165622 130294 165678 130350
rect 165250 130170 165306 130226
rect 165374 130170 165430 130226
rect 165498 130170 165554 130226
rect 165622 130170 165678 130226
rect 165250 130046 165306 130102
rect 165374 130046 165430 130102
rect 165498 130046 165554 130102
rect 165622 130046 165678 130102
rect 165250 129922 165306 129978
rect 165374 129922 165430 129978
rect 165498 129922 165554 129978
rect 165622 129922 165678 129978
rect 165250 112294 165306 112350
rect 165374 112294 165430 112350
rect 165498 112294 165554 112350
rect 165622 112294 165678 112350
rect 165250 112170 165306 112226
rect 165374 112170 165430 112226
rect 165498 112170 165554 112226
rect 165622 112170 165678 112226
rect 165250 112046 165306 112102
rect 165374 112046 165430 112102
rect 165498 112046 165554 112102
rect 165622 112046 165678 112102
rect 165250 111922 165306 111978
rect 165374 111922 165430 111978
rect 165498 111922 165554 111978
rect 165622 111922 165678 111978
rect 168970 154294 169026 154350
rect 169094 154294 169150 154350
rect 169218 154294 169274 154350
rect 169342 154294 169398 154350
rect 168970 154170 169026 154226
rect 169094 154170 169150 154226
rect 169218 154170 169274 154226
rect 169342 154170 169398 154226
rect 168970 154046 169026 154102
rect 169094 154046 169150 154102
rect 169218 154046 169274 154102
rect 169342 154046 169398 154102
rect 168970 153922 169026 153978
rect 169094 153922 169150 153978
rect 169218 153922 169274 153978
rect 169342 153922 169398 153978
rect 168970 136294 169026 136350
rect 169094 136294 169150 136350
rect 169218 136294 169274 136350
rect 169342 136294 169398 136350
rect 168970 136170 169026 136226
rect 169094 136170 169150 136226
rect 169218 136170 169274 136226
rect 169342 136170 169398 136226
rect 168970 136046 169026 136102
rect 169094 136046 169150 136102
rect 169218 136046 169274 136102
rect 169342 136046 169398 136102
rect 168970 135922 169026 135978
rect 169094 135922 169150 135978
rect 169218 135922 169274 135978
rect 169342 135922 169398 135978
rect 168970 118294 169026 118350
rect 169094 118294 169150 118350
rect 169218 118294 169274 118350
rect 169342 118294 169398 118350
rect 168970 118170 169026 118226
rect 169094 118170 169150 118226
rect 169218 118170 169274 118226
rect 169342 118170 169398 118226
rect 168970 118046 169026 118102
rect 169094 118046 169150 118102
rect 169218 118046 169274 118102
rect 169342 118046 169398 118102
rect 168970 117922 169026 117978
rect 169094 117922 169150 117978
rect 169218 117922 169274 117978
rect 169342 117922 169398 117978
rect 183250 148294 183306 148350
rect 183374 148294 183430 148350
rect 183498 148294 183554 148350
rect 183622 148294 183678 148350
rect 183250 148170 183306 148226
rect 183374 148170 183430 148226
rect 183498 148170 183554 148226
rect 183622 148170 183678 148226
rect 183250 148046 183306 148102
rect 183374 148046 183430 148102
rect 183498 148046 183554 148102
rect 183622 148046 183678 148102
rect 183250 147922 183306 147978
rect 183374 147922 183430 147978
rect 183498 147922 183554 147978
rect 183622 147922 183678 147978
rect 183250 130294 183306 130350
rect 183374 130294 183430 130350
rect 183498 130294 183554 130350
rect 183622 130294 183678 130350
rect 183250 130170 183306 130226
rect 183374 130170 183430 130226
rect 183498 130170 183554 130226
rect 183622 130170 183678 130226
rect 183250 130046 183306 130102
rect 183374 130046 183430 130102
rect 183498 130046 183554 130102
rect 183622 130046 183678 130102
rect 183250 129922 183306 129978
rect 183374 129922 183430 129978
rect 183498 129922 183554 129978
rect 183622 129922 183678 129978
rect 183250 112294 183306 112350
rect 183374 112294 183430 112350
rect 183498 112294 183554 112350
rect 183622 112294 183678 112350
rect 183250 112170 183306 112226
rect 183374 112170 183430 112226
rect 183498 112170 183554 112226
rect 183622 112170 183678 112226
rect 183250 112046 183306 112102
rect 183374 112046 183430 112102
rect 183498 112046 183554 112102
rect 183622 112046 183678 112102
rect 183250 111922 183306 111978
rect 183374 111922 183430 111978
rect 183498 111922 183554 111978
rect 183622 111922 183678 111978
rect 42970 100294 43026 100350
rect 43094 100294 43150 100350
rect 43218 100294 43274 100350
rect 43342 100294 43398 100350
rect 42970 100170 43026 100226
rect 43094 100170 43150 100226
rect 43218 100170 43274 100226
rect 43342 100170 43398 100226
rect 42970 100046 43026 100102
rect 43094 100046 43150 100102
rect 43218 100046 43274 100102
rect 43342 100046 43398 100102
rect 42970 99922 43026 99978
rect 43094 99922 43150 99978
rect 43218 99922 43274 99978
rect 43342 99922 43398 99978
rect 42970 82294 43026 82350
rect 43094 82294 43150 82350
rect 43218 82294 43274 82350
rect 43342 82294 43398 82350
rect 42970 82170 43026 82226
rect 43094 82170 43150 82226
rect 43218 82170 43274 82226
rect 43342 82170 43398 82226
rect 42970 82046 43026 82102
rect 43094 82046 43150 82102
rect 43218 82046 43274 82102
rect 43342 82046 43398 82102
rect 42970 81922 43026 81978
rect 43094 81922 43150 81978
rect 43218 81922 43274 81978
rect 43342 81922 43398 81978
rect 39250 58294 39306 58350
rect 39374 58294 39430 58350
rect 39498 58294 39554 58350
rect 39622 58294 39678 58350
rect 39250 58170 39306 58226
rect 39374 58170 39430 58226
rect 39498 58170 39554 58226
rect 39622 58170 39678 58226
rect 39250 58046 39306 58102
rect 39374 58046 39430 58102
rect 39498 58046 39554 58102
rect 39622 58046 39678 58102
rect 39250 57922 39306 57978
rect 39374 57922 39430 57978
rect 39498 57922 39554 57978
rect 39622 57922 39678 57978
rect 39250 40294 39306 40350
rect 39374 40294 39430 40350
rect 39498 40294 39554 40350
rect 39622 40294 39678 40350
rect 39250 40170 39306 40226
rect 39374 40170 39430 40226
rect 39498 40170 39554 40226
rect 39622 40170 39678 40226
rect 39250 40046 39306 40102
rect 39374 40046 39430 40102
rect 39498 40046 39554 40102
rect 39622 40046 39678 40102
rect 39250 39922 39306 39978
rect 39374 39922 39430 39978
rect 39498 39922 39554 39978
rect 39622 39922 39678 39978
rect 39250 22294 39306 22350
rect 39374 22294 39430 22350
rect 39498 22294 39554 22350
rect 39622 22294 39678 22350
rect 39250 22170 39306 22226
rect 39374 22170 39430 22226
rect 39498 22170 39554 22226
rect 39622 22170 39678 22226
rect 39250 22046 39306 22102
rect 39374 22046 39430 22102
rect 39498 22046 39554 22102
rect 39622 22046 39678 22102
rect 39250 21922 39306 21978
rect 39374 21922 39430 21978
rect 39498 21922 39554 21978
rect 39622 21922 39678 21978
rect 24970 -1176 25026 -1120
rect 25094 -1176 25150 -1120
rect 25218 -1176 25274 -1120
rect 25342 -1176 25398 -1120
rect 24970 -1300 25026 -1244
rect 25094 -1300 25150 -1244
rect 25218 -1300 25274 -1244
rect 25342 -1300 25398 -1244
rect 24970 -1424 25026 -1368
rect 25094 -1424 25150 -1368
rect 25218 -1424 25274 -1368
rect 25342 -1424 25398 -1368
rect 24970 -1548 25026 -1492
rect 25094 -1548 25150 -1492
rect 25218 -1548 25274 -1492
rect 25342 -1548 25398 -1492
rect 183250 94294 183306 94350
rect 183374 94294 183430 94350
rect 183498 94294 183554 94350
rect 183622 94294 183678 94350
rect 183250 94170 183306 94226
rect 183374 94170 183430 94226
rect 183498 94170 183554 94226
rect 183622 94170 183678 94226
rect 183250 94046 183306 94102
rect 183374 94046 183430 94102
rect 183498 94046 183554 94102
rect 183622 94046 183678 94102
rect 183250 93922 183306 93978
rect 183374 93922 183430 93978
rect 183498 93922 183554 93978
rect 183622 93922 183678 93978
rect 57250 76294 57306 76350
rect 57374 76294 57430 76350
rect 57498 76294 57554 76350
rect 57622 76294 57678 76350
rect 57250 76170 57306 76226
rect 57374 76170 57430 76226
rect 57498 76170 57554 76226
rect 57622 76170 57678 76226
rect 57250 76046 57306 76102
rect 57374 76046 57430 76102
rect 57498 76046 57554 76102
rect 57622 76046 57678 76102
rect 57250 75922 57306 75978
rect 57374 75922 57430 75978
rect 57498 75922 57554 75978
rect 57622 75922 57678 75978
rect 42970 64294 43026 64350
rect 43094 64294 43150 64350
rect 43218 64294 43274 64350
rect 43342 64294 43398 64350
rect 42970 64170 43026 64226
rect 43094 64170 43150 64226
rect 43218 64170 43274 64226
rect 43342 64170 43398 64226
rect 42970 64046 43026 64102
rect 43094 64046 43150 64102
rect 43218 64046 43274 64102
rect 43342 64046 43398 64102
rect 42970 63922 43026 63978
rect 43094 63922 43150 63978
rect 43218 63922 43274 63978
rect 43342 63922 43398 63978
rect 42970 46294 43026 46350
rect 43094 46294 43150 46350
rect 43218 46294 43274 46350
rect 43342 46294 43398 46350
rect 42970 46170 43026 46226
rect 43094 46170 43150 46226
rect 43218 46170 43274 46226
rect 43342 46170 43398 46226
rect 42970 46046 43026 46102
rect 43094 46046 43150 46102
rect 43218 46046 43274 46102
rect 43342 46046 43398 46102
rect 42970 45922 43026 45978
rect 43094 45922 43150 45978
rect 43218 45922 43274 45978
rect 43342 45922 43398 45978
rect 42970 28294 43026 28350
rect 43094 28294 43150 28350
rect 43218 28294 43274 28350
rect 43342 28294 43398 28350
rect 42970 28170 43026 28226
rect 43094 28170 43150 28226
rect 43218 28170 43274 28226
rect 43342 28170 43398 28226
rect 42970 28046 43026 28102
rect 43094 28046 43150 28102
rect 43218 28046 43274 28102
rect 43342 28046 43398 28102
rect 42970 27922 43026 27978
rect 43094 27922 43150 27978
rect 43218 27922 43274 27978
rect 43342 27922 43398 27978
rect 39250 4294 39306 4350
rect 39374 4294 39430 4350
rect 39498 4294 39554 4350
rect 39622 4294 39678 4350
rect 39250 4170 39306 4226
rect 39374 4170 39430 4226
rect 39498 4170 39554 4226
rect 39622 4170 39678 4226
rect 39250 4046 39306 4102
rect 39374 4046 39430 4102
rect 39498 4046 39554 4102
rect 39622 4046 39678 4102
rect 39250 3922 39306 3978
rect 39374 3922 39430 3978
rect 39498 3922 39554 3978
rect 39622 3922 39678 3978
rect 39250 -216 39306 -160
rect 39374 -216 39430 -160
rect 39498 -216 39554 -160
rect 39622 -216 39678 -160
rect 39250 -340 39306 -284
rect 39374 -340 39430 -284
rect 39498 -340 39554 -284
rect 39622 -340 39678 -284
rect 39250 -464 39306 -408
rect 39374 -464 39430 -408
rect 39498 -464 39554 -408
rect 39622 -464 39678 -408
rect 39250 -588 39306 -532
rect 39374 -588 39430 -532
rect 39498 -588 39554 -532
rect 39622 -588 39678 -532
rect 57250 58294 57306 58350
rect 57374 58294 57430 58350
rect 57498 58294 57554 58350
rect 57622 58294 57678 58350
rect 57250 58170 57306 58226
rect 57374 58170 57430 58226
rect 57498 58170 57554 58226
rect 57622 58170 57678 58226
rect 57250 58046 57306 58102
rect 57374 58046 57430 58102
rect 57498 58046 57554 58102
rect 57622 58046 57678 58102
rect 57250 57922 57306 57978
rect 57374 57922 57430 57978
rect 57498 57922 57554 57978
rect 57622 57922 57678 57978
rect 57250 40294 57306 40350
rect 57374 40294 57430 40350
rect 57498 40294 57554 40350
rect 57622 40294 57678 40350
rect 57250 40170 57306 40226
rect 57374 40170 57430 40226
rect 57498 40170 57554 40226
rect 57622 40170 57678 40226
rect 57250 40046 57306 40102
rect 57374 40046 57430 40102
rect 57498 40046 57554 40102
rect 57622 40046 57678 40102
rect 57250 39922 57306 39978
rect 57374 39922 57430 39978
rect 57498 39922 57554 39978
rect 57622 39922 57678 39978
rect 57250 22294 57306 22350
rect 57374 22294 57430 22350
rect 57498 22294 57554 22350
rect 57622 22294 57678 22350
rect 57250 22170 57306 22226
rect 57374 22170 57430 22226
rect 57498 22170 57554 22226
rect 57622 22170 57678 22226
rect 57250 22046 57306 22102
rect 57374 22046 57430 22102
rect 57498 22046 57554 22102
rect 57622 22046 57678 22102
rect 57250 21922 57306 21978
rect 57374 21922 57430 21978
rect 57498 21922 57554 21978
rect 57622 21922 57678 21978
rect 42970 10294 43026 10350
rect 43094 10294 43150 10350
rect 43218 10294 43274 10350
rect 43342 10294 43398 10350
rect 42970 10170 43026 10226
rect 43094 10170 43150 10226
rect 43218 10170 43274 10226
rect 43342 10170 43398 10226
rect 42970 10046 43026 10102
rect 43094 10046 43150 10102
rect 43218 10046 43274 10102
rect 43342 10046 43398 10102
rect 42970 9922 43026 9978
rect 43094 9922 43150 9978
rect 43218 9922 43274 9978
rect 43342 9922 43398 9978
rect 42970 -1176 43026 -1120
rect 43094 -1176 43150 -1120
rect 43218 -1176 43274 -1120
rect 43342 -1176 43398 -1120
rect 42970 -1300 43026 -1244
rect 43094 -1300 43150 -1244
rect 43218 -1300 43274 -1244
rect 43342 -1300 43398 -1244
rect 42970 -1424 43026 -1368
rect 43094 -1424 43150 -1368
rect 43218 -1424 43274 -1368
rect 43342 -1424 43398 -1368
rect 42970 -1548 43026 -1492
rect 43094 -1548 43150 -1492
rect 43218 -1548 43274 -1492
rect 43342 -1548 43398 -1492
rect 60970 64294 61026 64350
rect 61094 64294 61150 64350
rect 61218 64294 61274 64350
rect 61342 64294 61398 64350
rect 60970 64170 61026 64226
rect 61094 64170 61150 64226
rect 61218 64170 61274 64226
rect 61342 64170 61398 64226
rect 60970 64046 61026 64102
rect 61094 64046 61150 64102
rect 61218 64046 61274 64102
rect 61342 64046 61398 64102
rect 60970 63922 61026 63978
rect 61094 63922 61150 63978
rect 61218 63922 61274 63978
rect 61342 63922 61398 63978
rect 75250 76294 75306 76350
rect 75374 76294 75430 76350
rect 75498 76294 75554 76350
rect 75622 76294 75678 76350
rect 75250 76170 75306 76226
rect 75374 76170 75430 76226
rect 75498 76170 75554 76226
rect 75622 76170 75678 76226
rect 75250 76046 75306 76102
rect 75374 76046 75430 76102
rect 75498 76046 75554 76102
rect 75622 76046 75678 76102
rect 75250 75922 75306 75978
rect 75374 75922 75430 75978
rect 75498 75922 75554 75978
rect 75622 75922 75678 75978
rect 75250 58294 75306 58350
rect 75374 58294 75430 58350
rect 75498 58294 75554 58350
rect 75622 58294 75678 58350
rect 75250 58170 75306 58226
rect 75374 58170 75430 58226
rect 75498 58170 75554 58226
rect 75622 58170 75678 58226
rect 75250 58046 75306 58102
rect 75374 58046 75430 58102
rect 75498 58046 75554 58102
rect 75622 58046 75678 58102
rect 75250 57922 75306 57978
rect 75374 57922 75430 57978
rect 75498 57922 75554 57978
rect 75622 57922 75678 57978
rect 60970 46294 61026 46350
rect 61094 46294 61150 46350
rect 61218 46294 61274 46350
rect 61342 46294 61398 46350
rect 60970 46170 61026 46226
rect 61094 46170 61150 46226
rect 61218 46170 61274 46226
rect 61342 46170 61398 46226
rect 60970 46046 61026 46102
rect 61094 46046 61150 46102
rect 61218 46046 61274 46102
rect 61342 46046 61398 46102
rect 60970 45922 61026 45978
rect 61094 45922 61150 45978
rect 61218 45922 61274 45978
rect 61342 45922 61398 45978
rect 60970 28294 61026 28350
rect 61094 28294 61150 28350
rect 61218 28294 61274 28350
rect 61342 28294 61398 28350
rect 60970 28170 61026 28226
rect 61094 28170 61150 28226
rect 61218 28170 61274 28226
rect 61342 28170 61398 28226
rect 60970 28046 61026 28102
rect 61094 28046 61150 28102
rect 61218 28046 61274 28102
rect 61342 28046 61398 28102
rect 60970 27922 61026 27978
rect 61094 27922 61150 27978
rect 61218 27922 61274 27978
rect 61342 27922 61398 27978
rect 57250 4294 57306 4350
rect 57374 4294 57430 4350
rect 57498 4294 57554 4350
rect 57622 4294 57678 4350
rect 57250 4170 57306 4226
rect 57374 4170 57430 4226
rect 57498 4170 57554 4226
rect 57622 4170 57678 4226
rect 57250 4046 57306 4102
rect 57374 4046 57430 4102
rect 57498 4046 57554 4102
rect 57622 4046 57678 4102
rect 57250 3922 57306 3978
rect 57374 3922 57430 3978
rect 57498 3922 57554 3978
rect 57622 3922 57678 3978
rect 57250 -216 57306 -160
rect 57374 -216 57430 -160
rect 57498 -216 57554 -160
rect 57622 -216 57678 -160
rect 57250 -340 57306 -284
rect 57374 -340 57430 -284
rect 57498 -340 57554 -284
rect 57622 -340 57678 -284
rect 57250 -464 57306 -408
rect 57374 -464 57430 -408
rect 57498 -464 57554 -408
rect 57622 -464 57678 -408
rect 57250 -588 57306 -532
rect 57374 -588 57430 -532
rect 57498 -588 57554 -532
rect 57622 -588 57678 -532
rect 75250 40294 75306 40350
rect 75374 40294 75430 40350
rect 75498 40294 75554 40350
rect 75622 40294 75678 40350
rect 75250 40170 75306 40226
rect 75374 40170 75430 40226
rect 75498 40170 75554 40226
rect 75622 40170 75678 40226
rect 75250 40046 75306 40102
rect 75374 40046 75430 40102
rect 75498 40046 75554 40102
rect 75622 40046 75678 40102
rect 75250 39922 75306 39978
rect 75374 39922 75430 39978
rect 75498 39922 75554 39978
rect 75622 39922 75678 39978
rect 75250 22294 75306 22350
rect 75374 22294 75430 22350
rect 75498 22294 75554 22350
rect 75622 22294 75678 22350
rect 75250 22170 75306 22226
rect 75374 22170 75430 22226
rect 75498 22170 75554 22226
rect 75622 22170 75678 22226
rect 75250 22046 75306 22102
rect 75374 22046 75430 22102
rect 75498 22046 75554 22102
rect 75622 22046 75678 22102
rect 75250 21922 75306 21978
rect 75374 21922 75430 21978
rect 75498 21922 75554 21978
rect 75622 21922 75678 21978
rect 60970 10294 61026 10350
rect 61094 10294 61150 10350
rect 61218 10294 61274 10350
rect 61342 10294 61398 10350
rect 60970 10170 61026 10226
rect 61094 10170 61150 10226
rect 61218 10170 61274 10226
rect 61342 10170 61398 10226
rect 60970 10046 61026 10102
rect 61094 10046 61150 10102
rect 61218 10046 61274 10102
rect 61342 10046 61398 10102
rect 60970 9922 61026 9978
rect 61094 9922 61150 9978
rect 61218 9922 61274 9978
rect 61342 9922 61398 9978
rect 60970 -1176 61026 -1120
rect 61094 -1176 61150 -1120
rect 61218 -1176 61274 -1120
rect 61342 -1176 61398 -1120
rect 60970 -1300 61026 -1244
rect 61094 -1300 61150 -1244
rect 61218 -1300 61274 -1244
rect 61342 -1300 61398 -1244
rect 60970 -1424 61026 -1368
rect 61094 -1424 61150 -1368
rect 61218 -1424 61274 -1368
rect 61342 -1424 61398 -1368
rect 60970 -1548 61026 -1492
rect 61094 -1548 61150 -1492
rect 61218 -1548 61274 -1492
rect 61342 -1548 61398 -1492
rect 75250 4294 75306 4350
rect 75374 4294 75430 4350
rect 75498 4294 75554 4350
rect 75622 4294 75678 4350
rect 75250 4170 75306 4226
rect 75374 4170 75430 4226
rect 75498 4170 75554 4226
rect 75622 4170 75678 4226
rect 75250 4046 75306 4102
rect 75374 4046 75430 4102
rect 75498 4046 75554 4102
rect 75622 4046 75678 4102
rect 75250 3922 75306 3978
rect 75374 3922 75430 3978
rect 75498 3922 75554 3978
rect 75622 3922 75678 3978
rect 75250 -216 75306 -160
rect 75374 -216 75430 -160
rect 75498 -216 75554 -160
rect 75622 -216 75678 -160
rect 75250 -340 75306 -284
rect 75374 -340 75430 -284
rect 75498 -340 75554 -284
rect 75622 -340 75678 -284
rect 75250 -464 75306 -408
rect 75374 -464 75430 -408
rect 75498 -464 75554 -408
rect 75622 -464 75678 -408
rect 75250 -588 75306 -532
rect 75374 -588 75430 -532
rect 75498 -588 75554 -532
rect 75622 -588 75678 -532
rect 78970 64294 79026 64350
rect 79094 64294 79150 64350
rect 79218 64294 79274 64350
rect 79342 64294 79398 64350
rect 78970 64170 79026 64226
rect 79094 64170 79150 64226
rect 79218 64170 79274 64226
rect 79342 64170 79398 64226
rect 78970 64046 79026 64102
rect 79094 64046 79150 64102
rect 79218 64046 79274 64102
rect 79342 64046 79398 64102
rect 78970 63922 79026 63978
rect 79094 63922 79150 63978
rect 79218 63922 79274 63978
rect 79342 63922 79398 63978
rect 78970 46294 79026 46350
rect 79094 46294 79150 46350
rect 79218 46294 79274 46350
rect 79342 46294 79398 46350
rect 78970 46170 79026 46226
rect 79094 46170 79150 46226
rect 79218 46170 79274 46226
rect 79342 46170 79398 46226
rect 78970 46046 79026 46102
rect 79094 46046 79150 46102
rect 79218 46046 79274 46102
rect 79342 46046 79398 46102
rect 78970 45922 79026 45978
rect 79094 45922 79150 45978
rect 79218 45922 79274 45978
rect 79342 45922 79398 45978
rect 78970 28294 79026 28350
rect 79094 28294 79150 28350
rect 79218 28294 79274 28350
rect 79342 28294 79398 28350
rect 78970 28170 79026 28226
rect 79094 28170 79150 28226
rect 79218 28170 79274 28226
rect 79342 28170 79398 28226
rect 78970 28046 79026 28102
rect 79094 28046 79150 28102
rect 79218 28046 79274 28102
rect 79342 28046 79398 28102
rect 78970 27922 79026 27978
rect 79094 27922 79150 27978
rect 79218 27922 79274 27978
rect 79342 27922 79398 27978
rect 78970 10294 79026 10350
rect 79094 10294 79150 10350
rect 79218 10294 79274 10350
rect 79342 10294 79398 10350
rect 78970 10170 79026 10226
rect 79094 10170 79150 10226
rect 79218 10170 79274 10226
rect 79342 10170 79398 10226
rect 78970 10046 79026 10102
rect 79094 10046 79150 10102
rect 79218 10046 79274 10102
rect 79342 10046 79398 10102
rect 78970 9922 79026 9978
rect 79094 9922 79150 9978
rect 79218 9922 79274 9978
rect 79342 9922 79398 9978
rect 78970 -1176 79026 -1120
rect 79094 -1176 79150 -1120
rect 79218 -1176 79274 -1120
rect 79342 -1176 79398 -1120
rect 78970 -1300 79026 -1244
rect 79094 -1300 79150 -1244
rect 79218 -1300 79274 -1244
rect 79342 -1300 79398 -1244
rect 78970 -1424 79026 -1368
rect 79094 -1424 79150 -1368
rect 79218 -1424 79274 -1368
rect 79342 -1424 79398 -1368
rect 78970 -1548 79026 -1492
rect 79094 -1548 79150 -1492
rect 79218 -1548 79274 -1492
rect 79342 -1548 79398 -1492
rect 93250 76294 93306 76350
rect 93374 76294 93430 76350
rect 93498 76294 93554 76350
rect 93622 76294 93678 76350
rect 93250 76170 93306 76226
rect 93374 76170 93430 76226
rect 93498 76170 93554 76226
rect 93622 76170 93678 76226
rect 93250 76046 93306 76102
rect 93374 76046 93430 76102
rect 93498 76046 93554 76102
rect 93622 76046 93678 76102
rect 93250 75922 93306 75978
rect 93374 75922 93430 75978
rect 93498 75922 93554 75978
rect 93622 75922 93678 75978
rect 93250 58294 93306 58350
rect 93374 58294 93430 58350
rect 93498 58294 93554 58350
rect 93622 58294 93678 58350
rect 93250 58170 93306 58226
rect 93374 58170 93430 58226
rect 93498 58170 93554 58226
rect 93622 58170 93678 58226
rect 93250 58046 93306 58102
rect 93374 58046 93430 58102
rect 93498 58046 93554 58102
rect 93622 58046 93678 58102
rect 93250 57922 93306 57978
rect 93374 57922 93430 57978
rect 93498 57922 93554 57978
rect 93622 57922 93678 57978
rect 93250 40294 93306 40350
rect 93374 40294 93430 40350
rect 93498 40294 93554 40350
rect 93622 40294 93678 40350
rect 93250 40170 93306 40226
rect 93374 40170 93430 40226
rect 93498 40170 93554 40226
rect 93622 40170 93678 40226
rect 93250 40046 93306 40102
rect 93374 40046 93430 40102
rect 93498 40046 93554 40102
rect 93622 40046 93678 40102
rect 93250 39922 93306 39978
rect 93374 39922 93430 39978
rect 93498 39922 93554 39978
rect 93622 39922 93678 39978
rect 93250 22294 93306 22350
rect 93374 22294 93430 22350
rect 93498 22294 93554 22350
rect 93622 22294 93678 22350
rect 93250 22170 93306 22226
rect 93374 22170 93430 22226
rect 93498 22170 93554 22226
rect 93622 22170 93678 22226
rect 93250 22046 93306 22102
rect 93374 22046 93430 22102
rect 93498 22046 93554 22102
rect 93622 22046 93678 22102
rect 93250 21922 93306 21978
rect 93374 21922 93430 21978
rect 93498 21922 93554 21978
rect 93622 21922 93678 21978
rect 93250 4294 93306 4350
rect 93374 4294 93430 4350
rect 93498 4294 93554 4350
rect 93622 4294 93678 4350
rect 93250 4170 93306 4226
rect 93374 4170 93430 4226
rect 93498 4170 93554 4226
rect 93622 4170 93678 4226
rect 93250 4046 93306 4102
rect 93374 4046 93430 4102
rect 93498 4046 93554 4102
rect 93622 4046 93678 4102
rect 93250 3922 93306 3978
rect 93374 3922 93430 3978
rect 93498 3922 93554 3978
rect 93622 3922 93678 3978
rect 93250 -216 93306 -160
rect 93374 -216 93430 -160
rect 93498 -216 93554 -160
rect 93622 -216 93678 -160
rect 93250 -340 93306 -284
rect 93374 -340 93430 -284
rect 93498 -340 93554 -284
rect 93622 -340 93678 -284
rect 93250 -464 93306 -408
rect 93374 -464 93430 -408
rect 93498 -464 93554 -408
rect 93622 -464 93678 -408
rect 93250 -588 93306 -532
rect 93374 -588 93430 -532
rect 93498 -588 93554 -532
rect 93622 -588 93678 -532
rect 96970 64294 97026 64350
rect 97094 64294 97150 64350
rect 97218 64294 97274 64350
rect 97342 64294 97398 64350
rect 96970 64170 97026 64226
rect 97094 64170 97150 64226
rect 97218 64170 97274 64226
rect 97342 64170 97398 64226
rect 96970 64046 97026 64102
rect 97094 64046 97150 64102
rect 97218 64046 97274 64102
rect 97342 64046 97398 64102
rect 96970 63922 97026 63978
rect 97094 63922 97150 63978
rect 97218 63922 97274 63978
rect 97342 63922 97398 63978
rect 96970 46294 97026 46350
rect 97094 46294 97150 46350
rect 97218 46294 97274 46350
rect 97342 46294 97398 46350
rect 96970 46170 97026 46226
rect 97094 46170 97150 46226
rect 97218 46170 97274 46226
rect 97342 46170 97398 46226
rect 96970 46046 97026 46102
rect 97094 46046 97150 46102
rect 97218 46046 97274 46102
rect 97342 46046 97398 46102
rect 96970 45922 97026 45978
rect 97094 45922 97150 45978
rect 97218 45922 97274 45978
rect 97342 45922 97398 45978
rect 96970 28294 97026 28350
rect 97094 28294 97150 28350
rect 97218 28294 97274 28350
rect 97342 28294 97398 28350
rect 96970 28170 97026 28226
rect 97094 28170 97150 28226
rect 97218 28170 97274 28226
rect 97342 28170 97398 28226
rect 96970 28046 97026 28102
rect 97094 28046 97150 28102
rect 97218 28046 97274 28102
rect 97342 28046 97398 28102
rect 96970 27922 97026 27978
rect 97094 27922 97150 27978
rect 97218 27922 97274 27978
rect 97342 27922 97398 27978
rect 96970 10294 97026 10350
rect 97094 10294 97150 10350
rect 97218 10294 97274 10350
rect 97342 10294 97398 10350
rect 96970 10170 97026 10226
rect 97094 10170 97150 10226
rect 97218 10170 97274 10226
rect 97342 10170 97398 10226
rect 96970 10046 97026 10102
rect 97094 10046 97150 10102
rect 97218 10046 97274 10102
rect 97342 10046 97398 10102
rect 96970 9922 97026 9978
rect 97094 9922 97150 9978
rect 97218 9922 97274 9978
rect 97342 9922 97398 9978
rect 96970 -1176 97026 -1120
rect 97094 -1176 97150 -1120
rect 97218 -1176 97274 -1120
rect 97342 -1176 97398 -1120
rect 96970 -1300 97026 -1244
rect 97094 -1300 97150 -1244
rect 97218 -1300 97274 -1244
rect 97342 -1300 97398 -1244
rect 96970 -1424 97026 -1368
rect 97094 -1424 97150 -1368
rect 97218 -1424 97274 -1368
rect 97342 -1424 97398 -1368
rect 96970 -1548 97026 -1492
rect 97094 -1548 97150 -1492
rect 97218 -1548 97274 -1492
rect 97342 -1548 97398 -1492
rect 111250 76294 111306 76350
rect 111374 76294 111430 76350
rect 111498 76294 111554 76350
rect 111622 76294 111678 76350
rect 111250 76170 111306 76226
rect 111374 76170 111430 76226
rect 111498 76170 111554 76226
rect 111622 76170 111678 76226
rect 111250 76046 111306 76102
rect 111374 76046 111430 76102
rect 111498 76046 111554 76102
rect 111622 76046 111678 76102
rect 111250 75922 111306 75978
rect 111374 75922 111430 75978
rect 111498 75922 111554 75978
rect 111622 75922 111678 75978
rect 111250 58294 111306 58350
rect 111374 58294 111430 58350
rect 111498 58294 111554 58350
rect 111622 58294 111678 58350
rect 111250 58170 111306 58226
rect 111374 58170 111430 58226
rect 111498 58170 111554 58226
rect 111622 58170 111678 58226
rect 111250 58046 111306 58102
rect 111374 58046 111430 58102
rect 111498 58046 111554 58102
rect 111622 58046 111678 58102
rect 111250 57922 111306 57978
rect 111374 57922 111430 57978
rect 111498 57922 111554 57978
rect 111622 57922 111678 57978
rect 111250 40294 111306 40350
rect 111374 40294 111430 40350
rect 111498 40294 111554 40350
rect 111622 40294 111678 40350
rect 111250 40170 111306 40226
rect 111374 40170 111430 40226
rect 111498 40170 111554 40226
rect 111622 40170 111678 40226
rect 111250 40046 111306 40102
rect 111374 40046 111430 40102
rect 111498 40046 111554 40102
rect 111622 40046 111678 40102
rect 111250 39922 111306 39978
rect 111374 39922 111430 39978
rect 111498 39922 111554 39978
rect 111622 39922 111678 39978
rect 111250 22294 111306 22350
rect 111374 22294 111430 22350
rect 111498 22294 111554 22350
rect 111622 22294 111678 22350
rect 111250 22170 111306 22226
rect 111374 22170 111430 22226
rect 111498 22170 111554 22226
rect 111622 22170 111678 22226
rect 111250 22046 111306 22102
rect 111374 22046 111430 22102
rect 111498 22046 111554 22102
rect 111622 22046 111678 22102
rect 111250 21922 111306 21978
rect 111374 21922 111430 21978
rect 111498 21922 111554 21978
rect 111622 21922 111678 21978
rect 111250 4294 111306 4350
rect 111374 4294 111430 4350
rect 111498 4294 111554 4350
rect 111622 4294 111678 4350
rect 111250 4170 111306 4226
rect 111374 4170 111430 4226
rect 111498 4170 111554 4226
rect 111622 4170 111678 4226
rect 111250 4046 111306 4102
rect 111374 4046 111430 4102
rect 111498 4046 111554 4102
rect 111622 4046 111678 4102
rect 111250 3922 111306 3978
rect 111374 3922 111430 3978
rect 111498 3922 111554 3978
rect 111622 3922 111678 3978
rect 111250 -216 111306 -160
rect 111374 -216 111430 -160
rect 111498 -216 111554 -160
rect 111622 -216 111678 -160
rect 111250 -340 111306 -284
rect 111374 -340 111430 -284
rect 111498 -340 111554 -284
rect 111622 -340 111678 -284
rect 111250 -464 111306 -408
rect 111374 -464 111430 -408
rect 111498 -464 111554 -408
rect 111622 -464 111678 -408
rect 111250 -588 111306 -532
rect 111374 -588 111430 -532
rect 111498 -588 111554 -532
rect 111622 -588 111678 -532
rect 114970 64294 115026 64350
rect 115094 64294 115150 64350
rect 115218 64294 115274 64350
rect 115342 64294 115398 64350
rect 114970 64170 115026 64226
rect 115094 64170 115150 64226
rect 115218 64170 115274 64226
rect 115342 64170 115398 64226
rect 114970 64046 115026 64102
rect 115094 64046 115150 64102
rect 115218 64046 115274 64102
rect 115342 64046 115398 64102
rect 114970 63922 115026 63978
rect 115094 63922 115150 63978
rect 115218 63922 115274 63978
rect 115342 63922 115398 63978
rect 114970 46294 115026 46350
rect 115094 46294 115150 46350
rect 115218 46294 115274 46350
rect 115342 46294 115398 46350
rect 114970 46170 115026 46226
rect 115094 46170 115150 46226
rect 115218 46170 115274 46226
rect 115342 46170 115398 46226
rect 114970 46046 115026 46102
rect 115094 46046 115150 46102
rect 115218 46046 115274 46102
rect 115342 46046 115398 46102
rect 114970 45922 115026 45978
rect 115094 45922 115150 45978
rect 115218 45922 115274 45978
rect 115342 45922 115398 45978
rect 114970 28294 115026 28350
rect 115094 28294 115150 28350
rect 115218 28294 115274 28350
rect 115342 28294 115398 28350
rect 114970 28170 115026 28226
rect 115094 28170 115150 28226
rect 115218 28170 115274 28226
rect 115342 28170 115398 28226
rect 114970 28046 115026 28102
rect 115094 28046 115150 28102
rect 115218 28046 115274 28102
rect 115342 28046 115398 28102
rect 114970 27922 115026 27978
rect 115094 27922 115150 27978
rect 115218 27922 115274 27978
rect 115342 27922 115398 27978
rect 114970 10294 115026 10350
rect 115094 10294 115150 10350
rect 115218 10294 115274 10350
rect 115342 10294 115398 10350
rect 114970 10170 115026 10226
rect 115094 10170 115150 10226
rect 115218 10170 115274 10226
rect 115342 10170 115398 10226
rect 114970 10046 115026 10102
rect 115094 10046 115150 10102
rect 115218 10046 115274 10102
rect 115342 10046 115398 10102
rect 114970 9922 115026 9978
rect 115094 9922 115150 9978
rect 115218 9922 115274 9978
rect 115342 9922 115398 9978
rect 114970 -1176 115026 -1120
rect 115094 -1176 115150 -1120
rect 115218 -1176 115274 -1120
rect 115342 -1176 115398 -1120
rect 114970 -1300 115026 -1244
rect 115094 -1300 115150 -1244
rect 115218 -1300 115274 -1244
rect 115342 -1300 115398 -1244
rect 114970 -1424 115026 -1368
rect 115094 -1424 115150 -1368
rect 115218 -1424 115274 -1368
rect 115342 -1424 115398 -1368
rect 114970 -1548 115026 -1492
rect 115094 -1548 115150 -1492
rect 115218 -1548 115274 -1492
rect 115342 -1548 115398 -1492
rect 129250 76294 129306 76350
rect 129374 76294 129430 76350
rect 129498 76294 129554 76350
rect 129622 76294 129678 76350
rect 129250 76170 129306 76226
rect 129374 76170 129430 76226
rect 129498 76170 129554 76226
rect 129622 76170 129678 76226
rect 129250 76046 129306 76102
rect 129374 76046 129430 76102
rect 129498 76046 129554 76102
rect 129622 76046 129678 76102
rect 129250 75922 129306 75978
rect 129374 75922 129430 75978
rect 129498 75922 129554 75978
rect 129622 75922 129678 75978
rect 129250 58294 129306 58350
rect 129374 58294 129430 58350
rect 129498 58294 129554 58350
rect 129622 58294 129678 58350
rect 129250 58170 129306 58226
rect 129374 58170 129430 58226
rect 129498 58170 129554 58226
rect 129622 58170 129678 58226
rect 129250 58046 129306 58102
rect 129374 58046 129430 58102
rect 129498 58046 129554 58102
rect 129622 58046 129678 58102
rect 129250 57922 129306 57978
rect 129374 57922 129430 57978
rect 129498 57922 129554 57978
rect 129622 57922 129678 57978
rect 129250 40294 129306 40350
rect 129374 40294 129430 40350
rect 129498 40294 129554 40350
rect 129622 40294 129678 40350
rect 129250 40170 129306 40226
rect 129374 40170 129430 40226
rect 129498 40170 129554 40226
rect 129622 40170 129678 40226
rect 129250 40046 129306 40102
rect 129374 40046 129430 40102
rect 129498 40046 129554 40102
rect 129622 40046 129678 40102
rect 129250 39922 129306 39978
rect 129374 39922 129430 39978
rect 129498 39922 129554 39978
rect 129622 39922 129678 39978
rect 129250 22294 129306 22350
rect 129374 22294 129430 22350
rect 129498 22294 129554 22350
rect 129622 22294 129678 22350
rect 129250 22170 129306 22226
rect 129374 22170 129430 22226
rect 129498 22170 129554 22226
rect 129622 22170 129678 22226
rect 129250 22046 129306 22102
rect 129374 22046 129430 22102
rect 129498 22046 129554 22102
rect 129622 22046 129678 22102
rect 129250 21922 129306 21978
rect 129374 21922 129430 21978
rect 129498 21922 129554 21978
rect 129622 21922 129678 21978
rect 129250 4294 129306 4350
rect 129374 4294 129430 4350
rect 129498 4294 129554 4350
rect 129622 4294 129678 4350
rect 129250 4170 129306 4226
rect 129374 4170 129430 4226
rect 129498 4170 129554 4226
rect 129622 4170 129678 4226
rect 129250 4046 129306 4102
rect 129374 4046 129430 4102
rect 129498 4046 129554 4102
rect 129622 4046 129678 4102
rect 129250 3922 129306 3978
rect 129374 3922 129430 3978
rect 129498 3922 129554 3978
rect 129622 3922 129678 3978
rect 129250 -216 129306 -160
rect 129374 -216 129430 -160
rect 129498 -216 129554 -160
rect 129622 -216 129678 -160
rect 129250 -340 129306 -284
rect 129374 -340 129430 -284
rect 129498 -340 129554 -284
rect 129622 -340 129678 -284
rect 129250 -464 129306 -408
rect 129374 -464 129430 -408
rect 129498 -464 129554 -408
rect 129622 -464 129678 -408
rect 129250 -588 129306 -532
rect 129374 -588 129430 -532
rect 129498 -588 129554 -532
rect 129622 -588 129678 -532
rect 132970 64294 133026 64350
rect 133094 64294 133150 64350
rect 133218 64294 133274 64350
rect 133342 64294 133398 64350
rect 132970 64170 133026 64226
rect 133094 64170 133150 64226
rect 133218 64170 133274 64226
rect 133342 64170 133398 64226
rect 132970 64046 133026 64102
rect 133094 64046 133150 64102
rect 133218 64046 133274 64102
rect 133342 64046 133398 64102
rect 132970 63922 133026 63978
rect 133094 63922 133150 63978
rect 133218 63922 133274 63978
rect 133342 63922 133398 63978
rect 132970 46294 133026 46350
rect 133094 46294 133150 46350
rect 133218 46294 133274 46350
rect 133342 46294 133398 46350
rect 132970 46170 133026 46226
rect 133094 46170 133150 46226
rect 133218 46170 133274 46226
rect 133342 46170 133398 46226
rect 132970 46046 133026 46102
rect 133094 46046 133150 46102
rect 133218 46046 133274 46102
rect 133342 46046 133398 46102
rect 132970 45922 133026 45978
rect 133094 45922 133150 45978
rect 133218 45922 133274 45978
rect 133342 45922 133398 45978
rect 132970 28294 133026 28350
rect 133094 28294 133150 28350
rect 133218 28294 133274 28350
rect 133342 28294 133398 28350
rect 132970 28170 133026 28226
rect 133094 28170 133150 28226
rect 133218 28170 133274 28226
rect 133342 28170 133398 28226
rect 132970 28046 133026 28102
rect 133094 28046 133150 28102
rect 133218 28046 133274 28102
rect 133342 28046 133398 28102
rect 132970 27922 133026 27978
rect 133094 27922 133150 27978
rect 133218 27922 133274 27978
rect 133342 27922 133398 27978
rect 132970 10294 133026 10350
rect 133094 10294 133150 10350
rect 133218 10294 133274 10350
rect 133342 10294 133398 10350
rect 132970 10170 133026 10226
rect 133094 10170 133150 10226
rect 133218 10170 133274 10226
rect 133342 10170 133398 10226
rect 132970 10046 133026 10102
rect 133094 10046 133150 10102
rect 133218 10046 133274 10102
rect 133342 10046 133398 10102
rect 132970 9922 133026 9978
rect 133094 9922 133150 9978
rect 133218 9922 133274 9978
rect 133342 9922 133398 9978
rect 132970 -1176 133026 -1120
rect 133094 -1176 133150 -1120
rect 133218 -1176 133274 -1120
rect 133342 -1176 133398 -1120
rect 132970 -1300 133026 -1244
rect 133094 -1300 133150 -1244
rect 133218 -1300 133274 -1244
rect 133342 -1300 133398 -1244
rect 132970 -1424 133026 -1368
rect 133094 -1424 133150 -1368
rect 133218 -1424 133274 -1368
rect 133342 -1424 133398 -1368
rect 132970 -1548 133026 -1492
rect 133094 -1548 133150 -1492
rect 133218 -1548 133274 -1492
rect 133342 -1548 133398 -1492
rect 147250 76294 147306 76350
rect 147374 76294 147430 76350
rect 147498 76294 147554 76350
rect 147622 76294 147678 76350
rect 147250 76170 147306 76226
rect 147374 76170 147430 76226
rect 147498 76170 147554 76226
rect 147622 76170 147678 76226
rect 147250 76046 147306 76102
rect 147374 76046 147430 76102
rect 147498 76046 147554 76102
rect 147622 76046 147678 76102
rect 147250 75922 147306 75978
rect 147374 75922 147430 75978
rect 147498 75922 147554 75978
rect 147622 75922 147678 75978
rect 147250 58294 147306 58350
rect 147374 58294 147430 58350
rect 147498 58294 147554 58350
rect 147622 58294 147678 58350
rect 147250 58170 147306 58226
rect 147374 58170 147430 58226
rect 147498 58170 147554 58226
rect 147622 58170 147678 58226
rect 147250 58046 147306 58102
rect 147374 58046 147430 58102
rect 147498 58046 147554 58102
rect 147622 58046 147678 58102
rect 147250 57922 147306 57978
rect 147374 57922 147430 57978
rect 147498 57922 147554 57978
rect 147622 57922 147678 57978
rect 147250 40294 147306 40350
rect 147374 40294 147430 40350
rect 147498 40294 147554 40350
rect 147622 40294 147678 40350
rect 147250 40170 147306 40226
rect 147374 40170 147430 40226
rect 147498 40170 147554 40226
rect 147622 40170 147678 40226
rect 147250 40046 147306 40102
rect 147374 40046 147430 40102
rect 147498 40046 147554 40102
rect 147622 40046 147678 40102
rect 147250 39922 147306 39978
rect 147374 39922 147430 39978
rect 147498 39922 147554 39978
rect 147622 39922 147678 39978
rect 147250 22294 147306 22350
rect 147374 22294 147430 22350
rect 147498 22294 147554 22350
rect 147622 22294 147678 22350
rect 147250 22170 147306 22226
rect 147374 22170 147430 22226
rect 147498 22170 147554 22226
rect 147622 22170 147678 22226
rect 147250 22046 147306 22102
rect 147374 22046 147430 22102
rect 147498 22046 147554 22102
rect 147622 22046 147678 22102
rect 147250 21922 147306 21978
rect 147374 21922 147430 21978
rect 147498 21922 147554 21978
rect 147622 21922 147678 21978
rect 147250 4294 147306 4350
rect 147374 4294 147430 4350
rect 147498 4294 147554 4350
rect 147622 4294 147678 4350
rect 147250 4170 147306 4226
rect 147374 4170 147430 4226
rect 147498 4170 147554 4226
rect 147622 4170 147678 4226
rect 147250 4046 147306 4102
rect 147374 4046 147430 4102
rect 147498 4046 147554 4102
rect 147622 4046 147678 4102
rect 147250 3922 147306 3978
rect 147374 3922 147430 3978
rect 147498 3922 147554 3978
rect 147622 3922 147678 3978
rect 147250 -216 147306 -160
rect 147374 -216 147430 -160
rect 147498 -216 147554 -160
rect 147622 -216 147678 -160
rect 147250 -340 147306 -284
rect 147374 -340 147430 -284
rect 147498 -340 147554 -284
rect 147622 -340 147678 -284
rect 147250 -464 147306 -408
rect 147374 -464 147430 -408
rect 147498 -464 147554 -408
rect 147622 -464 147678 -408
rect 147250 -588 147306 -532
rect 147374 -588 147430 -532
rect 147498 -588 147554 -532
rect 147622 -588 147678 -532
rect 150970 64294 151026 64350
rect 151094 64294 151150 64350
rect 151218 64294 151274 64350
rect 151342 64294 151398 64350
rect 150970 64170 151026 64226
rect 151094 64170 151150 64226
rect 151218 64170 151274 64226
rect 151342 64170 151398 64226
rect 150970 64046 151026 64102
rect 151094 64046 151150 64102
rect 151218 64046 151274 64102
rect 151342 64046 151398 64102
rect 150970 63922 151026 63978
rect 151094 63922 151150 63978
rect 151218 63922 151274 63978
rect 151342 63922 151398 63978
rect 150970 46294 151026 46350
rect 151094 46294 151150 46350
rect 151218 46294 151274 46350
rect 151342 46294 151398 46350
rect 150970 46170 151026 46226
rect 151094 46170 151150 46226
rect 151218 46170 151274 46226
rect 151342 46170 151398 46226
rect 150970 46046 151026 46102
rect 151094 46046 151150 46102
rect 151218 46046 151274 46102
rect 151342 46046 151398 46102
rect 150970 45922 151026 45978
rect 151094 45922 151150 45978
rect 151218 45922 151274 45978
rect 151342 45922 151398 45978
rect 150970 28294 151026 28350
rect 151094 28294 151150 28350
rect 151218 28294 151274 28350
rect 151342 28294 151398 28350
rect 150970 28170 151026 28226
rect 151094 28170 151150 28226
rect 151218 28170 151274 28226
rect 151342 28170 151398 28226
rect 150970 28046 151026 28102
rect 151094 28046 151150 28102
rect 151218 28046 151274 28102
rect 151342 28046 151398 28102
rect 150970 27922 151026 27978
rect 151094 27922 151150 27978
rect 151218 27922 151274 27978
rect 151342 27922 151398 27978
rect 150970 10294 151026 10350
rect 151094 10294 151150 10350
rect 151218 10294 151274 10350
rect 151342 10294 151398 10350
rect 150970 10170 151026 10226
rect 151094 10170 151150 10226
rect 151218 10170 151274 10226
rect 151342 10170 151398 10226
rect 150970 10046 151026 10102
rect 151094 10046 151150 10102
rect 151218 10046 151274 10102
rect 151342 10046 151398 10102
rect 150970 9922 151026 9978
rect 151094 9922 151150 9978
rect 151218 9922 151274 9978
rect 151342 9922 151398 9978
rect 150970 -1176 151026 -1120
rect 151094 -1176 151150 -1120
rect 151218 -1176 151274 -1120
rect 151342 -1176 151398 -1120
rect 150970 -1300 151026 -1244
rect 151094 -1300 151150 -1244
rect 151218 -1300 151274 -1244
rect 151342 -1300 151398 -1244
rect 150970 -1424 151026 -1368
rect 151094 -1424 151150 -1368
rect 151218 -1424 151274 -1368
rect 151342 -1424 151398 -1368
rect 150970 -1548 151026 -1492
rect 151094 -1548 151150 -1492
rect 151218 -1548 151274 -1492
rect 151342 -1548 151398 -1492
rect 165250 76294 165306 76350
rect 165374 76294 165430 76350
rect 165498 76294 165554 76350
rect 165622 76294 165678 76350
rect 165250 76170 165306 76226
rect 165374 76170 165430 76226
rect 165498 76170 165554 76226
rect 165622 76170 165678 76226
rect 165250 76046 165306 76102
rect 165374 76046 165430 76102
rect 165498 76046 165554 76102
rect 165622 76046 165678 76102
rect 165250 75922 165306 75978
rect 165374 75922 165430 75978
rect 165498 75922 165554 75978
rect 165622 75922 165678 75978
rect 165250 58294 165306 58350
rect 165374 58294 165430 58350
rect 165498 58294 165554 58350
rect 165622 58294 165678 58350
rect 165250 58170 165306 58226
rect 165374 58170 165430 58226
rect 165498 58170 165554 58226
rect 165622 58170 165678 58226
rect 165250 58046 165306 58102
rect 165374 58046 165430 58102
rect 165498 58046 165554 58102
rect 165622 58046 165678 58102
rect 165250 57922 165306 57978
rect 165374 57922 165430 57978
rect 165498 57922 165554 57978
rect 165622 57922 165678 57978
rect 165250 40294 165306 40350
rect 165374 40294 165430 40350
rect 165498 40294 165554 40350
rect 165622 40294 165678 40350
rect 165250 40170 165306 40226
rect 165374 40170 165430 40226
rect 165498 40170 165554 40226
rect 165622 40170 165678 40226
rect 165250 40046 165306 40102
rect 165374 40046 165430 40102
rect 165498 40046 165554 40102
rect 165622 40046 165678 40102
rect 165250 39922 165306 39978
rect 165374 39922 165430 39978
rect 165498 39922 165554 39978
rect 165622 39922 165678 39978
rect 165250 22294 165306 22350
rect 165374 22294 165430 22350
rect 165498 22294 165554 22350
rect 165622 22294 165678 22350
rect 165250 22170 165306 22226
rect 165374 22170 165430 22226
rect 165498 22170 165554 22226
rect 165622 22170 165678 22226
rect 165250 22046 165306 22102
rect 165374 22046 165430 22102
rect 165498 22046 165554 22102
rect 165622 22046 165678 22102
rect 165250 21922 165306 21978
rect 165374 21922 165430 21978
rect 165498 21922 165554 21978
rect 165622 21922 165678 21978
rect 165250 4294 165306 4350
rect 165374 4294 165430 4350
rect 165498 4294 165554 4350
rect 165622 4294 165678 4350
rect 165250 4170 165306 4226
rect 165374 4170 165430 4226
rect 165498 4170 165554 4226
rect 165622 4170 165678 4226
rect 165250 4046 165306 4102
rect 165374 4046 165430 4102
rect 165498 4046 165554 4102
rect 165622 4046 165678 4102
rect 165250 3922 165306 3978
rect 165374 3922 165430 3978
rect 165498 3922 165554 3978
rect 165622 3922 165678 3978
rect 165250 -216 165306 -160
rect 165374 -216 165430 -160
rect 165498 -216 165554 -160
rect 165622 -216 165678 -160
rect 165250 -340 165306 -284
rect 165374 -340 165430 -284
rect 165498 -340 165554 -284
rect 165622 -340 165678 -284
rect 165250 -464 165306 -408
rect 165374 -464 165430 -408
rect 165498 -464 165554 -408
rect 165622 -464 165678 -408
rect 165250 -588 165306 -532
rect 165374 -588 165430 -532
rect 165498 -588 165554 -532
rect 165622 -588 165678 -532
rect 168970 64294 169026 64350
rect 169094 64294 169150 64350
rect 169218 64294 169274 64350
rect 169342 64294 169398 64350
rect 168970 64170 169026 64226
rect 169094 64170 169150 64226
rect 169218 64170 169274 64226
rect 169342 64170 169398 64226
rect 168970 64046 169026 64102
rect 169094 64046 169150 64102
rect 169218 64046 169274 64102
rect 169342 64046 169398 64102
rect 168970 63922 169026 63978
rect 169094 63922 169150 63978
rect 169218 63922 169274 63978
rect 169342 63922 169398 63978
rect 168970 46294 169026 46350
rect 169094 46294 169150 46350
rect 169218 46294 169274 46350
rect 169342 46294 169398 46350
rect 168970 46170 169026 46226
rect 169094 46170 169150 46226
rect 169218 46170 169274 46226
rect 169342 46170 169398 46226
rect 168970 46046 169026 46102
rect 169094 46046 169150 46102
rect 169218 46046 169274 46102
rect 169342 46046 169398 46102
rect 168970 45922 169026 45978
rect 169094 45922 169150 45978
rect 169218 45922 169274 45978
rect 169342 45922 169398 45978
rect 168970 28294 169026 28350
rect 169094 28294 169150 28350
rect 169218 28294 169274 28350
rect 169342 28294 169398 28350
rect 168970 28170 169026 28226
rect 169094 28170 169150 28226
rect 169218 28170 169274 28226
rect 169342 28170 169398 28226
rect 168970 28046 169026 28102
rect 169094 28046 169150 28102
rect 169218 28046 169274 28102
rect 169342 28046 169398 28102
rect 168970 27922 169026 27978
rect 169094 27922 169150 27978
rect 169218 27922 169274 27978
rect 169342 27922 169398 27978
rect 168970 10294 169026 10350
rect 169094 10294 169150 10350
rect 169218 10294 169274 10350
rect 169342 10294 169398 10350
rect 168970 10170 169026 10226
rect 169094 10170 169150 10226
rect 169218 10170 169274 10226
rect 169342 10170 169398 10226
rect 168970 10046 169026 10102
rect 169094 10046 169150 10102
rect 169218 10046 169274 10102
rect 169342 10046 169398 10102
rect 168970 9922 169026 9978
rect 169094 9922 169150 9978
rect 169218 9922 169274 9978
rect 169342 9922 169398 9978
rect 168970 -1176 169026 -1120
rect 169094 -1176 169150 -1120
rect 169218 -1176 169274 -1120
rect 169342 -1176 169398 -1120
rect 168970 -1300 169026 -1244
rect 169094 -1300 169150 -1244
rect 169218 -1300 169274 -1244
rect 169342 -1300 169398 -1244
rect 168970 -1424 169026 -1368
rect 169094 -1424 169150 -1368
rect 169218 -1424 169274 -1368
rect 169342 -1424 169398 -1368
rect 168970 -1548 169026 -1492
rect 169094 -1548 169150 -1492
rect 169218 -1548 169274 -1492
rect 169342 -1548 169398 -1492
rect 183250 76294 183306 76350
rect 183374 76294 183430 76350
rect 183498 76294 183554 76350
rect 183622 76294 183678 76350
rect 183250 76170 183306 76226
rect 183374 76170 183430 76226
rect 183498 76170 183554 76226
rect 183622 76170 183678 76226
rect 183250 76046 183306 76102
rect 183374 76046 183430 76102
rect 183498 76046 183554 76102
rect 183622 76046 183678 76102
rect 183250 75922 183306 75978
rect 183374 75922 183430 75978
rect 183498 75922 183554 75978
rect 183622 75922 183678 75978
rect 183250 58294 183306 58350
rect 183374 58294 183430 58350
rect 183498 58294 183554 58350
rect 183622 58294 183678 58350
rect 183250 58170 183306 58226
rect 183374 58170 183430 58226
rect 183498 58170 183554 58226
rect 183622 58170 183678 58226
rect 183250 58046 183306 58102
rect 183374 58046 183430 58102
rect 183498 58046 183554 58102
rect 183622 58046 183678 58102
rect 183250 57922 183306 57978
rect 183374 57922 183430 57978
rect 183498 57922 183554 57978
rect 183622 57922 183678 57978
rect 183250 40294 183306 40350
rect 183374 40294 183430 40350
rect 183498 40294 183554 40350
rect 183622 40294 183678 40350
rect 183250 40170 183306 40226
rect 183374 40170 183430 40226
rect 183498 40170 183554 40226
rect 183622 40170 183678 40226
rect 183250 40046 183306 40102
rect 183374 40046 183430 40102
rect 183498 40046 183554 40102
rect 183622 40046 183678 40102
rect 183250 39922 183306 39978
rect 183374 39922 183430 39978
rect 183498 39922 183554 39978
rect 183622 39922 183678 39978
rect 183250 22294 183306 22350
rect 183374 22294 183430 22350
rect 183498 22294 183554 22350
rect 183622 22294 183678 22350
rect 183250 22170 183306 22226
rect 183374 22170 183430 22226
rect 183498 22170 183554 22226
rect 183622 22170 183678 22226
rect 183250 22046 183306 22102
rect 183374 22046 183430 22102
rect 183498 22046 183554 22102
rect 183622 22046 183678 22102
rect 183250 21922 183306 21978
rect 183374 21922 183430 21978
rect 183498 21922 183554 21978
rect 183622 21922 183678 21978
rect 183250 4294 183306 4350
rect 183374 4294 183430 4350
rect 183498 4294 183554 4350
rect 183622 4294 183678 4350
rect 183250 4170 183306 4226
rect 183374 4170 183430 4226
rect 183498 4170 183554 4226
rect 183622 4170 183678 4226
rect 183250 4046 183306 4102
rect 183374 4046 183430 4102
rect 183498 4046 183554 4102
rect 183622 4046 183678 4102
rect 183250 3922 183306 3978
rect 183374 3922 183430 3978
rect 183498 3922 183554 3978
rect 183622 3922 183678 3978
rect 183250 -216 183306 -160
rect 183374 -216 183430 -160
rect 183498 -216 183554 -160
rect 183622 -216 183678 -160
rect 183250 -340 183306 -284
rect 183374 -340 183430 -284
rect 183498 -340 183554 -284
rect 183622 -340 183678 -284
rect 183250 -464 183306 -408
rect 183374 -464 183430 -408
rect 183498 -464 183554 -408
rect 183622 -464 183678 -408
rect 183250 -588 183306 -532
rect 183374 -588 183430 -532
rect 183498 -588 183554 -532
rect 183622 -588 183678 -532
rect 186970 154294 187026 154350
rect 187094 154294 187150 154350
rect 187218 154294 187274 154350
rect 187342 154294 187398 154350
rect 186970 154170 187026 154226
rect 187094 154170 187150 154226
rect 187218 154170 187274 154226
rect 187342 154170 187398 154226
rect 186970 154046 187026 154102
rect 187094 154046 187150 154102
rect 187218 154046 187274 154102
rect 187342 154046 187398 154102
rect 186970 153922 187026 153978
rect 187094 153922 187150 153978
rect 187218 153922 187274 153978
rect 187342 153922 187398 153978
rect 186970 136294 187026 136350
rect 187094 136294 187150 136350
rect 187218 136294 187274 136350
rect 187342 136294 187398 136350
rect 186970 136170 187026 136226
rect 187094 136170 187150 136226
rect 187218 136170 187274 136226
rect 187342 136170 187398 136226
rect 186970 136046 187026 136102
rect 187094 136046 187150 136102
rect 187218 136046 187274 136102
rect 187342 136046 187398 136102
rect 186970 135922 187026 135978
rect 187094 135922 187150 135978
rect 187218 135922 187274 135978
rect 187342 135922 187398 135978
rect 186970 118294 187026 118350
rect 187094 118294 187150 118350
rect 187218 118294 187274 118350
rect 187342 118294 187398 118350
rect 186970 118170 187026 118226
rect 187094 118170 187150 118226
rect 187218 118170 187274 118226
rect 187342 118170 187398 118226
rect 186970 118046 187026 118102
rect 187094 118046 187150 118102
rect 187218 118046 187274 118102
rect 187342 118046 187398 118102
rect 186970 117922 187026 117978
rect 187094 117922 187150 117978
rect 187218 117922 187274 117978
rect 187342 117922 187398 117978
rect 186970 100294 187026 100350
rect 187094 100294 187150 100350
rect 187218 100294 187274 100350
rect 187342 100294 187398 100350
rect 186970 100170 187026 100226
rect 187094 100170 187150 100226
rect 187218 100170 187274 100226
rect 187342 100170 187398 100226
rect 186970 100046 187026 100102
rect 187094 100046 187150 100102
rect 187218 100046 187274 100102
rect 187342 100046 187398 100102
rect 186970 99922 187026 99978
rect 187094 99922 187150 99978
rect 187218 99922 187274 99978
rect 187342 99922 187398 99978
rect 186970 82294 187026 82350
rect 187094 82294 187150 82350
rect 187218 82294 187274 82350
rect 187342 82294 187398 82350
rect 186970 82170 187026 82226
rect 187094 82170 187150 82226
rect 187218 82170 187274 82226
rect 187342 82170 187398 82226
rect 186970 82046 187026 82102
rect 187094 82046 187150 82102
rect 187218 82046 187274 82102
rect 187342 82046 187398 82102
rect 186970 81922 187026 81978
rect 187094 81922 187150 81978
rect 187218 81922 187274 81978
rect 187342 81922 187398 81978
rect 186970 64294 187026 64350
rect 187094 64294 187150 64350
rect 187218 64294 187274 64350
rect 187342 64294 187398 64350
rect 186970 64170 187026 64226
rect 187094 64170 187150 64226
rect 187218 64170 187274 64226
rect 187342 64170 187398 64226
rect 186970 64046 187026 64102
rect 187094 64046 187150 64102
rect 187218 64046 187274 64102
rect 187342 64046 187398 64102
rect 186970 63922 187026 63978
rect 187094 63922 187150 63978
rect 187218 63922 187274 63978
rect 187342 63922 187398 63978
rect 186970 46294 187026 46350
rect 187094 46294 187150 46350
rect 187218 46294 187274 46350
rect 187342 46294 187398 46350
rect 186970 46170 187026 46226
rect 187094 46170 187150 46226
rect 187218 46170 187274 46226
rect 187342 46170 187398 46226
rect 186970 46046 187026 46102
rect 187094 46046 187150 46102
rect 187218 46046 187274 46102
rect 187342 46046 187398 46102
rect 186970 45922 187026 45978
rect 187094 45922 187150 45978
rect 187218 45922 187274 45978
rect 187342 45922 187398 45978
rect 186970 28294 187026 28350
rect 187094 28294 187150 28350
rect 187218 28294 187274 28350
rect 187342 28294 187398 28350
rect 186970 28170 187026 28226
rect 187094 28170 187150 28226
rect 187218 28170 187274 28226
rect 187342 28170 187398 28226
rect 186970 28046 187026 28102
rect 187094 28046 187150 28102
rect 187218 28046 187274 28102
rect 187342 28046 187398 28102
rect 186970 27922 187026 27978
rect 187094 27922 187150 27978
rect 187218 27922 187274 27978
rect 187342 27922 187398 27978
rect 186970 10294 187026 10350
rect 187094 10294 187150 10350
rect 187218 10294 187274 10350
rect 187342 10294 187398 10350
rect 186970 10170 187026 10226
rect 187094 10170 187150 10226
rect 187218 10170 187274 10226
rect 187342 10170 187398 10226
rect 186970 10046 187026 10102
rect 187094 10046 187150 10102
rect 187218 10046 187274 10102
rect 187342 10046 187398 10102
rect 186970 9922 187026 9978
rect 187094 9922 187150 9978
rect 187218 9922 187274 9978
rect 187342 9922 187398 9978
rect 201250 580294 201306 580350
rect 201374 580294 201430 580350
rect 201498 580294 201554 580350
rect 201622 580294 201678 580350
rect 201250 580170 201306 580226
rect 201374 580170 201430 580226
rect 201498 580170 201554 580226
rect 201622 580170 201678 580226
rect 201250 580046 201306 580102
rect 201374 580046 201430 580102
rect 201498 580046 201554 580102
rect 201622 580046 201678 580102
rect 201250 579922 201306 579978
rect 201374 579922 201430 579978
rect 201498 579922 201554 579978
rect 201622 579922 201678 579978
rect 201250 562294 201306 562350
rect 201374 562294 201430 562350
rect 201498 562294 201554 562350
rect 201622 562294 201678 562350
rect 201250 562170 201306 562226
rect 201374 562170 201430 562226
rect 201498 562170 201554 562226
rect 201622 562170 201678 562226
rect 201250 562046 201306 562102
rect 201374 562046 201430 562102
rect 201498 562046 201554 562102
rect 201622 562046 201678 562102
rect 201250 561922 201306 561978
rect 201374 561922 201430 561978
rect 201498 561922 201554 561978
rect 201622 561922 201678 561978
rect 201250 544294 201306 544350
rect 201374 544294 201430 544350
rect 201498 544294 201554 544350
rect 201622 544294 201678 544350
rect 201250 544170 201306 544226
rect 201374 544170 201430 544226
rect 201498 544170 201554 544226
rect 201622 544170 201678 544226
rect 201250 544046 201306 544102
rect 201374 544046 201430 544102
rect 201498 544046 201554 544102
rect 201622 544046 201678 544102
rect 201250 543922 201306 543978
rect 201374 543922 201430 543978
rect 201498 543922 201554 543978
rect 201622 543922 201678 543978
rect 201250 526294 201306 526350
rect 201374 526294 201430 526350
rect 201498 526294 201554 526350
rect 201622 526294 201678 526350
rect 201250 526170 201306 526226
rect 201374 526170 201430 526226
rect 201498 526170 201554 526226
rect 201622 526170 201678 526226
rect 201250 526046 201306 526102
rect 201374 526046 201430 526102
rect 201498 526046 201554 526102
rect 201622 526046 201678 526102
rect 201250 525922 201306 525978
rect 201374 525922 201430 525978
rect 201498 525922 201554 525978
rect 201622 525922 201678 525978
rect 201250 508294 201306 508350
rect 201374 508294 201430 508350
rect 201498 508294 201554 508350
rect 201622 508294 201678 508350
rect 201250 508170 201306 508226
rect 201374 508170 201430 508226
rect 201498 508170 201554 508226
rect 201622 508170 201678 508226
rect 201250 508046 201306 508102
rect 201374 508046 201430 508102
rect 201498 508046 201554 508102
rect 201622 508046 201678 508102
rect 201250 507922 201306 507978
rect 201374 507922 201430 507978
rect 201498 507922 201554 507978
rect 201622 507922 201678 507978
rect 201250 490294 201306 490350
rect 201374 490294 201430 490350
rect 201498 490294 201554 490350
rect 201622 490294 201678 490350
rect 201250 490170 201306 490226
rect 201374 490170 201430 490226
rect 201498 490170 201554 490226
rect 201622 490170 201678 490226
rect 201250 490046 201306 490102
rect 201374 490046 201430 490102
rect 201498 490046 201554 490102
rect 201622 490046 201678 490102
rect 201250 489922 201306 489978
rect 201374 489922 201430 489978
rect 201498 489922 201554 489978
rect 201622 489922 201678 489978
rect 201250 472294 201306 472350
rect 201374 472294 201430 472350
rect 201498 472294 201554 472350
rect 201622 472294 201678 472350
rect 201250 472170 201306 472226
rect 201374 472170 201430 472226
rect 201498 472170 201554 472226
rect 201622 472170 201678 472226
rect 201250 472046 201306 472102
rect 201374 472046 201430 472102
rect 201498 472046 201554 472102
rect 201622 472046 201678 472102
rect 201250 471922 201306 471978
rect 201374 471922 201430 471978
rect 201498 471922 201554 471978
rect 201622 471922 201678 471978
rect 201250 454294 201306 454350
rect 201374 454294 201430 454350
rect 201498 454294 201554 454350
rect 201622 454294 201678 454350
rect 201250 454170 201306 454226
rect 201374 454170 201430 454226
rect 201498 454170 201554 454226
rect 201622 454170 201678 454226
rect 201250 454046 201306 454102
rect 201374 454046 201430 454102
rect 201498 454046 201554 454102
rect 201622 454046 201678 454102
rect 201250 453922 201306 453978
rect 201374 453922 201430 453978
rect 201498 453922 201554 453978
rect 201622 453922 201678 453978
rect 201250 436294 201306 436350
rect 201374 436294 201430 436350
rect 201498 436294 201554 436350
rect 201622 436294 201678 436350
rect 201250 436170 201306 436226
rect 201374 436170 201430 436226
rect 201498 436170 201554 436226
rect 201622 436170 201678 436226
rect 201250 436046 201306 436102
rect 201374 436046 201430 436102
rect 201498 436046 201554 436102
rect 201622 436046 201678 436102
rect 201250 435922 201306 435978
rect 201374 435922 201430 435978
rect 201498 435922 201554 435978
rect 201622 435922 201678 435978
rect 201250 418294 201306 418350
rect 201374 418294 201430 418350
rect 201498 418294 201554 418350
rect 201622 418294 201678 418350
rect 201250 418170 201306 418226
rect 201374 418170 201430 418226
rect 201498 418170 201554 418226
rect 201622 418170 201678 418226
rect 201250 418046 201306 418102
rect 201374 418046 201430 418102
rect 201498 418046 201554 418102
rect 201622 418046 201678 418102
rect 201250 417922 201306 417978
rect 201374 417922 201430 417978
rect 201498 417922 201554 417978
rect 201622 417922 201678 417978
rect 201250 400294 201306 400350
rect 201374 400294 201430 400350
rect 201498 400294 201554 400350
rect 201622 400294 201678 400350
rect 201250 400170 201306 400226
rect 201374 400170 201430 400226
rect 201498 400170 201554 400226
rect 201622 400170 201678 400226
rect 201250 400046 201306 400102
rect 201374 400046 201430 400102
rect 201498 400046 201554 400102
rect 201622 400046 201678 400102
rect 201250 399922 201306 399978
rect 201374 399922 201430 399978
rect 201498 399922 201554 399978
rect 201622 399922 201678 399978
rect 201250 382294 201306 382350
rect 201374 382294 201430 382350
rect 201498 382294 201554 382350
rect 201622 382294 201678 382350
rect 201250 382170 201306 382226
rect 201374 382170 201430 382226
rect 201498 382170 201554 382226
rect 201622 382170 201678 382226
rect 201250 382046 201306 382102
rect 201374 382046 201430 382102
rect 201498 382046 201554 382102
rect 201622 382046 201678 382102
rect 201250 381922 201306 381978
rect 201374 381922 201430 381978
rect 201498 381922 201554 381978
rect 201622 381922 201678 381978
rect 201250 364294 201306 364350
rect 201374 364294 201430 364350
rect 201498 364294 201554 364350
rect 201622 364294 201678 364350
rect 201250 364170 201306 364226
rect 201374 364170 201430 364226
rect 201498 364170 201554 364226
rect 201622 364170 201678 364226
rect 201250 364046 201306 364102
rect 201374 364046 201430 364102
rect 201498 364046 201554 364102
rect 201622 364046 201678 364102
rect 201250 363922 201306 363978
rect 201374 363922 201430 363978
rect 201498 363922 201554 363978
rect 201622 363922 201678 363978
rect 201250 346294 201306 346350
rect 201374 346294 201430 346350
rect 201498 346294 201554 346350
rect 201622 346294 201678 346350
rect 201250 346170 201306 346226
rect 201374 346170 201430 346226
rect 201498 346170 201554 346226
rect 201622 346170 201678 346226
rect 201250 346046 201306 346102
rect 201374 346046 201430 346102
rect 201498 346046 201554 346102
rect 201622 346046 201678 346102
rect 201250 345922 201306 345978
rect 201374 345922 201430 345978
rect 201498 345922 201554 345978
rect 201622 345922 201678 345978
rect 201250 328294 201306 328350
rect 201374 328294 201430 328350
rect 201498 328294 201554 328350
rect 201622 328294 201678 328350
rect 201250 328170 201306 328226
rect 201374 328170 201430 328226
rect 201498 328170 201554 328226
rect 201622 328170 201678 328226
rect 201250 328046 201306 328102
rect 201374 328046 201430 328102
rect 201498 328046 201554 328102
rect 201622 328046 201678 328102
rect 201250 327922 201306 327978
rect 201374 327922 201430 327978
rect 201498 327922 201554 327978
rect 201622 327922 201678 327978
rect 201250 310294 201306 310350
rect 201374 310294 201430 310350
rect 201498 310294 201554 310350
rect 201622 310294 201678 310350
rect 201250 310170 201306 310226
rect 201374 310170 201430 310226
rect 201498 310170 201554 310226
rect 201622 310170 201678 310226
rect 201250 310046 201306 310102
rect 201374 310046 201430 310102
rect 201498 310046 201554 310102
rect 201622 310046 201678 310102
rect 201250 309922 201306 309978
rect 201374 309922 201430 309978
rect 201498 309922 201554 309978
rect 201622 309922 201678 309978
rect 201250 292294 201306 292350
rect 201374 292294 201430 292350
rect 201498 292294 201554 292350
rect 201622 292294 201678 292350
rect 201250 292170 201306 292226
rect 201374 292170 201430 292226
rect 201498 292170 201554 292226
rect 201622 292170 201678 292226
rect 201250 292046 201306 292102
rect 201374 292046 201430 292102
rect 201498 292046 201554 292102
rect 201622 292046 201678 292102
rect 201250 291922 201306 291978
rect 201374 291922 201430 291978
rect 201498 291922 201554 291978
rect 201622 291922 201678 291978
rect 201250 274294 201306 274350
rect 201374 274294 201430 274350
rect 201498 274294 201554 274350
rect 201622 274294 201678 274350
rect 201250 274170 201306 274226
rect 201374 274170 201430 274226
rect 201498 274170 201554 274226
rect 201622 274170 201678 274226
rect 201250 274046 201306 274102
rect 201374 274046 201430 274102
rect 201498 274046 201554 274102
rect 201622 274046 201678 274102
rect 201250 273922 201306 273978
rect 201374 273922 201430 273978
rect 201498 273922 201554 273978
rect 201622 273922 201678 273978
rect 201250 256294 201306 256350
rect 201374 256294 201430 256350
rect 201498 256294 201554 256350
rect 201622 256294 201678 256350
rect 201250 256170 201306 256226
rect 201374 256170 201430 256226
rect 201498 256170 201554 256226
rect 201622 256170 201678 256226
rect 201250 256046 201306 256102
rect 201374 256046 201430 256102
rect 201498 256046 201554 256102
rect 201622 256046 201678 256102
rect 201250 255922 201306 255978
rect 201374 255922 201430 255978
rect 201498 255922 201554 255978
rect 201622 255922 201678 255978
rect 201250 238294 201306 238350
rect 201374 238294 201430 238350
rect 201498 238294 201554 238350
rect 201622 238294 201678 238350
rect 201250 238170 201306 238226
rect 201374 238170 201430 238226
rect 201498 238170 201554 238226
rect 201622 238170 201678 238226
rect 201250 238046 201306 238102
rect 201374 238046 201430 238102
rect 201498 238046 201554 238102
rect 201622 238046 201678 238102
rect 201250 237922 201306 237978
rect 201374 237922 201430 237978
rect 201498 237922 201554 237978
rect 201622 237922 201678 237978
rect 201250 220294 201306 220350
rect 201374 220294 201430 220350
rect 201498 220294 201554 220350
rect 201622 220294 201678 220350
rect 201250 220170 201306 220226
rect 201374 220170 201430 220226
rect 201498 220170 201554 220226
rect 201622 220170 201678 220226
rect 201250 220046 201306 220102
rect 201374 220046 201430 220102
rect 201498 220046 201554 220102
rect 201622 220046 201678 220102
rect 201250 219922 201306 219978
rect 201374 219922 201430 219978
rect 201498 219922 201554 219978
rect 201622 219922 201678 219978
rect 201250 202294 201306 202350
rect 201374 202294 201430 202350
rect 201498 202294 201554 202350
rect 201622 202294 201678 202350
rect 201250 202170 201306 202226
rect 201374 202170 201430 202226
rect 201498 202170 201554 202226
rect 201622 202170 201678 202226
rect 201250 202046 201306 202102
rect 201374 202046 201430 202102
rect 201498 202046 201554 202102
rect 201622 202046 201678 202102
rect 201250 201922 201306 201978
rect 201374 201922 201430 201978
rect 201498 201922 201554 201978
rect 201622 201922 201678 201978
rect 201250 184294 201306 184350
rect 201374 184294 201430 184350
rect 201498 184294 201554 184350
rect 201622 184294 201678 184350
rect 201250 184170 201306 184226
rect 201374 184170 201430 184226
rect 201498 184170 201554 184226
rect 201622 184170 201678 184226
rect 201250 184046 201306 184102
rect 201374 184046 201430 184102
rect 201498 184046 201554 184102
rect 201622 184046 201678 184102
rect 201250 183922 201306 183978
rect 201374 183922 201430 183978
rect 201498 183922 201554 183978
rect 201622 183922 201678 183978
rect 201250 166294 201306 166350
rect 201374 166294 201430 166350
rect 201498 166294 201554 166350
rect 201622 166294 201678 166350
rect 201250 166170 201306 166226
rect 201374 166170 201430 166226
rect 201498 166170 201554 166226
rect 201622 166170 201678 166226
rect 201250 166046 201306 166102
rect 201374 166046 201430 166102
rect 201498 166046 201554 166102
rect 201622 166046 201678 166102
rect 201250 165922 201306 165978
rect 201374 165922 201430 165978
rect 201498 165922 201554 165978
rect 201622 165922 201678 165978
rect 201250 148294 201306 148350
rect 201374 148294 201430 148350
rect 201498 148294 201554 148350
rect 201622 148294 201678 148350
rect 201250 148170 201306 148226
rect 201374 148170 201430 148226
rect 201498 148170 201554 148226
rect 201622 148170 201678 148226
rect 201250 148046 201306 148102
rect 201374 148046 201430 148102
rect 201498 148046 201554 148102
rect 201622 148046 201678 148102
rect 201250 147922 201306 147978
rect 201374 147922 201430 147978
rect 201498 147922 201554 147978
rect 201622 147922 201678 147978
rect 201250 130294 201306 130350
rect 201374 130294 201430 130350
rect 201498 130294 201554 130350
rect 201622 130294 201678 130350
rect 201250 130170 201306 130226
rect 201374 130170 201430 130226
rect 201498 130170 201554 130226
rect 201622 130170 201678 130226
rect 201250 130046 201306 130102
rect 201374 130046 201430 130102
rect 201498 130046 201554 130102
rect 201622 130046 201678 130102
rect 201250 129922 201306 129978
rect 201374 129922 201430 129978
rect 201498 129922 201554 129978
rect 201622 129922 201678 129978
rect 201250 112294 201306 112350
rect 201374 112294 201430 112350
rect 201498 112294 201554 112350
rect 201622 112294 201678 112350
rect 201250 112170 201306 112226
rect 201374 112170 201430 112226
rect 201498 112170 201554 112226
rect 201622 112170 201678 112226
rect 201250 112046 201306 112102
rect 201374 112046 201430 112102
rect 201498 112046 201554 112102
rect 201622 112046 201678 112102
rect 201250 111922 201306 111978
rect 201374 111922 201430 111978
rect 201498 111922 201554 111978
rect 201622 111922 201678 111978
rect 201250 94294 201306 94350
rect 201374 94294 201430 94350
rect 201498 94294 201554 94350
rect 201622 94294 201678 94350
rect 201250 94170 201306 94226
rect 201374 94170 201430 94226
rect 201498 94170 201554 94226
rect 201622 94170 201678 94226
rect 201250 94046 201306 94102
rect 201374 94046 201430 94102
rect 201498 94046 201554 94102
rect 201622 94046 201678 94102
rect 201250 93922 201306 93978
rect 201374 93922 201430 93978
rect 201498 93922 201554 93978
rect 201622 93922 201678 93978
rect 201250 76294 201306 76350
rect 201374 76294 201430 76350
rect 201498 76294 201554 76350
rect 201622 76294 201678 76350
rect 201250 76170 201306 76226
rect 201374 76170 201430 76226
rect 201498 76170 201554 76226
rect 201622 76170 201678 76226
rect 201250 76046 201306 76102
rect 201374 76046 201430 76102
rect 201498 76046 201554 76102
rect 201622 76046 201678 76102
rect 201250 75922 201306 75978
rect 201374 75922 201430 75978
rect 201498 75922 201554 75978
rect 201622 75922 201678 75978
rect 201250 58294 201306 58350
rect 201374 58294 201430 58350
rect 201498 58294 201554 58350
rect 201622 58294 201678 58350
rect 201250 58170 201306 58226
rect 201374 58170 201430 58226
rect 201498 58170 201554 58226
rect 201622 58170 201678 58226
rect 201250 58046 201306 58102
rect 201374 58046 201430 58102
rect 201498 58046 201554 58102
rect 201622 58046 201678 58102
rect 201250 57922 201306 57978
rect 201374 57922 201430 57978
rect 201498 57922 201554 57978
rect 201622 57922 201678 57978
rect 201250 40294 201306 40350
rect 201374 40294 201430 40350
rect 201498 40294 201554 40350
rect 201622 40294 201678 40350
rect 201250 40170 201306 40226
rect 201374 40170 201430 40226
rect 201498 40170 201554 40226
rect 201622 40170 201678 40226
rect 201250 40046 201306 40102
rect 201374 40046 201430 40102
rect 201498 40046 201554 40102
rect 201622 40046 201678 40102
rect 201250 39922 201306 39978
rect 201374 39922 201430 39978
rect 201498 39922 201554 39978
rect 201622 39922 201678 39978
rect 201250 22294 201306 22350
rect 201374 22294 201430 22350
rect 201498 22294 201554 22350
rect 201622 22294 201678 22350
rect 201250 22170 201306 22226
rect 201374 22170 201430 22226
rect 201498 22170 201554 22226
rect 201622 22170 201678 22226
rect 201250 22046 201306 22102
rect 201374 22046 201430 22102
rect 201498 22046 201554 22102
rect 201622 22046 201678 22102
rect 201250 21922 201306 21978
rect 201374 21922 201430 21978
rect 201498 21922 201554 21978
rect 201622 21922 201678 21978
rect 201250 4294 201306 4350
rect 201374 4294 201430 4350
rect 201498 4294 201554 4350
rect 201622 4294 201678 4350
rect 201250 4170 201306 4226
rect 201374 4170 201430 4226
rect 201498 4170 201554 4226
rect 201622 4170 201678 4226
rect 201250 4046 201306 4102
rect 201374 4046 201430 4102
rect 201498 4046 201554 4102
rect 201622 4046 201678 4102
rect 201250 3922 201306 3978
rect 201374 3922 201430 3978
rect 201498 3922 201554 3978
rect 201622 3922 201678 3978
rect 186970 -1176 187026 -1120
rect 187094 -1176 187150 -1120
rect 187218 -1176 187274 -1120
rect 187342 -1176 187398 -1120
rect 186970 -1300 187026 -1244
rect 187094 -1300 187150 -1244
rect 187218 -1300 187274 -1244
rect 187342 -1300 187398 -1244
rect 186970 -1424 187026 -1368
rect 187094 -1424 187150 -1368
rect 187218 -1424 187274 -1368
rect 187342 -1424 187398 -1368
rect 186970 -1548 187026 -1492
rect 187094 -1548 187150 -1492
rect 187218 -1548 187274 -1492
rect 187342 -1548 187398 -1492
rect 201250 -216 201306 -160
rect 201374 -216 201430 -160
rect 201498 -216 201554 -160
rect 201622 -216 201678 -160
rect 201250 -340 201306 -284
rect 201374 -340 201430 -284
rect 201498 -340 201554 -284
rect 201622 -340 201678 -284
rect 201250 -464 201306 -408
rect 201374 -464 201430 -408
rect 201498 -464 201554 -408
rect 201622 -464 201678 -408
rect 201250 -588 201306 -532
rect 201374 -588 201430 -532
rect 201498 -588 201554 -532
rect 201622 -588 201678 -532
rect 204970 598116 205026 598172
rect 205094 598116 205150 598172
rect 205218 598116 205274 598172
rect 205342 598116 205398 598172
rect 204970 597992 205026 598048
rect 205094 597992 205150 598048
rect 205218 597992 205274 598048
rect 205342 597992 205398 598048
rect 204970 597868 205026 597924
rect 205094 597868 205150 597924
rect 205218 597868 205274 597924
rect 205342 597868 205398 597924
rect 204970 597744 205026 597800
rect 205094 597744 205150 597800
rect 205218 597744 205274 597800
rect 205342 597744 205398 597800
rect 204970 586294 205026 586350
rect 205094 586294 205150 586350
rect 205218 586294 205274 586350
rect 205342 586294 205398 586350
rect 204970 586170 205026 586226
rect 205094 586170 205150 586226
rect 205218 586170 205274 586226
rect 205342 586170 205398 586226
rect 204970 586046 205026 586102
rect 205094 586046 205150 586102
rect 205218 586046 205274 586102
rect 205342 586046 205398 586102
rect 204970 585922 205026 585978
rect 205094 585922 205150 585978
rect 205218 585922 205274 585978
rect 205342 585922 205398 585978
rect 204970 568294 205026 568350
rect 205094 568294 205150 568350
rect 205218 568294 205274 568350
rect 205342 568294 205398 568350
rect 204970 568170 205026 568226
rect 205094 568170 205150 568226
rect 205218 568170 205274 568226
rect 205342 568170 205398 568226
rect 204970 568046 205026 568102
rect 205094 568046 205150 568102
rect 205218 568046 205274 568102
rect 205342 568046 205398 568102
rect 204970 567922 205026 567978
rect 205094 567922 205150 567978
rect 205218 567922 205274 567978
rect 205342 567922 205398 567978
rect 204970 550294 205026 550350
rect 205094 550294 205150 550350
rect 205218 550294 205274 550350
rect 205342 550294 205398 550350
rect 204970 550170 205026 550226
rect 205094 550170 205150 550226
rect 205218 550170 205274 550226
rect 205342 550170 205398 550226
rect 204970 550046 205026 550102
rect 205094 550046 205150 550102
rect 205218 550046 205274 550102
rect 205342 550046 205398 550102
rect 204970 549922 205026 549978
rect 205094 549922 205150 549978
rect 205218 549922 205274 549978
rect 205342 549922 205398 549978
rect 204970 532294 205026 532350
rect 205094 532294 205150 532350
rect 205218 532294 205274 532350
rect 205342 532294 205398 532350
rect 204970 532170 205026 532226
rect 205094 532170 205150 532226
rect 205218 532170 205274 532226
rect 205342 532170 205398 532226
rect 204970 532046 205026 532102
rect 205094 532046 205150 532102
rect 205218 532046 205274 532102
rect 205342 532046 205398 532102
rect 204970 531922 205026 531978
rect 205094 531922 205150 531978
rect 205218 531922 205274 531978
rect 205342 531922 205398 531978
rect 204970 514294 205026 514350
rect 205094 514294 205150 514350
rect 205218 514294 205274 514350
rect 205342 514294 205398 514350
rect 204970 514170 205026 514226
rect 205094 514170 205150 514226
rect 205218 514170 205274 514226
rect 205342 514170 205398 514226
rect 204970 514046 205026 514102
rect 205094 514046 205150 514102
rect 205218 514046 205274 514102
rect 205342 514046 205398 514102
rect 204970 513922 205026 513978
rect 205094 513922 205150 513978
rect 205218 513922 205274 513978
rect 205342 513922 205398 513978
rect 204970 496294 205026 496350
rect 205094 496294 205150 496350
rect 205218 496294 205274 496350
rect 205342 496294 205398 496350
rect 204970 496170 205026 496226
rect 205094 496170 205150 496226
rect 205218 496170 205274 496226
rect 205342 496170 205398 496226
rect 204970 496046 205026 496102
rect 205094 496046 205150 496102
rect 205218 496046 205274 496102
rect 205342 496046 205398 496102
rect 204970 495922 205026 495978
rect 205094 495922 205150 495978
rect 205218 495922 205274 495978
rect 205342 495922 205398 495978
rect 204970 478294 205026 478350
rect 205094 478294 205150 478350
rect 205218 478294 205274 478350
rect 205342 478294 205398 478350
rect 204970 478170 205026 478226
rect 205094 478170 205150 478226
rect 205218 478170 205274 478226
rect 205342 478170 205398 478226
rect 204970 478046 205026 478102
rect 205094 478046 205150 478102
rect 205218 478046 205274 478102
rect 205342 478046 205398 478102
rect 204970 477922 205026 477978
rect 205094 477922 205150 477978
rect 205218 477922 205274 477978
rect 205342 477922 205398 477978
rect 204970 460294 205026 460350
rect 205094 460294 205150 460350
rect 205218 460294 205274 460350
rect 205342 460294 205398 460350
rect 204970 460170 205026 460226
rect 205094 460170 205150 460226
rect 205218 460170 205274 460226
rect 205342 460170 205398 460226
rect 204970 460046 205026 460102
rect 205094 460046 205150 460102
rect 205218 460046 205274 460102
rect 205342 460046 205398 460102
rect 204970 459922 205026 459978
rect 205094 459922 205150 459978
rect 205218 459922 205274 459978
rect 205342 459922 205398 459978
rect 219250 597156 219306 597212
rect 219374 597156 219430 597212
rect 219498 597156 219554 597212
rect 219622 597156 219678 597212
rect 219250 597032 219306 597088
rect 219374 597032 219430 597088
rect 219498 597032 219554 597088
rect 219622 597032 219678 597088
rect 219250 596908 219306 596964
rect 219374 596908 219430 596964
rect 219498 596908 219554 596964
rect 219622 596908 219678 596964
rect 219250 596784 219306 596840
rect 219374 596784 219430 596840
rect 219498 596784 219554 596840
rect 219622 596784 219678 596840
rect 219250 580294 219306 580350
rect 219374 580294 219430 580350
rect 219498 580294 219554 580350
rect 219622 580294 219678 580350
rect 219250 580170 219306 580226
rect 219374 580170 219430 580226
rect 219498 580170 219554 580226
rect 219622 580170 219678 580226
rect 219250 580046 219306 580102
rect 219374 580046 219430 580102
rect 219498 580046 219554 580102
rect 219622 580046 219678 580102
rect 219250 579922 219306 579978
rect 219374 579922 219430 579978
rect 219498 579922 219554 579978
rect 219622 579922 219678 579978
rect 219250 562294 219306 562350
rect 219374 562294 219430 562350
rect 219498 562294 219554 562350
rect 219622 562294 219678 562350
rect 219250 562170 219306 562226
rect 219374 562170 219430 562226
rect 219498 562170 219554 562226
rect 219622 562170 219678 562226
rect 219250 562046 219306 562102
rect 219374 562046 219430 562102
rect 219498 562046 219554 562102
rect 219622 562046 219678 562102
rect 219250 561922 219306 561978
rect 219374 561922 219430 561978
rect 219498 561922 219554 561978
rect 219622 561922 219678 561978
rect 219250 544294 219306 544350
rect 219374 544294 219430 544350
rect 219498 544294 219554 544350
rect 219622 544294 219678 544350
rect 219250 544170 219306 544226
rect 219374 544170 219430 544226
rect 219498 544170 219554 544226
rect 219622 544170 219678 544226
rect 219250 544046 219306 544102
rect 219374 544046 219430 544102
rect 219498 544046 219554 544102
rect 219622 544046 219678 544102
rect 219250 543922 219306 543978
rect 219374 543922 219430 543978
rect 219498 543922 219554 543978
rect 219622 543922 219678 543978
rect 219250 526294 219306 526350
rect 219374 526294 219430 526350
rect 219498 526294 219554 526350
rect 219622 526294 219678 526350
rect 219250 526170 219306 526226
rect 219374 526170 219430 526226
rect 219498 526170 219554 526226
rect 219622 526170 219678 526226
rect 219250 526046 219306 526102
rect 219374 526046 219430 526102
rect 219498 526046 219554 526102
rect 219622 526046 219678 526102
rect 219250 525922 219306 525978
rect 219374 525922 219430 525978
rect 219498 525922 219554 525978
rect 219622 525922 219678 525978
rect 219250 508294 219306 508350
rect 219374 508294 219430 508350
rect 219498 508294 219554 508350
rect 219622 508294 219678 508350
rect 219250 508170 219306 508226
rect 219374 508170 219430 508226
rect 219498 508170 219554 508226
rect 219622 508170 219678 508226
rect 219250 508046 219306 508102
rect 219374 508046 219430 508102
rect 219498 508046 219554 508102
rect 219622 508046 219678 508102
rect 219250 507922 219306 507978
rect 219374 507922 219430 507978
rect 219498 507922 219554 507978
rect 219622 507922 219678 507978
rect 219250 490294 219306 490350
rect 219374 490294 219430 490350
rect 219498 490294 219554 490350
rect 219622 490294 219678 490350
rect 219250 490170 219306 490226
rect 219374 490170 219430 490226
rect 219498 490170 219554 490226
rect 219622 490170 219678 490226
rect 219250 490046 219306 490102
rect 219374 490046 219430 490102
rect 219498 490046 219554 490102
rect 219622 490046 219678 490102
rect 219250 489922 219306 489978
rect 219374 489922 219430 489978
rect 219498 489922 219554 489978
rect 219622 489922 219678 489978
rect 219250 472294 219306 472350
rect 219374 472294 219430 472350
rect 219498 472294 219554 472350
rect 219622 472294 219678 472350
rect 219250 472170 219306 472226
rect 219374 472170 219430 472226
rect 219498 472170 219554 472226
rect 219622 472170 219678 472226
rect 219250 472046 219306 472102
rect 219374 472046 219430 472102
rect 219498 472046 219554 472102
rect 219622 472046 219678 472102
rect 219250 471922 219306 471978
rect 219374 471922 219430 471978
rect 219498 471922 219554 471978
rect 219622 471922 219678 471978
rect 222970 598116 223026 598172
rect 223094 598116 223150 598172
rect 223218 598116 223274 598172
rect 223342 598116 223398 598172
rect 222970 597992 223026 598048
rect 223094 597992 223150 598048
rect 223218 597992 223274 598048
rect 223342 597992 223398 598048
rect 222970 597868 223026 597924
rect 223094 597868 223150 597924
rect 223218 597868 223274 597924
rect 223342 597868 223398 597924
rect 222970 597744 223026 597800
rect 223094 597744 223150 597800
rect 223218 597744 223274 597800
rect 223342 597744 223398 597800
rect 222970 586294 223026 586350
rect 223094 586294 223150 586350
rect 223218 586294 223274 586350
rect 223342 586294 223398 586350
rect 222970 586170 223026 586226
rect 223094 586170 223150 586226
rect 223218 586170 223274 586226
rect 223342 586170 223398 586226
rect 222970 586046 223026 586102
rect 223094 586046 223150 586102
rect 223218 586046 223274 586102
rect 223342 586046 223398 586102
rect 222970 585922 223026 585978
rect 223094 585922 223150 585978
rect 223218 585922 223274 585978
rect 223342 585922 223398 585978
rect 222970 568294 223026 568350
rect 223094 568294 223150 568350
rect 223218 568294 223274 568350
rect 223342 568294 223398 568350
rect 222970 568170 223026 568226
rect 223094 568170 223150 568226
rect 223218 568170 223274 568226
rect 223342 568170 223398 568226
rect 222970 568046 223026 568102
rect 223094 568046 223150 568102
rect 223218 568046 223274 568102
rect 223342 568046 223398 568102
rect 222970 567922 223026 567978
rect 223094 567922 223150 567978
rect 223218 567922 223274 567978
rect 223342 567922 223398 567978
rect 222970 550294 223026 550350
rect 223094 550294 223150 550350
rect 223218 550294 223274 550350
rect 223342 550294 223398 550350
rect 222970 550170 223026 550226
rect 223094 550170 223150 550226
rect 223218 550170 223274 550226
rect 223342 550170 223398 550226
rect 222970 550046 223026 550102
rect 223094 550046 223150 550102
rect 223218 550046 223274 550102
rect 223342 550046 223398 550102
rect 222970 549922 223026 549978
rect 223094 549922 223150 549978
rect 223218 549922 223274 549978
rect 223342 549922 223398 549978
rect 222970 532294 223026 532350
rect 223094 532294 223150 532350
rect 223218 532294 223274 532350
rect 223342 532294 223398 532350
rect 222970 532170 223026 532226
rect 223094 532170 223150 532226
rect 223218 532170 223274 532226
rect 223342 532170 223398 532226
rect 222970 532046 223026 532102
rect 223094 532046 223150 532102
rect 223218 532046 223274 532102
rect 223342 532046 223398 532102
rect 222970 531922 223026 531978
rect 223094 531922 223150 531978
rect 223218 531922 223274 531978
rect 223342 531922 223398 531978
rect 222970 514294 223026 514350
rect 223094 514294 223150 514350
rect 223218 514294 223274 514350
rect 223342 514294 223398 514350
rect 222970 514170 223026 514226
rect 223094 514170 223150 514226
rect 223218 514170 223274 514226
rect 223342 514170 223398 514226
rect 222970 514046 223026 514102
rect 223094 514046 223150 514102
rect 223218 514046 223274 514102
rect 223342 514046 223398 514102
rect 222970 513922 223026 513978
rect 223094 513922 223150 513978
rect 223218 513922 223274 513978
rect 223342 513922 223398 513978
rect 222970 496294 223026 496350
rect 223094 496294 223150 496350
rect 223218 496294 223274 496350
rect 223342 496294 223398 496350
rect 222970 496170 223026 496226
rect 223094 496170 223150 496226
rect 223218 496170 223274 496226
rect 223342 496170 223398 496226
rect 222970 496046 223026 496102
rect 223094 496046 223150 496102
rect 223218 496046 223274 496102
rect 223342 496046 223398 496102
rect 222970 495922 223026 495978
rect 223094 495922 223150 495978
rect 223218 495922 223274 495978
rect 223342 495922 223398 495978
rect 222970 478294 223026 478350
rect 223094 478294 223150 478350
rect 223218 478294 223274 478350
rect 223342 478294 223398 478350
rect 222970 478170 223026 478226
rect 223094 478170 223150 478226
rect 223218 478170 223274 478226
rect 223342 478170 223398 478226
rect 222970 478046 223026 478102
rect 223094 478046 223150 478102
rect 223218 478046 223274 478102
rect 223342 478046 223398 478102
rect 222970 477922 223026 477978
rect 223094 477922 223150 477978
rect 223218 477922 223274 477978
rect 223342 477922 223398 477978
rect 222970 460294 223026 460350
rect 223094 460294 223150 460350
rect 223218 460294 223274 460350
rect 223342 460294 223398 460350
rect 222970 460170 223026 460226
rect 223094 460170 223150 460226
rect 223218 460170 223274 460226
rect 223342 460170 223398 460226
rect 222970 460046 223026 460102
rect 223094 460046 223150 460102
rect 223218 460046 223274 460102
rect 223342 460046 223398 460102
rect 222970 459922 223026 459978
rect 223094 459922 223150 459978
rect 223218 459922 223274 459978
rect 223342 459922 223398 459978
rect 237250 597156 237306 597212
rect 237374 597156 237430 597212
rect 237498 597156 237554 597212
rect 237622 597156 237678 597212
rect 237250 597032 237306 597088
rect 237374 597032 237430 597088
rect 237498 597032 237554 597088
rect 237622 597032 237678 597088
rect 237250 596908 237306 596964
rect 237374 596908 237430 596964
rect 237498 596908 237554 596964
rect 237622 596908 237678 596964
rect 237250 596784 237306 596840
rect 237374 596784 237430 596840
rect 237498 596784 237554 596840
rect 237622 596784 237678 596840
rect 237250 580294 237306 580350
rect 237374 580294 237430 580350
rect 237498 580294 237554 580350
rect 237622 580294 237678 580350
rect 237250 580170 237306 580226
rect 237374 580170 237430 580226
rect 237498 580170 237554 580226
rect 237622 580170 237678 580226
rect 237250 580046 237306 580102
rect 237374 580046 237430 580102
rect 237498 580046 237554 580102
rect 237622 580046 237678 580102
rect 237250 579922 237306 579978
rect 237374 579922 237430 579978
rect 237498 579922 237554 579978
rect 237622 579922 237678 579978
rect 237250 562294 237306 562350
rect 237374 562294 237430 562350
rect 237498 562294 237554 562350
rect 237622 562294 237678 562350
rect 237250 562170 237306 562226
rect 237374 562170 237430 562226
rect 237498 562170 237554 562226
rect 237622 562170 237678 562226
rect 237250 562046 237306 562102
rect 237374 562046 237430 562102
rect 237498 562046 237554 562102
rect 237622 562046 237678 562102
rect 237250 561922 237306 561978
rect 237374 561922 237430 561978
rect 237498 561922 237554 561978
rect 237622 561922 237678 561978
rect 237250 544294 237306 544350
rect 237374 544294 237430 544350
rect 237498 544294 237554 544350
rect 237622 544294 237678 544350
rect 237250 544170 237306 544226
rect 237374 544170 237430 544226
rect 237498 544170 237554 544226
rect 237622 544170 237678 544226
rect 237250 544046 237306 544102
rect 237374 544046 237430 544102
rect 237498 544046 237554 544102
rect 237622 544046 237678 544102
rect 237250 543922 237306 543978
rect 237374 543922 237430 543978
rect 237498 543922 237554 543978
rect 237622 543922 237678 543978
rect 237250 526294 237306 526350
rect 237374 526294 237430 526350
rect 237498 526294 237554 526350
rect 237622 526294 237678 526350
rect 237250 526170 237306 526226
rect 237374 526170 237430 526226
rect 237498 526170 237554 526226
rect 237622 526170 237678 526226
rect 237250 526046 237306 526102
rect 237374 526046 237430 526102
rect 237498 526046 237554 526102
rect 237622 526046 237678 526102
rect 237250 525922 237306 525978
rect 237374 525922 237430 525978
rect 237498 525922 237554 525978
rect 237622 525922 237678 525978
rect 237250 508294 237306 508350
rect 237374 508294 237430 508350
rect 237498 508294 237554 508350
rect 237622 508294 237678 508350
rect 237250 508170 237306 508226
rect 237374 508170 237430 508226
rect 237498 508170 237554 508226
rect 237622 508170 237678 508226
rect 237250 508046 237306 508102
rect 237374 508046 237430 508102
rect 237498 508046 237554 508102
rect 237622 508046 237678 508102
rect 237250 507922 237306 507978
rect 237374 507922 237430 507978
rect 237498 507922 237554 507978
rect 237622 507922 237678 507978
rect 237250 490294 237306 490350
rect 237374 490294 237430 490350
rect 237498 490294 237554 490350
rect 237622 490294 237678 490350
rect 237250 490170 237306 490226
rect 237374 490170 237430 490226
rect 237498 490170 237554 490226
rect 237622 490170 237678 490226
rect 237250 490046 237306 490102
rect 237374 490046 237430 490102
rect 237498 490046 237554 490102
rect 237622 490046 237678 490102
rect 237250 489922 237306 489978
rect 237374 489922 237430 489978
rect 237498 489922 237554 489978
rect 237622 489922 237678 489978
rect 237250 472294 237306 472350
rect 237374 472294 237430 472350
rect 237498 472294 237554 472350
rect 237622 472294 237678 472350
rect 237250 472170 237306 472226
rect 237374 472170 237430 472226
rect 237498 472170 237554 472226
rect 237622 472170 237678 472226
rect 237250 472046 237306 472102
rect 237374 472046 237430 472102
rect 237498 472046 237554 472102
rect 237622 472046 237678 472102
rect 237250 471922 237306 471978
rect 237374 471922 237430 471978
rect 237498 471922 237554 471978
rect 237622 471922 237678 471978
rect 240970 598116 241026 598172
rect 241094 598116 241150 598172
rect 241218 598116 241274 598172
rect 241342 598116 241398 598172
rect 240970 597992 241026 598048
rect 241094 597992 241150 598048
rect 241218 597992 241274 598048
rect 241342 597992 241398 598048
rect 240970 597868 241026 597924
rect 241094 597868 241150 597924
rect 241218 597868 241274 597924
rect 241342 597868 241398 597924
rect 240970 597744 241026 597800
rect 241094 597744 241150 597800
rect 241218 597744 241274 597800
rect 241342 597744 241398 597800
rect 240970 586294 241026 586350
rect 241094 586294 241150 586350
rect 241218 586294 241274 586350
rect 241342 586294 241398 586350
rect 240970 586170 241026 586226
rect 241094 586170 241150 586226
rect 241218 586170 241274 586226
rect 241342 586170 241398 586226
rect 240970 586046 241026 586102
rect 241094 586046 241150 586102
rect 241218 586046 241274 586102
rect 241342 586046 241398 586102
rect 240970 585922 241026 585978
rect 241094 585922 241150 585978
rect 241218 585922 241274 585978
rect 241342 585922 241398 585978
rect 240970 568294 241026 568350
rect 241094 568294 241150 568350
rect 241218 568294 241274 568350
rect 241342 568294 241398 568350
rect 240970 568170 241026 568226
rect 241094 568170 241150 568226
rect 241218 568170 241274 568226
rect 241342 568170 241398 568226
rect 240970 568046 241026 568102
rect 241094 568046 241150 568102
rect 241218 568046 241274 568102
rect 241342 568046 241398 568102
rect 240970 567922 241026 567978
rect 241094 567922 241150 567978
rect 241218 567922 241274 567978
rect 241342 567922 241398 567978
rect 240970 550294 241026 550350
rect 241094 550294 241150 550350
rect 241218 550294 241274 550350
rect 241342 550294 241398 550350
rect 240970 550170 241026 550226
rect 241094 550170 241150 550226
rect 241218 550170 241274 550226
rect 241342 550170 241398 550226
rect 240970 550046 241026 550102
rect 241094 550046 241150 550102
rect 241218 550046 241274 550102
rect 241342 550046 241398 550102
rect 240970 549922 241026 549978
rect 241094 549922 241150 549978
rect 241218 549922 241274 549978
rect 241342 549922 241398 549978
rect 240970 532294 241026 532350
rect 241094 532294 241150 532350
rect 241218 532294 241274 532350
rect 241342 532294 241398 532350
rect 240970 532170 241026 532226
rect 241094 532170 241150 532226
rect 241218 532170 241274 532226
rect 241342 532170 241398 532226
rect 240970 532046 241026 532102
rect 241094 532046 241150 532102
rect 241218 532046 241274 532102
rect 241342 532046 241398 532102
rect 240970 531922 241026 531978
rect 241094 531922 241150 531978
rect 241218 531922 241274 531978
rect 241342 531922 241398 531978
rect 240970 514294 241026 514350
rect 241094 514294 241150 514350
rect 241218 514294 241274 514350
rect 241342 514294 241398 514350
rect 240970 514170 241026 514226
rect 241094 514170 241150 514226
rect 241218 514170 241274 514226
rect 241342 514170 241398 514226
rect 240970 514046 241026 514102
rect 241094 514046 241150 514102
rect 241218 514046 241274 514102
rect 241342 514046 241398 514102
rect 240970 513922 241026 513978
rect 241094 513922 241150 513978
rect 241218 513922 241274 513978
rect 241342 513922 241398 513978
rect 240970 496294 241026 496350
rect 241094 496294 241150 496350
rect 241218 496294 241274 496350
rect 241342 496294 241398 496350
rect 240970 496170 241026 496226
rect 241094 496170 241150 496226
rect 241218 496170 241274 496226
rect 241342 496170 241398 496226
rect 240970 496046 241026 496102
rect 241094 496046 241150 496102
rect 241218 496046 241274 496102
rect 241342 496046 241398 496102
rect 240970 495922 241026 495978
rect 241094 495922 241150 495978
rect 241218 495922 241274 495978
rect 241342 495922 241398 495978
rect 240970 478294 241026 478350
rect 241094 478294 241150 478350
rect 241218 478294 241274 478350
rect 241342 478294 241398 478350
rect 240970 478170 241026 478226
rect 241094 478170 241150 478226
rect 241218 478170 241274 478226
rect 241342 478170 241398 478226
rect 240970 478046 241026 478102
rect 241094 478046 241150 478102
rect 241218 478046 241274 478102
rect 241342 478046 241398 478102
rect 240970 477922 241026 477978
rect 241094 477922 241150 477978
rect 241218 477922 241274 477978
rect 241342 477922 241398 477978
rect 240970 460294 241026 460350
rect 241094 460294 241150 460350
rect 241218 460294 241274 460350
rect 241342 460294 241398 460350
rect 240970 460170 241026 460226
rect 241094 460170 241150 460226
rect 241218 460170 241274 460226
rect 241342 460170 241398 460226
rect 240970 460046 241026 460102
rect 241094 460046 241150 460102
rect 241218 460046 241274 460102
rect 241342 460046 241398 460102
rect 240970 459922 241026 459978
rect 241094 459922 241150 459978
rect 241218 459922 241274 459978
rect 241342 459922 241398 459978
rect 255250 597156 255306 597212
rect 255374 597156 255430 597212
rect 255498 597156 255554 597212
rect 255622 597156 255678 597212
rect 255250 597032 255306 597088
rect 255374 597032 255430 597088
rect 255498 597032 255554 597088
rect 255622 597032 255678 597088
rect 255250 596908 255306 596964
rect 255374 596908 255430 596964
rect 255498 596908 255554 596964
rect 255622 596908 255678 596964
rect 255250 596784 255306 596840
rect 255374 596784 255430 596840
rect 255498 596784 255554 596840
rect 255622 596784 255678 596840
rect 255250 580294 255306 580350
rect 255374 580294 255430 580350
rect 255498 580294 255554 580350
rect 255622 580294 255678 580350
rect 255250 580170 255306 580226
rect 255374 580170 255430 580226
rect 255498 580170 255554 580226
rect 255622 580170 255678 580226
rect 255250 580046 255306 580102
rect 255374 580046 255430 580102
rect 255498 580046 255554 580102
rect 255622 580046 255678 580102
rect 255250 579922 255306 579978
rect 255374 579922 255430 579978
rect 255498 579922 255554 579978
rect 255622 579922 255678 579978
rect 255250 562294 255306 562350
rect 255374 562294 255430 562350
rect 255498 562294 255554 562350
rect 255622 562294 255678 562350
rect 255250 562170 255306 562226
rect 255374 562170 255430 562226
rect 255498 562170 255554 562226
rect 255622 562170 255678 562226
rect 255250 562046 255306 562102
rect 255374 562046 255430 562102
rect 255498 562046 255554 562102
rect 255622 562046 255678 562102
rect 255250 561922 255306 561978
rect 255374 561922 255430 561978
rect 255498 561922 255554 561978
rect 255622 561922 255678 561978
rect 255250 544294 255306 544350
rect 255374 544294 255430 544350
rect 255498 544294 255554 544350
rect 255622 544294 255678 544350
rect 255250 544170 255306 544226
rect 255374 544170 255430 544226
rect 255498 544170 255554 544226
rect 255622 544170 255678 544226
rect 255250 544046 255306 544102
rect 255374 544046 255430 544102
rect 255498 544046 255554 544102
rect 255622 544046 255678 544102
rect 255250 543922 255306 543978
rect 255374 543922 255430 543978
rect 255498 543922 255554 543978
rect 255622 543922 255678 543978
rect 255250 526294 255306 526350
rect 255374 526294 255430 526350
rect 255498 526294 255554 526350
rect 255622 526294 255678 526350
rect 255250 526170 255306 526226
rect 255374 526170 255430 526226
rect 255498 526170 255554 526226
rect 255622 526170 255678 526226
rect 255250 526046 255306 526102
rect 255374 526046 255430 526102
rect 255498 526046 255554 526102
rect 255622 526046 255678 526102
rect 255250 525922 255306 525978
rect 255374 525922 255430 525978
rect 255498 525922 255554 525978
rect 255622 525922 255678 525978
rect 255250 508294 255306 508350
rect 255374 508294 255430 508350
rect 255498 508294 255554 508350
rect 255622 508294 255678 508350
rect 255250 508170 255306 508226
rect 255374 508170 255430 508226
rect 255498 508170 255554 508226
rect 255622 508170 255678 508226
rect 255250 508046 255306 508102
rect 255374 508046 255430 508102
rect 255498 508046 255554 508102
rect 255622 508046 255678 508102
rect 255250 507922 255306 507978
rect 255374 507922 255430 507978
rect 255498 507922 255554 507978
rect 255622 507922 255678 507978
rect 255250 490294 255306 490350
rect 255374 490294 255430 490350
rect 255498 490294 255554 490350
rect 255622 490294 255678 490350
rect 255250 490170 255306 490226
rect 255374 490170 255430 490226
rect 255498 490170 255554 490226
rect 255622 490170 255678 490226
rect 255250 490046 255306 490102
rect 255374 490046 255430 490102
rect 255498 490046 255554 490102
rect 255622 490046 255678 490102
rect 255250 489922 255306 489978
rect 255374 489922 255430 489978
rect 255498 489922 255554 489978
rect 255622 489922 255678 489978
rect 255250 472294 255306 472350
rect 255374 472294 255430 472350
rect 255498 472294 255554 472350
rect 255622 472294 255678 472350
rect 255250 472170 255306 472226
rect 255374 472170 255430 472226
rect 255498 472170 255554 472226
rect 255622 472170 255678 472226
rect 255250 472046 255306 472102
rect 255374 472046 255430 472102
rect 255498 472046 255554 472102
rect 255622 472046 255678 472102
rect 255250 471922 255306 471978
rect 255374 471922 255430 471978
rect 255498 471922 255554 471978
rect 255622 471922 255678 471978
rect 258970 598116 259026 598172
rect 259094 598116 259150 598172
rect 259218 598116 259274 598172
rect 259342 598116 259398 598172
rect 258970 597992 259026 598048
rect 259094 597992 259150 598048
rect 259218 597992 259274 598048
rect 259342 597992 259398 598048
rect 258970 597868 259026 597924
rect 259094 597868 259150 597924
rect 259218 597868 259274 597924
rect 259342 597868 259398 597924
rect 258970 597744 259026 597800
rect 259094 597744 259150 597800
rect 259218 597744 259274 597800
rect 259342 597744 259398 597800
rect 258970 586294 259026 586350
rect 259094 586294 259150 586350
rect 259218 586294 259274 586350
rect 259342 586294 259398 586350
rect 258970 586170 259026 586226
rect 259094 586170 259150 586226
rect 259218 586170 259274 586226
rect 259342 586170 259398 586226
rect 258970 586046 259026 586102
rect 259094 586046 259150 586102
rect 259218 586046 259274 586102
rect 259342 586046 259398 586102
rect 258970 585922 259026 585978
rect 259094 585922 259150 585978
rect 259218 585922 259274 585978
rect 259342 585922 259398 585978
rect 258970 568294 259026 568350
rect 259094 568294 259150 568350
rect 259218 568294 259274 568350
rect 259342 568294 259398 568350
rect 258970 568170 259026 568226
rect 259094 568170 259150 568226
rect 259218 568170 259274 568226
rect 259342 568170 259398 568226
rect 258970 568046 259026 568102
rect 259094 568046 259150 568102
rect 259218 568046 259274 568102
rect 259342 568046 259398 568102
rect 258970 567922 259026 567978
rect 259094 567922 259150 567978
rect 259218 567922 259274 567978
rect 259342 567922 259398 567978
rect 258970 550294 259026 550350
rect 259094 550294 259150 550350
rect 259218 550294 259274 550350
rect 259342 550294 259398 550350
rect 258970 550170 259026 550226
rect 259094 550170 259150 550226
rect 259218 550170 259274 550226
rect 259342 550170 259398 550226
rect 258970 550046 259026 550102
rect 259094 550046 259150 550102
rect 259218 550046 259274 550102
rect 259342 550046 259398 550102
rect 258970 549922 259026 549978
rect 259094 549922 259150 549978
rect 259218 549922 259274 549978
rect 259342 549922 259398 549978
rect 258970 532294 259026 532350
rect 259094 532294 259150 532350
rect 259218 532294 259274 532350
rect 259342 532294 259398 532350
rect 258970 532170 259026 532226
rect 259094 532170 259150 532226
rect 259218 532170 259274 532226
rect 259342 532170 259398 532226
rect 258970 532046 259026 532102
rect 259094 532046 259150 532102
rect 259218 532046 259274 532102
rect 259342 532046 259398 532102
rect 258970 531922 259026 531978
rect 259094 531922 259150 531978
rect 259218 531922 259274 531978
rect 259342 531922 259398 531978
rect 258970 514294 259026 514350
rect 259094 514294 259150 514350
rect 259218 514294 259274 514350
rect 259342 514294 259398 514350
rect 258970 514170 259026 514226
rect 259094 514170 259150 514226
rect 259218 514170 259274 514226
rect 259342 514170 259398 514226
rect 258970 514046 259026 514102
rect 259094 514046 259150 514102
rect 259218 514046 259274 514102
rect 259342 514046 259398 514102
rect 258970 513922 259026 513978
rect 259094 513922 259150 513978
rect 259218 513922 259274 513978
rect 259342 513922 259398 513978
rect 258970 496294 259026 496350
rect 259094 496294 259150 496350
rect 259218 496294 259274 496350
rect 259342 496294 259398 496350
rect 258970 496170 259026 496226
rect 259094 496170 259150 496226
rect 259218 496170 259274 496226
rect 259342 496170 259398 496226
rect 258970 496046 259026 496102
rect 259094 496046 259150 496102
rect 259218 496046 259274 496102
rect 259342 496046 259398 496102
rect 258970 495922 259026 495978
rect 259094 495922 259150 495978
rect 259218 495922 259274 495978
rect 259342 495922 259398 495978
rect 258970 478294 259026 478350
rect 259094 478294 259150 478350
rect 259218 478294 259274 478350
rect 259342 478294 259398 478350
rect 258970 478170 259026 478226
rect 259094 478170 259150 478226
rect 259218 478170 259274 478226
rect 259342 478170 259398 478226
rect 258970 478046 259026 478102
rect 259094 478046 259150 478102
rect 259218 478046 259274 478102
rect 259342 478046 259398 478102
rect 258970 477922 259026 477978
rect 259094 477922 259150 477978
rect 259218 477922 259274 477978
rect 259342 477922 259398 477978
rect 258970 460294 259026 460350
rect 259094 460294 259150 460350
rect 259218 460294 259274 460350
rect 259342 460294 259398 460350
rect 258970 460170 259026 460226
rect 259094 460170 259150 460226
rect 259218 460170 259274 460226
rect 259342 460170 259398 460226
rect 258970 460046 259026 460102
rect 259094 460046 259150 460102
rect 259218 460046 259274 460102
rect 259342 460046 259398 460102
rect 258970 459922 259026 459978
rect 259094 459922 259150 459978
rect 259218 459922 259274 459978
rect 259342 459922 259398 459978
rect 273250 597156 273306 597212
rect 273374 597156 273430 597212
rect 273498 597156 273554 597212
rect 273622 597156 273678 597212
rect 273250 597032 273306 597088
rect 273374 597032 273430 597088
rect 273498 597032 273554 597088
rect 273622 597032 273678 597088
rect 273250 596908 273306 596964
rect 273374 596908 273430 596964
rect 273498 596908 273554 596964
rect 273622 596908 273678 596964
rect 273250 596784 273306 596840
rect 273374 596784 273430 596840
rect 273498 596784 273554 596840
rect 273622 596784 273678 596840
rect 273250 580294 273306 580350
rect 273374 580294 273430 580350
rect 273498 580294 273554 580350
rect 273622 580294 273678 580350
rect 273250 580170 273306 580226
rect 273374 580170 273430 580226
rect 273498 580170 273554 580226
rect 273622 580170 273678 580226
rect 273250 580046 273306 580102
rect 273374 580046 273430 580102
rect 273498 580046 273554 580102
rect 273622 580046 273678 580102
rect 273250 579922 273306 579978
rect 273374 579922 273430 579978
rect 273498 579922 273554 579978
rect 273622 579922 273678 579978
rect 273250 562294 273306 562350
rect 273374 562294 273430 562350
rect 273498 562294 273554 562350
rect 273622 562294 273678 562350
rect 273250 562170 273306 562226
rect 273374 562170 273430 562226
rect 273498 562170 273554 562226
rect 273622 562170 273678 562226
rect 273250 562046 273306 562102
rect 273374 562046 273430 562102
rect 273498 562046 273554 562102
rect 273622 562046 273678 562102
rect 273250 561922 273306 561978
rect 273374 561922 273430 561978
rect 273498 561922 273554 561978
rect 273622 561922 273678 561978
rect 273250 544294 273306 544350
rect 273374 544294 273430 544350
rect 273498 544294 273554 544350
rect 273622 544294 273678 544350
rect 273250 544170 273306 544226
rect 273374 544170 273430 544226
rect 273498 544170 273554 544226
rect 273622 544170 273678 544226
rect 273250 544046 273306 544102
rect 273374 544046 273430 544102
rect 273498 544046 273554 544102
rect 273622 544046 273678 544102
rect 273250 543922 273306 543978
rect 273374 543922 273430 543978
rect 273498 543922 273554 543978
rect 273622 543922 273678 543978
rect 273250 526294 273306 526350
rect 273374 526294 273430 526350
rect 273498 526294 273554 526350
rect 273622 526294 273678 526350
rect 273250 526170 273306 526226
rect 273374 526170 273430 526226
rect 273498 526170 273554 526226
rect 273622 526170 273678 526226
rect 273250 526046 273306 526102
rect 273374 526046 273430 526102
rect 273498 526046 273554 526102
rect 273622 526046 273678 526102
rect 273250 525922 273306 525978
rect 273374 525922 273430 525978
rect 273498 525922 273554 525978
rect 273622 525922 273678 525978
rect 273250 508294 273306 508350
rect 273374 508294 273430 508350
rect 273498 508294 273554 508350
rect 273622 508294 273678 508350
rect 273250 508170 273306 508226
rect 273374 508170 273430 508226
rect 273498 508170 273554 508226
rect 273622 508170 273678 508226
rect 273250 508046 273306 508102
rect 273374 508046 273430 508102
rect 273498 508046 273554 508102
rect 273622 508046 273678 508102
rect 273250 507922 273306 507978
rect 273374 507922 273430 507978
rect 273498 507922 273554 507978
rect 273622 507922 273678 507978
rect 273250 490294 273306 490350
rect 273374 490294 273430 490350
rect 273498 490294 273554 490350
rect 273622 490294 273678 490350
rect 273250 490170 273306 490226
rect 273374 490170 273430 490226
rect 273498 490170 273554 490226
rect 273622 490170 273678 490226
rect 273250 490046 273306 490102
rect 273374 490046 273430 490102
rect 273498 490046 273554 490102
rect 273622 490046 273678 490102
rect 273250 489922 273306 489978
rect 273374 489922 273430 489978
rect 273498 489922 273554 489978
rect 273622 489922 273678 489978
rect 273250 472294 273306 472350
rect 273374 472294 273430 472350
rect 273498 472294 273554 472350
rect 273622 472294 273678 472350
rect 273250 472170 273306 472226
rect 273374 472170 273430 472226
rect 273498 472170 273554 472226
rect 273622 472170 273678 472226
rect 273250 472046 273306 472102
rect 273374 472046 273430 472102
rect 273498 472046 273554 472102
rect 273622 472046 273678 472102
rect 273250 471922 273306 471978
rect 273374 471922 273430 471978
rect 273498 471922 273554 471978
rect 273622 471922 273678 471978
rect 276970 598116 277026 598172
rect 277094 598116 277150 598172
rect 277218 598116 277274 598172
rect 277342 598116 277398 598172
rect 276970 597992 277026 598048
rect 277094 597992 277150 598048
rect 277218 597992 277274 598048
rect 277342 597992 277398 598048
rect 276970 597868 277026 597924
rect 277094 597868 277150 597924
rect 277218 597868 277274 597924
rect 277342 597868 277398 597924
rect 276970 597744 277026 597800
rect 277094 597744 277150 597800
rect 277218 597744 277274 597800
rect 277342 597744 277398 597800
rect 276970 586294 277026 586350
rect 277094 586294 277150 586350
rect 277218 586294 277274 586350
rect 277342 586294 277398 586350
rect 276970 586170 277026 586226
rect 277094 586170 277150 586226
rect 277218 586170 277274 586226
rect 277342 586170 277398 586226
rect 276970 586046 277026 586102
rect 277094 586046 277150 586102
rect 277218 586046 277274 586102
rect 277342 586046 277398 586102
rect 276970 585922 277026 585978
rect 277094 585922 277150 585978
rect 277218 585922 277274 585978
rect 277342 585922 277398 585978
rect 276970 568294 277026 568350
rect 277094 568294 277150 568350
rect 277218 568294 277274 568350
rect 277342 568294 277398 568350
rect 276970 568170 277026 568226
rect 277094 568170 277150 568226
rect 277218 568170 277274 568226
rect 277342 568170 277398 568226
rect 276970 568046 277026 568102
rect 277094 568046 277150 568102
rect 277218 568046 277274 568102
rect 277342 568046 277398 568102
rect 276970 567922 277026 567978
rect 277094 567922 277150 567978
rect 277218 567922 277274 567978
rect 277342 567922 277398 567978
rect 276970 550294 277026 550350
rect 277094 550294 277150 550350
rect 277218 550294 277274 550350
rect 277342 550294 277398 550350
rect 276970 550170 277026 550226
rect 277094 550170 277150 550226
rect 277218 550170 277274 550226
rect 277342 550170 277398 550226
rect 276970 550046 277026 550102
rect 277094 550046 277150 550102
rect 277218 550046 277274 550102
rect 277342 550046 277398 550102
rect 276970 549922 277026 549978
rect 277094 549922 277150 549978
rect 277218 549922 277274 549978
rect 277342 549922 277398 549978
rect 276970 532294 277026 532350
rect 277094 532294 277150 532350
rect 277218 532294 277274 532350
rect 277342 532294 277398 532350
rect 276970 532170 277026 532226
rect 277094 532170 277150 532226
rect 277218 532170 277274 532226
rect 277342 532170 277398 532226
rect 276970 532046 277026 532102
rect 277094 532046 277150 532102
rect 277218 532046 277274 532102
rect 277342 532046 277398 532102
rect 276970 531922 277026 531978
rect 277094 531922 277150 531978
rect 277218 531922 277274 531978
rect 277342 531922 277398 531978
rect 276970 514294 277026 514350
rect 277094 514294 277150 514350
rect 277218 514294 277274 514350
rect 277342 514294 277398 514350
rect 276970 514170 277026 514226
rect 277094 514170 277150 514226
rect 277218 514170 277274 514226
rect 277342 514170 277398 514226
rect 276970 514046 277026 514102
rect 277094 514046 277150 514102
rect 277218 514046 277274 514102
rect 277342 514046 277398 514102
rect 276970 513922 277026 513978
rect 277094 513922 277150 513978
rect 277218 513922 277274 513978
rect 277342 513922 277398 513978
rect 276970 496294 277026 496350
rect 277094 496294 277150 496350
rect 277218 496294 277274 496350
rect 277342 496294 277398 496350
rect 276970 496170 277026 496226
rect 277094 496170 277150 496226
rect 277218 496170 277274 496226
rect 277342 496170 277398 496226
rect 276970 496046 277026 496102
rect 277094 496046 277150 496102
rect 277218 496046 277274 496102
rect 277342 496046 277398 496102
rect 276970 495922 277026 495978
rect 277094 495922 277150 495978
rect 277218 495922 277274 495978
rect 277342 495922 277398 495978
rect 276970 478294 277026 478350
rect 277094 478294 277150 478350
rect 277218 478294 277274 478350
rect 277342 478294 277398 478350
rect 276970 478170 277026 478226
rect 277094 478170 277150 478226
rect 277218 478170 277274 478226
rect 277342 478170 277398 478226
rect 276970 478046 277026 478102
rect 277094 478046 277150 478102
rect 277218 478046 277274 478102
rect 277342 478046 277398 478102
rect 276970 477922 277026 477978
rect 277094 477922 277150 477978
rect 277218 477922 277274 477978
rect 277342 477922 277398 477978
rect 276970 460294 277026 460350
rect 277094 460294 277150 460350
rect 277218 460294 277274 460350
rect 277342 460294 277398 460350
rect 276970 460170 277026 460226
rect 277094 460170 277150 460226
rect 277218 460170 277274 460226
rect 277342 460170 277398 460226
rect 276970 460046 277026 460102
rect 277094 460046 277150 460102
rect 277218 460046 277274 460102
rect 277342 460046 277398 460102
rect 276970 459922 277026 459978
rect 277094 459922 277150 459978
rect 277218 459922 277274 459978
rect 277342 459922 277398 459978
rect 291250 597156 291306 597212
rect 291374 597156 291430 597212
rect 291498 597156 291554 597212
rect 291622 597156 291678 597212
rect 291250 597032 291306 597088
rect 291374 597032 291430 597088
rect 291498 597032 291554 597088
rect 291622 597032 291678 597088
rect 291250 596908 291306 596964
rect 291374 596908 291430 596964
rect 291498 596908 291554 596964
rect 291622 596908 291678 596964
rect 291250 596784 291306 596840
rect 291374 596784 291430 596840
rect 291498 596784 291554 596840
rect 291622 596784 291678 596840
rect 291250 580294 291306 580350
rect 291374 580294 291430 580350
rect 291498 580294 291554 580350
rect 291622 580294 291678 580350
rect 291250 580170 291306 580226
rect 291374 580170 291430 580226
rect 291498 580170 291554 580226
rect 291622 580170 291678 580226
rect 291250 580046 291306 580102
rect 291374 580046 291430 580102
rect 291498 580046 291554 580102
rect 291622 580046 291678 580102
rect 291250 579922 291306 579978
rect 291374 579922 291430 579978
rect 291498 579922 291554 579978
rect 291622 579922 291678 579978
rect 291250 562294 291306 562350
rect 291374 562294 291430 562350
rect 291498 562294 291554 562350
rect 291622 562294 291678 562350
rect 291250 562170 291306 562226
rect 291374 562170 291430 562226
rect 291498 562170 291554 562226
rect 291622 562170 291678 562226
rect 291250 562046 291306 562102
rect 291374 562046 291430 562102
rect 291498 562046 291554 562102
rect 291622 562046 291678 562102
rect 291250 561922 291306 561978
rect 291374 561922 291430 561978
rect 291498 561922 291554 561978
rect 291622 561922 291678 561978
rect 291250 544294 291306 544350
rect 291374 544294 291430 544350
rect 291498 544294 291554 544350
rect 291622 544294 291678 544350
rect 291250 544170 291306 544226
rect 291374 544170 291430 544226
rect 291498 544170 291554 544226
rect 291622 544170 291678 544226
rect 291250 544046 291306 544102
rect 291374 544046 291430 544102
rect 291498 544046 291554 544102
rect 291622 544046 291678 544102
rect 291250 543922 291306 543978
rect 291374 543922 291430 543978
rect 291498 543922 291554 543978
rect 291622 543922 291678 543978
rect 291250 526294 291306 526350
rect 291374 526294 291430 526350
rect 291498 526294 291554 526350
rect 291622 526294 291678 526350
rect 291250 526170 291306 526226
rect 291374 526170 291430 526226
rect 291498 526170 291554 526226
rect 291622 526170 291678 526226
rect 291250 526046 291306 526102
rect 291374 526046 291430 526102
rect 291498 526046 291554 526102
rect 291622 526046 291678 526102
rect 291250 525922 291306 525978
rect 291374 525922 291430 525978
rect 291498 525922 291554 525978
rect 291622 525922 291678 525978
rect 291250 508294 291306 508350
rect 291374 508294 291430 508350
rect 291498 508294 291554 508350
rect 291622 508294 291678 508350
rect 291250 508170 291306 508226
rect 291374 508170 291430 508226
rect 291498 508170 291554 508226
rect 291622 508170 291678 508226
rect 291250 508046 291306 508102
rect 291374 508046 291430 508102
rect 291498 508046 291554 508102
rect 291622 508046 291678 508102
rect 291250 507922 291306 507978
rect 291374 507922 291430 507978
rect 291498 507922 291554 507978
rect 291622 507922 291678 507978
rect 291250 490294 291306 490350
rect 291374 490294 291430 490350
rect 291498 490294 291554 490350
rect 291622 490294 291678 490350
rect 291250 490170 291306 490226
rect 291374 490170 291430 490226
rect 291498 490170 291554 490226
rect 291622 490170 291678 490226
rect 291250 490046 291306 490102
rect 291374 490046 291430 490102
rect 291498 490046 291554 490102
rect 291622 490046 291678 490102
rect 291250 489922 291306 489978
rect 291374 489922 291430 489978
rect 291498 489922 291554 489978
rect 291622 489922 291678 489978
rect 291250 472294 291306 472350
rect 291374 472294 291430 472350
rect 291498 472294 291554 472350
rect 291622 472294 291678 472350
rect 291250 472170 291306 472226
rect 291374 472170 291430 472226
rect 291498 472170 291554 472226
rect 291622 472170 291678 472226
rect 291250 472046 291306 472102
rect 291374 472046 291430 472102
rect 291498 472046 291554 472102
rect 291622 472046 291678 472102
rect 291250 471922 291306 471978
rect 291374 471922 291430 471978
rect 291498 471922 291554 471978
rect 291622 471922 291678 471978
rect 294970 598116 295026 598172
rect 295094 598116 295150 598172
rect 295218 598116 295274 598172
rect 295342 598116 295398 598172
rect 294970 597992 295026 598048
rect 295094 597992 295150 598048
rect 295218 597992 295274 598048
rect 295342 597992 295398 598048
rect 294970 597868 295026 597924
rect 295094 597868 295150 597924
rect 295218 597868 295274 597924
rect 295342 597868 295398 597924
rect 294970 597744 295026 597800
rect 295094 597744 295150 597800
rect 295218 597744 295274 597800
rect 295342 597744 295398 597800
rect 294970 586294 295026 586350
rect 295094 586294 295150 586350
rect 295218 586294 295274 586350
rect 295342 586294 295398 586350
rect 294970 586170 295026 586226
rect 295094 586170 295150 586226
rect 295218 586170 295274 586226
rect 295342 586170 295398 586226
rect 294970 586046 295026 586102
rect 295094 586046 295150 586102
rect 295218 586046 295274 586102
rect 295342 586046 295398 586102
rect 294970 585922 295026 585978
rect 295094 585922 295150 585978
rect 295218 585922 295274 585978
rect 295342 585922 295398 585978
rect 294970 568294 295026 568350
rect 295094 568294 295150 568350
rect 295218 568294 295274 568350
rect 295342 568294 295398 568350
rect 294970 568170 295026 568226
rect 295094 568170 295150 568226
rect 295218 568170 295274 568226
rect 295342 568170 295398 568226
rect 294970 568046 295026 568102
rect 295094 568046 295150 568102
rect 295218 568046 295274 568102
rect 295342 568046 295398 568102
rect 294970 567922 295026 567978
rect 295094 567922 295150 567978
rect 295218 567922 295274 567978
rect 295342 567922 295398 567978
rect 294970 550294 295026 550350
rect 295094 550294 295150 550350
rect 295218 550294 295274 550350
rect 295342 550294 295398 550350
rect 294970 550170 295026 550226
rect 295094 550170 295150 550226
rect 295218 550170 295274 550226
rect 295342 550170 295398 550226
rect 294970 550046 295026 550102
rect 295094 550046 295150 550102
rect 295218 550046 295274 550102
rect 295342 550046 295398 550102
rect 294970 549922 295026 549978
rect 295094 549922 295150 549978
rect 295218 549922 295274 549978
rect 295342 549922 295398 549978
rect 294970 532294 295026 532350
rect 295094 532294 295150 532350
rect 295218 532294 295274 532350
rect 295342 532294 295398 532350
rect 294970 532170 295026 532226
rect 295094 532170 295150 532226
rect 295218 532170 295274 532226
rect 295342 532170 295398 532226
rect 294970 532046 295026 532102
rect 295094 532046 295150 532102
rect 295218 532046 295274 532102
rect 295342 532046 295398 532102
rect 294970 531922 295026 531978
rect 295094 531922 295150 531978
rect 295218 531922 295274 531978
rect 295342 531922 295398 531978
rect 294970 514294 295026 514350
rect 295094 514294 295150 514350
rect 295218 514294 295274 514350
rect 295342 514294 295398 514350
rect 294970 514170 295026 514226
rect 295094 514170 295150 514226
rect 295218 514170 295274 514226
rect 295342 514170 295398 514226
rect 294970 514046 295026 514102
rect 295094 514046 295150 514102
rect 295218 514046 295274 514102
rect 295342 514046 295398 514102
rect 294970 513922 295026 513978
rect 295094 513922 295150 513978
rect 295218 513922 295274 513978
rect 295342 513922 295398 513978
rect 294970 496294 295026 496350
rect 295094 496294 295150 496350
rect 295218 496294 295274 496350
rect 295342 496294 295398 496350
rect 294970 496170 295026 496226
rect 295094 496170 295150 496226
rect 295218 496170 295274 496226
rect 295342 496170 295398 496226
rect 294970 496046 295026 496102
rect 295094 496046 295150 496102
rect 295218 496046 295274 496102
rect 295342 496046 295398 496102
rect 294970 495922 295026 495978
rect 295094 495922 295150 495978
rect 295218 495922 295274 495978
rect 295342 495922 295398 495978
rect 294970 478294 295026 478350
rect 295094 478294 295150 478350
rect 295218 478294 295274 478350
rect 295342 478294 295398 478350
rect 294970 478170 295026 478226
rect 295094 478170 295150 478226
rect 295218 478170 295274 478226
rect 295342 478170 295398 478226
rect 294970 478046 295026 478102
rect 295094 478046 295150 478102
rect 295218 478046 295274 478102
rect 295342 478046 295398 478102
rect 294970 477922 295026 477978
rect 295094 477922 295150 477978
rect 295218 477922 295274 477978
rect 295342 477922 295398 477978
rect 294970 460294 295026 460350
rect 295094 460294 295150 460350
rect 295218 460294 295274 460350
rect 295342 460294 295398 460350
rect 294970 460170 295026 460226
rect 295094 460170 295150 460226
rect 295218 460170 295274 460226
rect 295342 460170 295398 460226
rect 294970 460046 295026 460102
rect 295094 460046 295150 460102
rect 295218 460046 295274 460102
rect 295342 460046 295398 460102
rect 294970 459922 295026 459978
rect 295094 459922 295150 459978
rect 295218 459922 295274 459978
rect 295342 459922 295398 459978
rect 309250 597156 309306 597212
rect 309374 597156 309430 597212
rect 309498 597156 309554 597212
rect 309622 597156 309678 597212
rect 309250 597032 309306 597088
rect 309374 597032 309430 597088
rect 309498 597032 309554 597088
rect 309622 597032 309678 597088
rect 309250 596908 309306 596964
rect 309374 596908 309430 596964
rect 309498 596908 309554 596964
rect 309622 596908 309678 596964
rect 309250 596784 309306 596840
rect 309374 596784 309430 596840
rect 309498 596784 309554 596840
rect 309622 596784 309678 596840
rect 309250 580294 309306 580350
rect 309374 580294 309430 580350
rect 309498 580294 309554 580350
rect 309622 580294 309678 580350
rect 309250 580170 309306 580226
rect 309374 580170 309430 580226
rect 309498 580170 309554 580226
rect 309622 580170 309678 580226
rect 309250 580046 309306 580102
rect 309374 580046 309430 580102
rect 309498 580046 309554 580102
rect 309622 580046 309678 580102
rect 309250 579922 309306 579978
rect 309374 579922 309430 579978
rect 309498 579922 309554 579978
rect 309622 579922 309678 579978
rect 309250 562294 309306 562350
rect 309374 562294 309430 562350
rect 309498 562294 309554 562350
rect 309622 562294 309678 562350
rect 309250 562170 309306 562226
rect 309374 562170 309430 562226
rect 309498 562170 309554 562226
rect 309622 562170 309678 562226
rect 309250 562046 309306 562102
rect 309374 562046 309430 562102
rect 309498 562046 309554 562102
rect 309622 562046 309678 562102
rect 309250 561922 309306 561978
rect 309374 561922 309430 561978
rect 309498 561922 309554 561978
rect 309622 561922 309678 561978
rect 309250 544294 309306 544350
rect 309374 544294 309430 544350
rect 309498 544294 309554 544350
rect 309622 544294 309678 544350
rect 309250 544170 309306 544226
rect 309374 544170 309430 544226
rect 309498 544170 309554 544226
rect 309622 544170 309678 544226
rect 309250 544046 309306 544102
rect 309374 544046 309430 544102
rect 309498 544046 309554 544102
rect 309622 544046 309678 544102
rect 309250 543922 309306 543978
rect 309374 543922 309430 543978
rect 309498 543922 309554 543978
rect 309622 543922 309678 543978
rect 309250 526294 309306 526350
rect 309374 526294 309430 526350
rect 309498 526294 309554 526350
rect 309622 526294 309678 526350
rect 309250 526170 309306 526226
rect 309374 526170 309430 526226
rect 309498 526170 309554 526226
rect 309622 526170 309678 526226
rect 309250 526046 309306 526102
rect 309374 526046 309430 526102
rect 309498 526046 309554 526102
rect 309622 526046 309678 526102
rect 309250 525922 309306 525978
rect 309374 525922 309430 525978
rect 309498 525922 309554 525978
rect 309622 525922 309678 525978
rect 309250 508294 309306 508350
rect 309374 508294 309430 508350
rect 309498 508294 309554 508350
rect 309622 508294 309678 508350
rect 309250 508170 309306 508226
rect 309374 508170 309430 508226
rect 309498 508170 309554 508226
rect 309622 508170 309678 508226
rect 309250 508046 309306 508102
rect 309374 508046 309430 508102
rect 309498 508046 309554 508102
rect 309622 508046 309678 508102
rect 309250 507922 309306 507978
rect 309374 507922 309430 507978
rect 309498 507922 309554 507978
rect 309622 507922 309678 507978
rect 309250 490294 309306 490350
rect 309374 490294 309430 490350
rect 309498 490294 309554 490350
rect 309622 490294 309678 490350
rect 309250 490170 309306 490226
rect 309374 490170 309430 490226
rect 309498 490170 309554 490226
rect 309622 490170 309678 490226
rect 309250 490046 309306 490102
rect 309374 490046 309430 490102
rect 309498 490046 309554 490102
rect 309622 490046 309678 490102
rect 309250 489922 309306 489978
rect 309374 489922 309430 489978
rect 309498 489922 309554 489978
rect 309622 489922 309678 489978
rect 309250 472294 309306 472350
rect 309374 472294 309430 472350
rect 309498 472294 309554 472350
rect 309622 472294 309678 472350
rect 309250 472170 309306 472226
rect 309374 472170 309430 472226
rect 309498 472170 309554 472226
rect 309622 472170 309678 472226
rect 309250 472046 309306 472102
rect 309374 472046 309430 472102
rect 309498 472046 309554 472102
rect 309622 472046 309678 472102
rect 309250 471922 309306 471978
rect 309374 471922 309430 471978
rect 309498 471922 309554 471978
rect 309622 471922 309678 471978
rect 312970 598116 313026 598172
rect 313094 598116 313150 598172
rect 313218 598116 313274 598172
rect 313342 598116 313398 598172
rect 312970 597992 313026 598048
rect 313094 597992 313150 598048
rect 313218 597992 313274 598048
rect 313342 597992 313398 598048
rect 312970 597868 313026 597924
rect 313094 597868 313150 597924
rect 313218 597868 313274 597924
rect 313342 597868 313398 597924
rect 312970 597744 313026 597800
rect 313094 597744 313150 597800
rect 313218 597744 313274 597800
rect 313342 597744 313398 597800
rect 312970 586294 313026 586350
rect 313094 586294 313150 586350
rect 313218 586294 313274 586350
rect 313342 586294 313398 586350
rect 312970 586170 313026 586226
rect 313094 586170 313150 586226
rect 313218 586170 313274 586226
rect 313342 586170 313398 586226
rect 312970 586046 313026 586102
rect 313094 586046 313150 586102
rect 313218 586046 313274 586102
rect 313342 586046 313398 586102
rect 312970 585922 313026 585978
rect 313094 585922 313150 585978
rect 313218 585922 313274 585978
rect 313342 585922 313398 585978
rect 312970 568294 313026 568350
rect 313094 568294 313150 568350
rect 313218 568294 313274 568350
rect 313342 568294 313398 568350
rect 312970 568170 313026 568226
rect 313094 568170 313150 568226
rect 313218 568170 313274 568226
rect 313342 568170 313398 568226
rect 312970 568046 313026 568102
rect 313094 568046 313150 568102
rect 313218 568046 313274 568102
rect 313342 568046 313398 568102
rect 312970 567922 313026 567978
rect 313094 567922 313150 567978
rect 313218 567922 313274 567978
rect 313342 567922 313398 567978
rect 312970 550294 313026 550350
rect 313094 550294 313150 550350
rect 313218 550294 313274 550350
rect 313342 550294 313398 550350
rect 312970 550170 313026 550226
rect 313094 550170 313150 550226
rect 313218 550170 313274 550226
rect 313342 550170 313398 550226
rect 312970 550046 313026 550102
rect 313094 550046 313150 550102
rect 313218 550046 313274 550102
rect 313342 550046 313398 550102
rect 312970 549922 313026 549978
rect 313094 549922 313150 549978
rect 313218 549922 313274 549978
rect 313342 549922 313398 549978
rect 312970 532294 313026 532350
rect 313094 532294 313150 532350
rect 313218 532294 313274 532350
rect 313342 532294 313398 532350
rect 312970 532170 313026 532226
rect 313094 532170 313150 532226
rect 313218 532170 313274 532226
rect 313342 532170 313398 532226
rect 312970 532046 313026 532102
rect 313094 532046 313150 532102
rect 313218 532046 313274 532102
rect 313342 532046 313398 532102
rect 312970 531922 313026 531978
rect 313094 531922 313150 531978
rect 313218 531922 313274 531978
rect 313342 531922 313398 531978
rect 312970 514294 313026 514350
rect 313094 514294 313150 514350
rect 313218 514294 313274 514350
rect 313342 514294 313398 514350
rect 312970 514170 313026 514226
rect 313094 514170 313150 514226
rect 313218 514170 313274 514226
rect 313342 514170 313398 514226
rect 312970 514046 313026 514102
rect 313094 514046 313150 514102
rect 313218 514046 313274 514102
rect 313342 514046 313398 514102
rect 312970 513922 313026 513978
rect 313094 513922 313150 513978
rect 313218 513922 313274 513978
rect 313342 513922 313398 513978
rect 312970 496294 313026 496350
rect 313094 496294 313150 496350
rect 313218 496294 313274 496350
rect 313342 496294 313398 496350
rect 312970 496170 313026 496226
rect 313094 496170 313150 496226
rect 313218 496170 313274 496226
rect 313342 496170 313398 496226
rect 312970 496046 313026 496102
rect 313094 496046 313150 496102
rect 313218 496046 313274 496102
rect 313342 496046 313398 496102
rect 312970 495922 313026 495978
rect 313094 495922 313150 495978
rect 313218 495922 313274 495978
rect 313342 495922 313398 495978
rect 312970 478294 313026 478350
rect 313094 478294 313150 478350
rect 313218 478294 313274 478350
rect 313342 478294 313398 478350
rect 312970 478170 313026 478226
rect 313094 478170 313150 478226
rect 313218 478170 313274 478226
rect 313342 478170 313398 478226
rect 312970 478046 313026 478102
rect 313094 478046 313150 478102
rect 313218 478046 313274 478102
rect 313342 478046 313398 478102
rect 312970 477922 313026 477978
rect 313094 477922 313150 477978
rect 313218 477922 313274 477978
rect 313342 477922 313398 477978
rect 312970 460294 313026 460350
rect 313094 460294 313150 460350
rect 313218 460294 313274 460350
rect 313342 460294 313398 460350
rect 312970 460170 313026 460226
rect 313094 460170 313150 460226
rect 313218 460170 313274 460226
rect 313342 460170 313398 460226
rect 312970 460046 313026 460102
rect 313094 460046 313150 460102
rect 313218 460046 313274 460102
rect 313342 460046 313398 460102
rect 312970 459922 313026 459978
rect 313094 459922 313150 459978
rect 313218 459922 313274 459978
rect 313342 459922 313398 459978
rect 327250 597156 327306 597212
rect 327374 597156 327430 597212
rect 327498 597156 327554 597212
rect 327622 597156 327678 597212
rect 327250 597032 327306 597088
rect 327374 597032 327430 597088
rect 327498 597032 327554 597088
rect 327622 597032 327678 597088
rect 327250 596908 327306 596964
rect 327374 596908 327430 596964
rect 327498 596908 327554 596964
rect 327622 596908 327678 596964
rect 327250 596784 327306 596840
rect 327374 596784 327430 596840
rect 327498 596784 327554 596840
rect 327622 596784 327678 596840
rect 327250 580294 327306 580350
rect 327374 580294 327430 580350
rect 327498 580294 327554 580350
rect 327622 580294 327678 580350
rect 327250 580170 327306 580226
rect 327374 580170 327430 580226
rect 327498 580170 327554 580226
rect 327622 580170 327678 580226
rect 327250 580046 327306 580102
rect 327374 580046 327430 580102
rect 327498 580046 327554 580102
rect 327622 580046 327678 580102
rect 327250 579922 327306 579978
rect 327374 579922 327430 579978
rect 327498 579922 327554 579978
rect 327622 579922 327678 579978
rect 327250 562294 327306 562350
rect 327374 562294 327430 562350
rect 327498 562294 327554 562350
rect 327622 562294 327678 562350
rect 327250 562170 327306 562226
rect 327374 562170 327430 562226
rect 327498 562170 327554 562226
rect 327622 562170 327678 562226
rect 327250 562046 327306 562102
rect 327374 562046 327430 562102
rect 327498 562046 327554 562102
rect 327622 562046 327678 562102
rect 327250 561922 327306 561978
rect 327374 561922 327430 561978
rect 327498 561922 327554 561978
rect 327622 561922 327678 561978
rect 327250 544294 327306 544350
rect 327374 544294 327430 544350
rect 327498 544294 327554 544350
rect 327622 544294 327678 544350
rect 327250 544170 327306 544226
rect 327374 544170 327430 544226
rect 327498 544170 327554 544226
rect 327622 544170 327678 544226
rect 327250 544046 327306 544102
rect 327374 544046 327430 544102
rect 327498 544046 327554 544102
rect 327622 544046 327678 544102
rect 327250 543922 327306 543978
rect 327374 543922 327430 543978
rect 327498 543922 327554 543978
rect 327622 543922 327678 543978
rect 327250 526294 327306 526350
rect 327374 526294 327430 526350
rect 327498 526294 327554 526350
rect 327622 526294 327678 526350
rect 327250 526170 327306 526226
rect 327374 526170 327430 526226
rect 327498 526170 327554 526226
rect 327622 526170 327678 526226
rect 327250 526046 327306 526102
rect 327374 526046 327430 526102
rect 327498 526046 327554 526102
rect 327622 526046 327678 526102
rect 327250 525922 327306 525978
rect 327374 525922 327430 525978
rect 327498 525922 327554 525978
rect 327622 525922 327678 525978
rect 327250 508294 327306 508350
rect 327374 508294 327430 508350
rect 327498 508294 327554 508350
rect 327622 508294 327678 508350
rect 327250 508170 327306 508226
rect 327374 508170 327430 508226
rect 327498 508170 327554 508226
rect 327622 508170 327678 508226
rect 327250 508046 327306 508102
rect 327374 508046 327430 508102
rect 327498 508046 327554 508102
rect 327622 508046 327678 508102
rect 327250 507922 327306 507978
rect 327374 507922 327430 507978
rect 327498 507922 327554 507978
rect 327622 507922 327678 507978
rect 327250 490294 327306 490350
rect 327374 490294 327430 490350
rect 327498 490294 327554 490350
rect 327622 490294 327678 490350
rect 327250 490170 327306 490226
rect 327374 490170 327430 490226
rect 327498 490170 327554 490226
rect 327622 490170 327678 490226
rect 327250 490046 327306 490102
rect 327374 490046 327430 490102
rect 327498 490046 327554 490102
rect 327622 490046 327678 490102
rect 327250 489922 327306 489978
rect 327374 489922 327430 489978
rect 327498 489922 327554 489978
rect 327622 489922 327678 489978
rect 327250 472294 327306 472350
rect 327374 472294 327430 472350
rect 327498 472294 327554 472350
rect 327622 472294 327678 472350
rect 327250 472170 327306 472226
rect 327374 472170 327430 472226
rect 327498 472170 327554 472226
rect 327622 472170 327678 472226
rect 327250 472046 327306 472102
rect 327374 472046 327430 472102
rect 327498 472046 327554 472102
rect 327622 472046 327678 472102
rect 327250 471922 327306 471978
rect 327374 471922 327430 471978
rect 327498 471922 327554 471978
rect 327622 471922 327678 471978
rect 330970 598116 331026 598172
rect 331094 598116 331150 598172
rect 331218 598116 331274 598172
rect 331342 598116 331398 598172
rect 330970 597992 331026 598048
rect 331094 597992 331150 598048
rect 331218 597992 331274 598048
rect 331342 597992 331398 598048
rect 330970 597868 331026 597924
rect 331094 597868 331150 597924
rect 331218 597868 331274 597924
rect 331342 597868 331398 597924
rect 330970 597744 331026 597800
rect 331094 597744 331150 597800
rect 331218 597744 331274 597800
rect 331342 597744 331398 597800
rect 330970 586294 331026 586350
rect 331094 586294 331150 586350
rect 331218 586294 331274 586350
rect 331342 586294 331398 586350
rect 330970 586170 331026 586226
rect 331094 586170 331150 586226
rect 331218 586170 331274 586226
rect 331342 586170 331398 586226
rect 330970 586046 331026 586102
rect 331094 586046 331150 586102
rect 331218 586046 331274 586102
rect 331342 586046 331398 586102
rect 330970 585922 331026 585978
rect 331094 585922 331150 585978
rect 331218 585922 331274 585978
rect 331342 585922 331398 585978
rect 330970 568294 331026 568350
rect 331094 568294 331150 568350
rect 331218 568294 331274 568350
rect 331342 568294 331398 568350
rect 330970 568170 331026 568226
rect 331094 568170 331150 568226
rect 331218 568170 331274 568226
rect 331342 568170 331398 568226
rect 330970 568046 331026 568102
rect 331094 568046 331150 568102
rect 331218 568046 331274 568102
rect 331342 568046 331398 568102
rect 330970 567922 331026 567978
rect 331094 567922 331150 567978
rect 331218 567922 331274 567978
rect 331342 567922 331398 567978
rect 330970 550294 331026 550350
rect 331094 550294 331150 550350
rect 331218 550294 331274 550350
rect 331342 550294 331398 550350
rect 330970 550170 331026 550226
rect 331094 550170 331150 550226
rect 331218 550170 331274 550226
rect 331342 550170 331398 550226
rect 330970 550046 331026 550102
rect 331094 550046 331150 550102
rect 331218 550046 331274 550102
rect 331342 550046 331398 550102
rect 330970 549922 331026 549978
rect 331094 549922 331150 549978
rect 331218 549922 331274 549978
rect 331342 549922 331398 549978
rect 330970 532294 331026 532350
rect 331094 532294 331150 532350
rect 331218 532294 331274 532350
rect 331342 532294 331398 532350
rect 330970 532170 331026 532226
rect 331094 532170 331150 532226
rect 331218 532170 331274 532226
rect 331342 532170 331398 532226
rect 330970 532046 331026 532102
rect 331094 532046 331150 532102
rect 331218 532046 331274 532102
rect 331342 532046 331398 532102
rect 330970 531922 331026 531978
rect 331094 531922 331150 531978
rect 331218 531922 331274 531978
rect 331342 531922 331398 531978
rect 330970 514294 331026 514350
rect 331094 514294 331150 514350
rect 331218 514294 331274 514350
rect 331342 514294 331398 514350
rect 330970 514170 331026 514226
rect 331094 514170 331150 514226
rect 331218 514170 331274 514226
rect 331342 514170 331398 514226
rect 330970 514046 331026 514102
rect 331094 514046 331150 514102
rect 331218 514046 331274 514102
rect 331342 514046 331398 514102
rect 330970 513922 331026 513978
rect 331094 513922 331150 513978
rect 331218 513922 331274 513978
rect 331342 513922 331398 513978
rect 330970 496294 331026 496350
rect 331094 496294 331150 496350
rect 331218 496294 331274 496350
rect 331342 496294 331398 496350
rect 330970 496170 331026 496226
rect 331094 496170 331150 496226
rect 331218 496170 331274 496226
rect 331342 496170 331398 496226
rect 330970 496046 331026 496102
rect 331094 496046 331150 496102
rect 331218 496046 331274 496102
rect 331342 496046 331398 496102
rect 330970 495922 331026 495978
rect 331094 495922 331150 495978
rect 331218 495922 331274 495978
rect 331342 495922 331398 495978
rect 330970 478294 331026 478350
rect 331094 478294 331150 478350
rect 331218 478294 331274 478350
rect 331342 478294 331398 478350
rect 330970 478170 331026 478226
rect 331094 478170 331150 478226
rect 331218 478170 331274 478226
rect 331342 478170 331398 478226
rect 330970 478046 331026 478102
rect 331094 478046 331150 478102
rect 331218 478046 331274 478102
rect 331342 478046 331398 478102
rect 330970 477922 331026 477978
rect 331094 477922 331150 477978
rect 331218 477922 331274 477978
rect 331342 477922 331398 477978
rect 330970 460294 331026 460350
rect 331094 460294 331150 460350
rect 331218 460294 331274 460350
rect 331342 460294 331398 460350
rect 330970 460170 331026 460226
rect 331094 460170 331150 460226
rect 331218 460170 331274 460226
rect 331342 460170 331398 460226
rect 330970 460046 331026 460102
rect 331094 460046 331150 460102
rect 331218 460046 331274 460102
rect 331342 460046 331398 460102
rect 330970 459922 331026 459978
rect 331094 459922 331150 459978
rect 331218 459922 331274 459978
rect 331342 459922 331398 459978
rect 345250 597156 345306 597212
rect 345374 597156 345430 597212
rect 345498 597156 345554 597212
rect 345622 597156 345678 597212
rect 345250 597032 345306 597088
rect 345374 597032 345430 597088
rect 345498 597032 345554 597088
rect 345622 597032 345678 597088
rect 345250 596908 345306 596964
rect 345374 596908 345430 596964
rect 345498 596908 345554 596964
rect 345622 596908 345678 596964
rect 345250 596784 345306 596840
rect 345374 596784 345430 596840
rect 345498 596784 345554 596840
rect 345622 596784 345678 596840
rect 345250 580294 345306 580350
rect 345374 580294 345430 580350
rect 345498 580294 345554 580350
rect 345622 580294 345678 580350
rect 345250 580170 345306 580226
rect 345374 580170 345430 580226
rect 345498 580170 345554 580226
rect 345622 580170 345678 580226
rect 345250 580046 345306 580102
rect 345374 580046 345430 580102
rect 345498 580046 345554 580102
rect 345622 580046 345678 580102
rect 345250 579922 345306 579978
rect 345374 579922 345430 579978
rect 345498 579922 345554 579978
rect 345622 579922 345678 579978
rect 345250 562294 345306 562350
rect 345374 562294 345430 562350
rect 345498 562294 345554 562350
rect 345622 562294 345678 562350
rect 345250 562170 345306 562226
rect 345374 562170 345430 562226
rect 345498 562170 345554 562226
rect 345622 562170 345678 562226
rect 345250 562046 345306 562102
rect 345374 562046 345430 562102
rect 345498 562046 345554 562102
rect 345622 562046 345678 562102
rect 345250 561922 345306 561978
rect 345374 561922 345430 561978
rect 345498 561922 345554 561978
rect 345622 561922 345678 561978
rect 345250 544294 345306 544350
rect 345374 544294 345430 544350
rect 345498 544294 345554 544350
rect 345622 544294 345678 544350
rect 345250 544170 345306 544226
rect 345374 544170 345430 544226
rect 345498 544170 345554 544226
rect 345622 544170 345678 544226
rect 345250 544046 345306 544102
rect 345374 544046 345430 544102
rect 345498 544046 345554 544102
rect 345622 544046 345678 544102
rect 345250 543922 345306 543978
rect 345374 543922 345430 543978
rect 345498 543922 345554 543978
rect 345622 543922 345678 543978
rect 345250 526294 345306 526350
rect 345374 526294 345430 526350
rect 345498 526294 345554 526350
rect 345622 526294 345678 526350
rect 345250 526170 345306 526226
rect 345374 526170 345430 526226
rect 345498 526170 345554 526226
rect 345622 526170 345678 526226
rect 345250 526046 345306 526102
rect 345374 526046 345430 526102
rect 345498 526046 345554 526102
rect 345622 526046 345678 526102
rect 345250 525922 345306 525978
rect 345374 525922 345430 525978
rect 345498 525922 345554 525978
rect 345622 525922 345678 525978
rect 345250 508294 345306 508350
rect 345374 508294 345430 508350
rect 345498 508294 345554 508350
rect 345622 508294 345678 508350
rect 345250 508170 345306 508226
rect 345374 508170 345430 508226
rect 345498 508170 345554 508226
rect 345622 508170 345678 508226
rect 345250 508046 345306 508102
rect 345374 508046 345430 508102
rect 345498 508046 345554 508102
rect 345622 508046 345678 508102
rect 345250 507922 345306 507978
rect 345374 507922 345430 507978
rect 345498 507922 345554 507978
rect 345622 507922 345678 507978
rect 345250 490294 345306 490350
rect 345374 490294 345430 490350
rect 345498 490294 345554 490350
rect 345622 490294 345678 490350
rect 345250 490170 345306 490226
rect 345374 490170 345430 490226
rect 345498 490170 345554 490226
rect 345622 490170 345678 490226
rect 345250 490046 345306 490102
rect 345374 490046 345430 490102
rect 345498 490046 345554 490102
rect 345622 490046 345678 490102
rect 345250 489922 345306 489978
rect 345374 489922 345430 489978
rect 345498 489922 345554 489978
rect 345622 489922 345678 489978
rect 345250 472294 345306 472350
rect 345374 472294 345430 472350
rect 345498 472294 345554 472350
rect 345622 472294 345678 472350
rect 345250 472170 345306 472226
rect 345374 472170 345430 472226
rect 345498 472170 345554 472226
rect 345622 472170 345678 472226
rect 345250 472046 345306 472102
rect 345374 472046 345430 472102
rect 345498 472046 345554 472102
rect 345622 472046 345678 472102
rect 345250 471922 345306 471978
rect 345374 471922 345430 471978
rect 345498 471922 345554 471978
rect 345622 471922 345678 471978
rect 348970 598116 349026 598172
rect 349094 598116 349150 598172
rect 349218 598116 349274 598172
rect 349342 598116 349398 598172
rect 348970 597992 349026 598048
rect 349094 597992 349150 598048
rect 349218 597992 349274 598048
rect 349342 597992 349398 598048
rect 348970 597868 349026 597924
rect 349094 597868 349150 597924
rect 349218 597868 349274 597924
rect 349342 597868 349398 597924
rect 348970 597744 349026 597800
rect 349094 597744 349150 597800
rect 349218 597744 349274 597800
rect 349342 597744 349398 597800
rect 348970 586294 349026 586350
rect 349094 586294 349150 586350
rect 349218 586294 349274 586350
rect 349342 586294 349398 586350
rect 348970 586170 349026 586226
rect 349094 586170 349150 586226
rect 349218 586170 349274 586226
rect 349342 586170 349398 586226
rect 348970 586046 349026 586102
rect 349094 586046 349150 586102
rect 349218 586046 349274 586102
rect 349342 586046 349398 586102
rect 348970 585922 349026 585978
rect 349094 585922 349150 585978
rect 349218 585922 349274 585978
rect 349342 585922 349398 585978
rect 348970 568294 349026 568350
rect 349094 568294 349150 568350
rect 349218 568294 349274 568350
rect 349342 568294 349398 568350
rect 348970 568170 349026 568226
rect 349094 568170 349150 568226
rect 349218 568170 349274 568226
rect 349342 568170 349398 568226
rect 348970 568046 349026 568102
rect 349094 568046 349150 568102
rect 349218 568046 349274 568102
rect 349342 568046 349398 568102
rect 348970 567922 349026 567978
rect 349094 567922 349150 567978
rect 349218 567922 349274 567978
rect 349342 567922 349398 567978
rect 348970 550294 349026 550350
rect 349094 550294 349150 550350
rect 349218 550294 349274 550350
rect 349342 550294 349398 550350
rect 348970 550170 349026 550226
rect 349094 550170 349150 550226
rect 349218 550170 349274 550226
rect 349342 550170 349398 550226
rect 348970 550046 349026 550102
rect 349094 550046 349150 550102
rect 349218 550046 349274 550102
rect 349342 550046 349398 550102
rect 348970 549922 349026 549978
rect 349094 549922 349150 549978
rect 349218 549922 349274 549978
rect 349342 549922 349398 549978
rect 348970 532294 349026 532350
rect 349094 532294 349150 532350
rect 349218 532294 349274 532350
rect 349342 532294 349398 532350
rect 348970 532170 349026 532226
rect 349094 532170 349150 532226
rect 349218 532170 349274 532226
rect 349342 532170 349398 532226
rect 348970 532046 349026 532102
rect 349094 532046 349150 532102
rect 349218 532046 349274 532102
rect 349342 532046 349398 532102
rect 348970 531922 349026 531978
rect 349094 531922 349150 531978
rect 349218 531922 349274 531978
rect 349342 531922 349398 531978
rect 348970 514294 349026 514350
rect 349094 514294 349150 514350
rect 349218 514294 349274 514350
rect 349342 514294 349398 514350
rect 348970 514170 349026 514226
rect 349094 514170 349150 514226
rect 349218 514170 349274 514226
rect 349342 514170 349398 514226
rect 348970 514046 349026 514102
rect 349094 514046 349150 514102
rect 349218 514046 349274 514102
rect 349342 514046 349398 514102
rect 348970 513922 349026 513978
rect 349094 513922 349150 513978
rect 349218 513922 349274 513978
rect 349342 513922 349398 513978
rect 348970 496294 349026 496350
rect 349094 496294 349150 496350
rect 349218 496294 349274 496350
rect 349342 496294 349398 496350
rect 348970 496170 349026 496226
rect 349094 496170 349150 496226
rect 349218 496170 349274 496226
rect 349342 496170 349398 496226
rect 348970 496046 349026 496102
rect 349094 496046 349150 496102
rect 349218 496046 349274 496102
rect 349342 496046 349398 496102
rect 348970 495922 349026 495978
rect 349094 495922 349150 495978
rect 349218 495922 349274 495978
rect 349342 495922 349398 495978
rect 348970 478294 349026 478350
rect 349094 478294 349150 478350
rect 349218 478294 349274 478350
rect 349342 478294 349398 478350
rect 348970 478170 349026 478226
rect 349094 478170 349150 478226
rect 349218 478170 349274 478226
rect 349342 478170 349398 478226
rect 348970 478046 349026 478102
rect 349094 478046 349150 478102
rect 349218 478046 349274 478102
rect 349342 478046 349398 478102
rect 348970 477922 349026 477978
rect 349094 477922 349150 477978
rect 349218 477922 349274 477978
rect 349342 477922 349398 477978
rect 348970 460294 349026 460350
rect 349094 460294 349150 460350
rect 349218 460294 349274 460350
rect 349342 460294 349398 460350
rect 348970 460170 349026 460226
rect 349094 460170 349150 460226
rect 349218 460170 349274 460226
rect 349342 460170 349398 460226
rect 348970 460046 349026 460102
rect 349094 460046 349150 460102
rect 349218 460046 349274 460102
rect 349342 460046 349398 460102
rect 348970 459922 349026 459978
rect 349094 459922 349150 459978
rect 349218 459922 349274 459978
rect 349342 459922 349398 459978
rect 363250 597156 363306 597212
rect 363374 597156 363430 597212
rect 363498 597156 363554 597212
rect 363622 597156 363678 597212
rect 363250 597032 363306 597088
rect 363374 597032 363430 597088
rect 363498 597032 363554 597088
rect 363622 597032 363678 597088
rect 363250 596908 363306 596964
rect 363374 596908 363430 596964
rect 363498 596908 363554 596964
rect 363622 596908 363678 596964
rect 363250 596784 363306 596840
rect 363374 596784 363430 596840
rect 363498 596784 363554 596840
rect 363622 596784 363678 596840
rect 363250 580294 363306 580350
rect 363374 580294 363430 580350
rect 363498 580294 363554 580350
rect 363622 580294 363678 580350
rect 363250 580170 363306 580226
rect 363374 580170 363430 580226
rect 363498 580170 363554 580226
rect 363622 580170 363678 580226
rect 363250 580046 363306 580102
rect 363374 580046 363430 580102
rect 363498 580046 363554 580102
rect 363622 580046 363678 580102
rect 363250 579922 363306 579978
rect 363374 579922 363430 579978
rect 363498 579922 363554 579978
rect 363622 579922 363678 579978
rect 363250 562294 363306 562350
rect 363374 562294 363430 562350
rect 363498 562294 363554 562350
rect 363622 562294 363678 562350
rect 363250 562170 363306 562226
rect 363374 562170 363430 562226
rect 363498 562170 363554 562226
rect 363622 562170 363678 562226
rect 363250 562046 363306 562102
rect 363374 562046 363430 562102
rect 363498 562046 363554 562102
rect 363622 562046 363678 562102
rect 363250 561922 363306 561978
rect 363374 561922 363430 561978
rect 363498 561922 363554 561978
rect 363622 561922 363678 561978
rect 363250 544294 363306 544350
rect 363374 544294 363430 544350
rect 363498 544294 363554 544350
rect 363622 544294 363678 544350
rect 363250 544170 363306 544226
rect 363374 544170 363430 544226
rect 363498 544170 363554 544226
rect 363622 544170 363678 544226
rect 363250 544046 363306 544102
rect 363374 544046 363430 544102
rect 363498 544046 363554 544102
rect 363622 544046 363678 544102
rect 363250 543922 363306 543978
rect 363374 543922 363430 543978
rect 363498 543922 363554 543978
rect 363622 543922 363678 543978
rect 363250 526294 363306 526350
rect 363374 526294 363430 526350
rect 363498 526294 363554 526350
rect 363622 526294 363678 526350
rect 363250 526170 363306 526226
rect 363374 526170 363430 526226
rect 363498 526170 363554 526226
rect 363622 526170 363678 526226
rect 363250 526046 363306 526102
rect 363374 526046 363430 526102
rect 363498 526046 363554 526102
rect 363622 526046 363678 526102
rect 363250 525922 363306 525978
rect 363374 525922 363430 525978
rect 363498 525922 363554 525978
rect 363622 525922 363678 525978
rect 363250 508294 363306 508350
rect 363374 508294 363430 508350
rect 363498 508294 363554 508350
rect 363622 508294 363678 508350
rect 363250 508170 363306 508226
rect 363374 508170 363430 508226
rect 363498 508170 363554 508226
rect 363622 508170 363678 508226
rect 363250 508046 363306 508102
rect 363374 508046 363430 508102
rect 363498 508046 363554 508102
rect 363622 508046 363678 508102
rect 363250 507922 363306 507978
rect 363374 507922 363430 507978
rect 363498 507922 363554 507978
rect 363622 507922 363678 507978
rect 363250 490294 363306 490350
rect 363374 490294 363430 490350
rect 363498 490294 363554 490350
rect 363622 490294 363678 490350
rect 363250 490170 363306 490226
rect 363374 490170 363430 490226
rect 363498 490170 363554 490226
rect 363622 490170 363678 490226
rect 363250 490046 363306 490102
rect 363374 490046 363430 490102
rect 363498 490046 363554 490102
rect 363622 490046 363678 490102
rect 363250 489922 363306 489978
rect 363374 489922 363430 489978
rect 363498 489922 363554 489978
rect 363622 489922 363678 489978
rect 363250 472294 363306 472350
rect 363374 472294 363430 472350
rect 363498 472294 363554 472350
rect 363622 472294 363678 472350
rect 363250 472170 363306 472226
rect 363374 472170 363430 472226
rect 363498 472170 363554 472226
rect 363622 472170 363678 472226
rect 363250 472046 363306 472102
rect 363374 472046 363430 472102
rect 363498 472046 363554 472102
rect 363622 472046 363678 472102
rect 363250 471922 363306 471978
rect 363374 471922 363430 471978
rect 363498 471922 363554 471978
rect 363622 471922 363678 471978
rect 366970 598116 367026 598172
rect 367094 598116 367150 598172
rect 367218 598116 367274 598172
rect 367342 598116 367398 598172
rect 366970 597992 367026 598048
rect 367094 597992 367150 598048
rect 367218 597992 367274 598048
rect 367342 597992 367398 598048
rect 366970 597868 367026 597924
rect 367094 597868 367150 597924
rect 367218 597868 367274 597924
rect 367342 597868 367398 597924
rect 366970 597744 367026 597800
rect 367094 597744 367150 597800
rect 367218 597744 367274 597800
rect 367342 597744 367398 597800
rect 366970 586294 367026 586350
rect 367094 586294 367150 586350
rect 367218 586294 367274 586350
rect 367342 586294 367398 586350
rect 366970 586170 367026 586226
rect 367094 586170 367150 586226
rect 367218 586170 367274 586226
rect 367342 586170 367398 586226
rect 366970 586046 367026 586102
rect 367094 586046 367150 586102
rect 367218 586046 367274 586102
rect 367342 586046 367398 586102
rect 366970 585922 367026 585978
rect 367094 585922 367150 585978
rect 367218 585922 367274 585978
rect 367342 585922 367398 585978
rect 366970 568294 367026 568350
rect 367094 568294 367150 568350
rect 367218 568294 367274 568350
rect 367342 568294 367398 568350
rect 366970 568170 367026 568226
rect 367094 568170 367150 568226
rect 367218 568170 367274 568226
rect 367342 568170 367398 568226
rect 366970 568046 367026 568102
rect 367094 568046 367150 568102
rect 367218 568046 367274 568102
rect 367342 568046 367398 568102
rect 366970 567922 367026 567978
rect 367094 567922 367150 567978
rect 367218 567922 367274 567978
rect 367342 567922 367398 567978
rect 366970 550294 367026 550350
rect 367094 550294 367150 550350
rect 367218 550294 367274 550350
rect 367342 550294 367398 550350
rect 366970 550170 367026 550226
rect 367094 550170 367150 550226
rect 367218 550170 367274 550226
rect 367342 550170 367398 550226
rect 366970 550046 367026 550102
rect 367094 550046 367150 550102
rect 367218 550046 367274 550102
rect 367342 550046 367398 550102
rect 366970 549922 367026 549978
rect 367094 549922 367150 549978
rect 367218 549922 367274 549978
rect 367342 549922 367398 549978
rect 366970 532294 367026 532350
rect 367094 532294 367150 532350
rect 367218 532294 367274 532350
rect 367342 532294 367398 532350
rect 366970 532170 367026 532226
rect 367094 532170 367150 532226
rect 367218 532170 367274 532226
rect 367342 532170 367398 532226
rect 366970 532046 367026 532102
rect 367094 532046 367150 532102
rect 367218 532046 367274 532102
rect 367342 532046 367398 532102
rect 366970 531922 367026 531978
rect 367094 531922 367150 531978
rect 367218 531922 367274 531978
rect 367342 531922 367398 531978
rect 366970 514294 367026 514350
rect 367094 514294 367150 514350
rect 367218 514294 367274 514350
rect 367342 514294 367398 514350
rect 366970 514170 367026 514226
rect 367094 514170 367150 514226
rect 367218 514170 367274 514226
rect 367342 514170 367398 514226
rect 366970 514046 367026 514102
rect 367094 514046 367150 514102
rect 367218 514046 367274 514102
rect 367342 514046 367398 514102
rect 366970 513922 367026 513978
rect 367094 513922 367150 513978
rect 367218 513922 367274 513978
rect 367342 513922 367398 513978
rect 366970 496294 367026 496350
rect 367094 496294 367150 496350
rect 367218 496294 367274 496350
rect 367342 496294 367398 496350
rect 366970 496170 367026 496226
rect 367094 496170 367150 496226
rect 367218 496170 367274 496226
rect 367342 496170 367398 496226
rect 366970 496046 367026 496102
rect 367094 496046 367150 496102
rect 367218 496046 367274 496102
rect 367342 496046 367398 496102
rect 366970 495922 367026 495978
rect 367094 495922 367150 495978
rect 367218 495922 367274 495978
rect 367342 495922 367398 495978
rect 366970 478294 367026 478350
rect 367094 478294 367150 478350
rect 367218 478294 367274 478350
rect 367342 478294 367398 478350
rect 366970 478170 367026 478226
rect 367094 478170 367150 478226
rect 367218 478170 367274 478226
rect 367342 478170 367398 478226
rect 366970 478046 367026 478102
rect 367094 478046 367150 478102
rect 367218 478046 367274 478102
rect 367342 478046 367398 478102
rect 366970 477922 367026 477978
rect 367094 477922 367150 477978
rect 367218 477922 367274 477978
rect 367342 477922 367398 477978
rect 366970 460294 367026 460350
rect 367094 460294 367150 460350
rect 367218 460294 367274 460350
rect 367342 460294 367398 460350
rect 366970 460170 367026 460226
rect 367094 460170 367150 460226
rect 367218 460170 367274 460226
rect 367342 460170 367398 460226
rect 366970 460046 367026 460102
rect 367094 460046 367150 460102
rect 367218 460046 367274 460102
rect 367342 460046 367398 460102
rect 366970 459922 367026 459978
rect 367094 459922 367150 459978
rect 367218 459922 367274 459978
rect 367342 459922 367398 459978
rect 381250 597156 381306 597212
rect 381374 597156 381430 597212
rect 381498 597156 381554 597212
rect 381622 597156 381678 597212
rect 381250 597032 381306 597088
rect 381374 597032 381430 597088
rect 381498 597032 381554 597088
rect 381622 597032 381678 597088
rect 381250 596908 381306 596964
rect 381374 596908 381430 596964
rect 381498 596908 381554 596964
rect 381622 596908 381678 596964
rect 381250 596784 381306 596840
rect 381374 596784 381430 596840
rect 381498 596784 381554 596840
rect 381622 596784 381678 596840
rect 381250 580294 381306 580350
rect 381374 580294 381430 580350
rect 381498 580294 381554 580350
rect 381622 580294 381678 580350
rect 381250 580170 381306 580226
rect 381374 580170 381430 580226
rect 381498 580170 381554 580226
rect 381622 580170 381678 580226
rect 381250 580046 381306 580102
rect 381374 580046 381430 580102
rect 381498 580046 381554 580102
rect 381622 580046 381678 580102
rect 381250 579922 381306 579978
rect 381374 579922 381430 579978
rect 381498 579922 381554 579978
rect 381622 579922 381678 579978
rect 381250 562294 381306 562350
rect 381374 562294 381430 562350
rect 381498 562294 381554 562350
rect 381622 562294 381678 562350
rect 381250 562170 381306 562226
rect 381374 562170 381430 562226
rect 381498 562170 381554 562226
rect 381622 562170 381678 562226
rect 381250 562046 381306 562102
rect 381374 562046 381430 562102
rect 381498 562046 381554 562102
rect 381622 562046 381678 562102
rect 381250 561922 381306 561978
rect 381374 561922 381430 561978
rect 381498 561922 381554 561978
rect 381622 561922 381678 561978
rect 381250 544294 381306 544350
rect 381374 544294 381430 544350
rect 381498 544294 381554 544350
rect 381622 544294 381678 544350
rect 381250 544170 381306 544226
rect 381374 544170 381430 544226
rect 381498 544170 381554 544226
rect 381622 544170 381678 544226
rect 381250 544046 381306 544102
rect 381374 544046 381430 544102
rect 381498 544046 381554 544102
rect 381622 544046 381678 544102
rect 381250 543922 381306 543978
rect 381374 543922 381430 543978
rect 381498 543922 381554 543978
rect 381622 543922 381678 543978
rect 381250 526294 381306 526350
rect 381374 526294 381430 526350
rect 381498 526294 381554 526350
rect 381622 526294 381678 526350
rect 381250 526170 381306 526226
rect 381374 526170 381430 526226
rect 381498 526170 381554 526226
rect 381622 526170 381678 526226
rect 381250 526046 381306 526102
rect 381374 526046 381430 526102
rect 381498 526046 381554 526102
rect 381622 526046 381678 526102
rect 381250 525922 381306 525978
rect 381374 525922 381430 525978
rect 381498 525922 381554 525978
rect 381622 525922 381678 525978
rect 381250 508294 381306 508350
rect 381374 508294 381430 508350
rect 381498 508294 381554 508350
rect 381622 508294 381678 508350
rect 381250 508170 381306 508226
rect 381374 508170 381430 508226
rect 381498 508170 381554 508226
rect 381622 508170 381678 508226
rect 381250 508046 381306 508102
rect 381374 508046 381430 508102
rect 381498 508046 381554 508102
rect 381622 508046 381678 508102
rect 381250 507922 381306 507978
rect 381374 507922 381430 507978
rect 381498 507922 381554 507978
rect 381622 507922 381678 507978
rect 381250 490294 381306 490350
rect 381374 490294 381430 490350
rect 381498 490294 381554 490350
rect 381622 490294 381678 490350
rect 381250 490170 381306 490226
rect 381374 490170 381430 490226
rect 381498 490170 381554 490226
rect 381622 490170 381678 490226
rect 381250 490046 381306 490102
rect 381374 490046 381430 490102
rect 381498 490046 381554 490102
rect 381622 490046 381678 490102
rect 381250 489922 381306 489978
rect 381374 489922 381430 489978
rect 381498 489922 381554 489978
rect 381622 489922 381678 489978
rect 381250 472294 381306 472350
rect 381374 472294 381430 472350
rect 381498 472294 381554 472350
rect 381622 472294 381678 472350
rect 381250 472170 381306 472226
rect 381374 472170 381430 472226
rect 381498 472170 381554 472226
rect 381622 472170 381678 472226
rect 381250 472046 381306 472102
rect 381374 472046 381430 472102
rect 381498 472046 381554 472102
rect 381622 472046 381678 472102
rect 381250 471922 381306 471978
rect 381374 471922 381430 471978
rect 381498 471922 381554 471978
rect 381622 471922 381678 471978
rect 204970 442294 205026 442350
rect 205094 442294 205150 442350
rect 205218 442294 205274 442350
rect 205342 442294 205398 442350
rect 204970 442170 205026 442226
rect 205094 442170 205150 442226
rect 205218 442170 205274 442226
rect 205342 442170 205398 442226
rect 204970 442046 205026 442102
rect 205094 442046 205150 442102
rect 205218 442046 205274 442102
rect 205342 442046 205398 442102
rect 204970 441922 205026 441978
rect 205094 441922 205150 441978
rect 205218 441922 205274 441978
rect 205342 441922 205398 441978
rect 204970 424294 205026 424350
rect 205094 424294 205150 424350
rect 205218 424294 205274 424350
rect 205342 424294 205398 424350
rect 204970 424170 205026 424226
rect 205094 424170 205150 424226
rect 205218 424170 205274 424226
rect 205342 424170 205398 424226
rect 204970 424046 205026 424102
rect 205094 424046 205150 424102
rect 205218 424046 205274 424102
rect 205342 424046 205398 424102
rect 204970 423922 205026 423978
rect 205094 423922 205150 423978
rect 205218 423922 205274 423978
rect 205342 423922 205398 423978
rect 204970 406294 205026 406350
rect 205094 406294 205150 406350
rect 205218 406294 205274 406350
rect 205342 406294 205398 406350
rect 204970 406170 205026 406226
rect 205094 406170 205150 406226
rect 205218 406170 205274 406226
rect 205342 406170 205398 406226
rect 204970 406046 205026 406102
rect 205094 406046 205150 406102
rect 205218 406046 205274 406102
rect 205342 406046 205398 406102
rect 204970 405922 205026 405978
rect 205094 405922 205150 405978
rect 205218 405922 205274 405978
rect 205342 405922 205398 405978
rect 204970 388294 205026 388350
rect 205094 388294 205150 388350
rect 205218 388294 205274 388350
rect 205342 388294 205398 388350
rect 204970 388170 205026 388226
rect 205094 388170 205150 388226
rect 205218 388170 205274 388226
rect 205342 388170 205398 388226
rect 204970 388046 205026 388102
rect 205094 388046 205150 388102
rect 205218 388046 205274 388102
rect 205342 388046 205398 388102
rect 204970 387922 205026 387978
rect 205094 387922 205150 387978
rect 205218 387922 205274 387978
rect 205342 387922 205398 387978
rect 204970 370294 205026 370350
rect 205094 370294 205150 370350
rect 205218 370294 205274 370350
rect 205342 370294 205398 370350
rect 204970 370170 205026 370226
rect 205094 370170 205150 370226
rect 205218 370170 205274 370226
rect 205342 370170 205398 370226
rect 204970 370046 205026 370102
rect 205094 370046 205150 370102
rect 205218 370046 205274 370102
rect 205342 370046 205398 370102
rect 204970 369922 205026 369978
rect 205094 369922 205150 369978
rect 205218 369922 205274 369978
rect 205342 369922 205398 369978
rect 204970 352294 205026 352350
rect 205094 352294 205150 352350
rect 205218 352294 205274 352350
rect 205342 352294 205398 352350
rect 204970 352170 205026 352226
rect 205094 352170 205150 352226
rect 205218 352170 205274 352226
rect 205342 352170 205398 352226
rect 204970 352046 205026 352102
rect 205094 352046 205150 352102
rect 205218 352046 205274 352102
rect 205342 352046 205398 352102
rect 204970 351922 205026 351978
rect 205094 351922 205150 351978
rect 205218 351922 205274 351978
rect 205342 351922 205398 351978
rect 204970 334294 205026 334350
rect 205094 334294 205150 334350
rect 205218 334294 205274 334350
rect 205342 334294 205398 334350
rect 204970 334170 205026 334226
rect 205094 334170 205150 334226
rect 205218 334170 205274 334226
rect 205342 334170 205398 334226
rect 204970 334046 205026 334102
rect 205094 334046 205150 334102
rect 205218 334046 205274 334102
rect 205342 334046 205398 334102
rect 204970 333922 205026 333978
rect 205094 333922 205150 333978
rect 205218 333922 205274 333978
rect 205342 333922 205398 333978
rect 381250 454294 381306 454350
rect 381374 454294 381430 454350
rect 381498 454294 381554 454350
rect 381622 454294 381678 454350
rect 381250 454170 381306 454226
rect 381374 454170 381430 454226
rect 381498 454170 381554 454226
rect 381622 454170 381678 454226
rect 381250 454046 381306 454102
rect 381374 454046 381430 454102
rect 381498 454046 381554 454102
rect 381622 454046 381678 454102
rect 381250 453922 381306 453978
rect 381374 453922 381430 453978
rect 381498 453922 381554 453978
rect 381622 453922 381678 453978
rect 381250 436294 381306 436350
rect 381374 436294 381430 436350
rect 381498 436294 381554 436350
rect 381622 436294 381678 436350
rect 381250 436170 381306 436226
rect 381374 436170 381430 436226
rect 381498 436170 381554 436226
rect 381622 436170 381678 436226
rect 381250 436046 381306 436102
rect 381374 436046 381430 436102
rect 381498 436046 381554 436102
rect 381622 436046 381678 436102
rect 381250 435922 381306 435978
rect 381374 435922 381430 435978
rect 381498 435922 381554 435978
rect 381622 435922 381678 435978
rect 381250 418294 381306 418350
rect 381374 418294 381430 418350
rect 381498 418294 381554 418350
rect 381622 418294 381678 418350
rect 381250 418170 381306 418226
rect 381374 418170 381430 418226
rect 381498 418170 381554 418226
rect 381622 418170 381678 418226
rect 381250 418046 381306 418102
rect 381374 418046 381430 418102
rect 381498 418046 381554 418102
rect 381622 418046 381678 418102
rect 381250 417922 381306 417978
rect 381374 417922 381430 417978
rect 381498 417922 381554 417978
rect 381622 417922 381678 417978
rect 381250 400294 381306 400350
rect 381374 400294 381430 400350
rect 381498 400294 381554 400350
rect 381622 400294 381678 400350
rect 381250 400170 381306 400226
rect 381374 400170 381430 400226
rect 381498 400170 381554 400226
rect 381622 400170 381678 400226
rect 381250 400046 381306 400102
rect 381374 400046 381430 400102
rect 381498 400046 381554 400102
rect 381622 400046 381678 400102
rect 381250 399922 381306 399978
rect 381374 399922 381430 399978
rect 381498 399922 381554 399978
rect 381622 399922 381678 399978
rect 381250 382294 381306 382350
rect 381374 382294 381430 382350
rect 381498 382294 381554 382350
rect 381622 382294 381678 382350
rect 381250 382170 381306 382226
rect 381374 382170 381430 382226
rect 381498 382170 381554 382226
rect 381622 382170 381678 382226
rect 381250 382046 381306 382102
rect 381374 382046 381430 382102
rect 381498 382046 381554 382102
rect 381622 382046 381678 382102
rect 381250 381922 381306 381978
rect 381374 381922 381430 381978
rect 381498 381922 381554 381978
rect 381622 381922 381678 381978
rect 381250 364294 381306 364350
rect 381374 364294 381430 364350
rect 381498 364294 381554 364350
rect 381622 364294 381678 364350
rect 381250 364170 381306 364226
rect 381374 364170 381430 364226
rect 381498 364170 381554 364226
rect 381622 364170 381678 364226
rect 381250 364046 381306 364102
rect 381374 364046 381430 364102
rect 381498 364046 381554 364102
rect 381622 364046 381678 364102
rect 381250 363922 381306 363978
rect 381374 363922 381430 363978
rect 381498 363922 381554 363978
rect 381622 363922 381678 363978
rect 381250 346294 381306 346350
rect 381374 346294 381430 346350
rect 381498 346294 381554 346350
rect 381622 346294 381678 346350
rect 381250 346170 381306 346226
rect 381374 346170 381430 346226
rect 381498 346170 381554 346226
rect 381622 346170 381678 346226
rect 381250 346046 381306 346102
rect 381374 346046 381430 346102
rect 381498 346046 381554 346102
rect 381622 346046 381678 346102
rect 381250 345922 381306 345978
rect 381374 345922 381430 345978
rect 381498 345922 381554 345978
rect 381622 345922 381678 345978
rect 381250 328294 381306 328350
rect 381374 328294 381430 328350
rect 381498 328294 381554 328350
rect 381622 328294 381678 328350
rect 381250 328170 381306 328226
rect 381374 328170 381430 328226
rect 381498 328170 381554 328226
rect 381622 328170 381678 328226
rect 381250 328046 381306 328102
rect 381374 328046 381430 328102
rect 381498 328046 381554 328102
rect 381622 328046 381678 328102
rect 381250 327922 381306 327978
rect 381374 327922 381430 327978
rect 381498 327922 381554 327978
rect 381622 327922 381678 327978
rect 204970 316294 205026 316350
rect 205094 316294 205150 316350
rect 205218 316294 205274 316350
rect 205342 316294 205398 316350
rect 204970 316170 205026 316226
rect 205094 316170 205150 316226
rect 205218 316170 205274 316226
rect 205342 316170 205398 316226
rect 204970 316046 205026 316102
rect 205094 316046 205150 316102
rect 205218 316046 205274 316102
rect 205342 316046 205398 316102
rect 204970 315922 205026 315978
rect 205094 315922 205150 315978
rect 205218 315922 205274 315978
rect 205342 315922 205398 315978
rect 204970 298294 205026 298350
rect 205094 298294 205150 298350
rect 205218 298294 205274 298350
rect 205342 298294 205398 298350
rect 222970 316294 223026 316350
rect 223094 316294 223150 316350
rect 223218 316294 223274 316350
rect 223342 316294 223398 316350
rect 222970 316170 223026 316226
rect 223094 316170 223150 316226
rect 223218 316170 223274 316226
rect 223342 316170 223398 316226
rect 222970 316046 223026 316102
rect 223094 316046 223150 316102
rect 223218 316046 223274 316102
rect 223342 316046 223398 316102
rect 222970 315922 223026 315978
rect 223094 315922 223150 315978
rect 223218 315922 223274 315978
rect 223342 315922 223398 315978
rect 222970 298366 223026 298422
rect 223094 298366 223150 298422
rect 223218 298366 223274 298422
rect 223342 298366 223398 298422
rect 240970 316294 241026 316350
rect 241094 316294 241150 316350
rect 241218 316294 241274 316350
rect 241342 316294 241398 316350
rect 240970 316170 241026 316226
rect 241094 316170 241150 316226
rect 241218 316170 241274 316226
rect 241342 316170 241398 316226
rect 240970 316046 241026 316102
rect 241094 316046 241150 316102
rect 241218 316046 241274 316102
rect 241342 316046 241398 316102
rect 240970 315922 241026 315978
rect 241094 315922 241150 315978
rect 241218 315922 241274 315978
rect 241342 315922 241398 315978
rect 240970 298366 241026 298422
rect 241094 298366 241150 298422
rect 241218 298366 241274 298422
rect 241342 298366 241398 298422
rect 258970 316294 259026 316350
rect 259094 316294 259150 316350
rect 259218 316294 259274 316350
rect 259342 316294 259398 316350
rect 258970 316170 259026 316226
rect 259094 316170 259150 316226
rect 259218 316170 259274 316226
rect 259342 316170 259398 316226
rect 258970 316046 259026 316102
rect 259094 316046 259150 316102
rect 259218 316046 259274 316102
rect 259342 316046 259398 316102
rect 258970 315922 259026 315978
rect 259094 315922 259150 315978
rect 259218 315922 259274 315978
rect 259342 315922 259398 315978
rect 258970 298366 259026 298422
rect 259094 298366 259150 298422
rect 259218 298366 259274 298422
rect 259342 298366 259398 298422
rect 276970 316294 277026 316350
rect 277094 316294 277150 316350
rect 277218 316294 277274 316350
rect 277342 316294 277398 316350
rect 276970 316170 277026 316226
rect 277094 316170 277150 316226
rect 277218 316170 277274 316226
rect 277342 316170 277398 316226
rect 276970 316046 277026 316102
rect 277094 316046 277150 316102
rect 277218 316046 277274 316102
rect 277342 316046 277398 316102
rect 276970 315922 277026 315978
rect 277094 315922 277150 315978
rect 277218 315922 277274 315978
rect 277342 315922 277398 315978
rect 276970 298366 277026 298422
rect 277094 298366 277150 298422
rect 277218 298366 277274 298422
rect 277342 298366 277398 298422
rect 294970 316294 295026 316350
rect 295094 316294 295150 316350
rect 295218 316294 295274 316350
rect 295342 316294 295398 316350
rect 294970 316170 295026 316226
rect 295094 316170 295150 316226
rect 295218 316170 295274 316226
rect 295342 316170 295398 316226
rect 294970 316046 295026 316102
rect 295094 316046 295150 316102
rect 295218 316046 295274 316102
rect 295342 316046 295398 316102
rect 294970 315922 295026 315978
rect 295094 315922 295150 315978
rect 295218 315922 295274 315978
rect 295342 315922 295398 315978
rect 294970 298366 295026 298422
rect 295094 298366 295150 298422
rect 295218 298366 295274 298422
rect 295342 298366 295398 298422
rect 312970 316294 313026 316350
rect 313094 316294 313150 316350
rect 313218 316294 313274 316350
rect 313342 316294 313398 316350
rect 312970 316170 313026 316226
rect 313094 316170 313150 316226
rect 313218 316170 313274 316226
rect 313342 316170 313398 316226
rect 312970 316046 313026 316102
rect 313094 316046 313150 316102
rect 313218 316046 313274 316102
rect 313342 316046 313398 316102
rect 312970 315922 313026 315978
rect 313094 315922 313150 315978
rect 313218 315922 313274 315978
rect 313342 315922 313398 315978
rect 312970 298366 313026 298422
rect 313094 298366 313150 298422
rect 313218 298366 313274 298422
rect 313342 298366 313398 298422
rect 330970 316294 331026 316350
rect 331094 316294 331150 316350
rect 331218 316294 331274 316350
rect 331342 316294 331398 316350
rect 330970 316170 331026 316226
rect 331094 316170 331150 316226
rect 331218 316170 331274 316226
rect 331342 316170 331398 316226
rect 330970 316046 331026 316102
rect 331094 316046 331150 316102
rect 331218 316046 331274 316102
rect 331342 316046 331398 316102
rect 330970 315922 331026 315978
rect 331094 315922 331150 315978
rect 331218 315922 331274 315978
rect 331342 315922 331398 315978
rect 330970 298366 331026 298422
rect 331094 298366 331150 298422
rect 331218 298366 331274 298422
rect 331342 298366 331398 298422
rect 348970 316294 349026 316350
rect 349094 316294 349150 316350
rect 349218 316294 349274 316350
rect 349342 316294 349398 316350
rect 348970 316170 349026 316226
rect 349094 316170 349150 316226
rect 349218 316170 349274 316226
rect 349342 316170 349398 316226
rect 348970 316046 349026 316102
rect 349094 316046 349150 316102
rect 349218 316046 349274 316102
rect 349342 316046 349398 316102
rect 348970 315922 349026 315978
rect 349094 315922 349150 315978
rect 349218 315922 349274 315978
rect 349342 315922 349398 315978
rect 348970 298366 349026 298422
rect 349094 298366 349150 298422
rect 349218 298366 349274 298422
rect 349342 298366 349398 298422
rect 366970 316294 367026 316350
rect 367094 316294 367150 316350
rect 367218 316294 367274 316350
rect 367342 316294 367398 316350
rect 366970 316170 367026 316226
rect 367094 316170 367150 316226
rect 367218 316170 367274 316226
rect 367342 316170 367398 316226
rect 366970 316046 367026 316102
rect 367094 316046 367150 316102
rect 367218 316046 367274 316102
rect 367342 316046 367398 316102
rect 366970 315922 367026 315978
rect 367094 315922 367150 315978
rect 367218 315922 367274 315978
rect 367342 315922 367398 315978
rect 381250 310294 381306 310350
rect 381374 310294 381430 310350
rect 381498 310294 381554 310350
rect 381622 310294 381678 310350
rect 381250 310170 381306 310226
rect 381374 310170 381430 310226
rect 381498 310170 381554 310226
rect 381622 310170 381678 310226
rect 381250 310046 381306 310102
rect 381374 310046 381430 310102
rect 381498 310046 381554 310102
rect 381622 310046 381678 310102
rect 366970 298366 367026 298422
rect 367094 298366 367150 298422
rect 367218 298366 367274 298422
rect 367342 298366 367398 298422
rect 204970 298170 205026 298226
rect 205094 298170 205150 298226
rect 205218 298170 205274 298226
rect 205342 298170 205398 298226
rect 204970 298046 205026 298102
rect 205094 298046 205150 298102
rect 205218 298046 205274 298102
rect 205342 298046 205398 298102
rect 204970 297922 205026 297978
rect 205094 297922 205150 297978
rect 205218 297922 205274 297978
rect 205342 297922 205398 297978
rect 204970 280294 205026 280350
rect 205094 280294 205150 280350
rect 205218 280294 205274 280350
rect 205342 280294 205398 280350
rect 204970 280170 205026 280226
rect 205094 280170 205150 280226
rect 205218 280170 205274 280226
rect 205342 280170 205398 280226
rect 204970 280046 205026 280102
rect 205094 280046 205150 280102
rect 205218 280046 205274 280102
rect 205342 280046 205398 280102
rect 204970 279922 205026 279978
rect 205094 279922 205150 279978
rect 205218 279922 205274 279978
rect 205342 279922 205398 279978
rect 204970 262294 205026 262350
rect 205094 262294 205150 262350
rect 205218 262294 205274 262350
rect 205342 262294 205398 262350
rect 204970 262170 205026 262226
rect 205094 262170 205150 262226
rect 205218 262170 205274 262226
rect 205342 262170 205398 262226
rect 204970 262046 205026 262102
rect 205094 262046 205150 262102
rect 205218 262046 205274 262102
rect 205342 262046 205398 262102
rect 204970 261922 205026 261978
rect 205094 261922 205150 261978
rect 205218 261922 205274 261978
rect 205342 261922 205398 261978
rect 204970 244294 205026 244350
rect 205094 244294 205150 244350
rect 205218 244294 205274 244350
rect 205342 244294 205398 244350
rect 204970 244170 205026 244226
rect 205094 244170 205150 244226
rect 205218 244170 205274 244226
rect 205342 244170 205398 244226
rect 204970 244046 205026 244102
rect 205094 244046 205150 244102
rect 205218 244046 205274 244102
rect 205342 244046 205398 244102
rect 204970 243922 205026 243978
rect 205094 243922 205150 243978
rect 205218 243922 205274 243978
rect 205342 243922 205398 243978
rect 204970 226294 205026 226350
rect 205094 226294 205150 226350
rect 205218 226294 205274 226350
rect 205342 226294 205398 226350
rect 204970 226170 205026 226226
rect 205094 226170 205150 226226
rect 205218 226170 205274 226226
rect 205342 226170 205398 226226
rect 204970 226046 205026 226102
rect 205094 226046 205150 226102
rect 205218 226046 205274 226102
rect 205342 226046 205398 226102
rect 204970 225922 205026 225978
rect 205094 225922 205150 225978
rect 205218 225922 205274 225978
rect 205342 225922 205398 225978
rect 204970 208294 205026 208350
rect 205094 208294 205150 208350
rect 205218 208294 205274 208350
rect 205342 208294 205398 208350
rect 204970 208170 205026 208226
rect 205094 208170 205150 208226
rect 205218 208170 205274 208226
rect 205342 208170 205398 208226
rect 204970 208046 205026 208102
rect 205094 208046 205150 208102
rect 205218 208046 205274 208102
rect 205342 208046 205398 208102
rect 204970 207922 205026 207978
rect 205094 207922 205150 207978
rect 205218 207922 205274 207978
rect 205342 207922 205398 207978
rect 204970 190294 205026 190350
rect 205094 190294 205150 190350
rect 205218 190294 205274 190350
rect 205342 190294 205398 190350
rect 204970 190170 205026 190226
rect 205094 190170 205150 190226
rect 205218 190170 205274 190226
rect 205342 190170 205398 190226
rect 204970 190046 205026 190102
rect 205094 190046 205150 190102
rect 205218 190046 205274 190102
rect 205342 190046 205398 190102
rect 204970 189922 205026 189978
rect 205094 189922 205150 189978
rect 205218 189922 205274 189978
rect 205342 189922 205398 189978
rect 204970 172294 205026 172350
rect 205094 172294 205150 172350
rect 205218 172294 205274 172350
rect 205342 172294 205398 172350
rect 204970 172170 205026 172226
rect 205094 172170 205150 172226
rect 205218 172170 205274 172226
rect 205342 172170 205398 172226
rect 204970 172046 205026 172102
rect 205094 172046 205150 172102
rect 205218 172046 205274 172102
rect 205342 172046 205398 172102
rect 204970 171922 205026 171978
rect 205094 171922 205150 171978
rect 205218 171922 205274 171978
rect 205342 171922 205398 171978
rect 204970 154294 205026 154350
rect 205094 154294 205150 154350
rect 205218 154294 205274 154350
rect 205342 154294 205398 154350
rect 204970 154170 205026 154226
rect 205094 154170 205150 154226
rect 205218 154170 205274 154226
rect 205342 154170 205398 154226
rect 204970 154046 205026 154102
rect 205094 154046 205150 154102
rect 205218 154046 205274 154102
rect 205342 154046 205398 154102
rect 204970 153922 205026 153978
rect 205094 153922 205150 153978
rect 205218 153922 205274 153978
rect 205342 153922 205398 153978
rect 219250 148366 219306 148422
rect 219374 148366 219430 148422
rect 219498 148366 219554 148422
rect 219622 148366 219678 148422
rect 222970 154294 223026 154350
rect 223094 154294 223150 154350
rect 223218 154294 223274 154350
rect 223342 154294 223398 154350
rect 222970 154170 223026 154226
rect 223094 154170 223150 154226
rect 223218 154170 223274 154226
rect 223342 154170 223398 154226
rect 222970 154046 223026 154102
rect 223094 154046 223150 154102
rect 223218 154046 223274 154102
rect 223342 154046 223398 154102
rect 222970 153922 223026 153978
rect 223094 153922 223150 153978
rect 223218 153922 223274 153978
rect 223342 153922 223398 153978
rect 237250 148366 237306 148422
rect 237374 148366 237430 148422
rect 237498 148366 237554 148422
rect 237622 148366 237678 148422
rect 240970 154294 241026 154350
rect 241094 154294 241150 154350
rect 241218 154294 241274 154350
rect 241342 154294 241398 154350
rect 240970 154170 241026 154226
rect 241094 154170 241150 154226
rect 241218 154170 241274 154226
rect 241342 154170 241398 154226
rect 240970 154046 241026 154102
rect 241094 154046 241150 154102
rect 241218 154046 241274 154102
rect 241342 154046 241398 154102
rect 240970 153922 241026 153978
rect 241094 153922 241150 153978
rect 241218 153922 241274 153978
rect 241342 153922 241398 153978
rect 255250 148366 255306 148422
rect 255374 148366 255430 148422
rect 255498 148366 255554 148422
rect 255622 148366 255678 148422
rect 258970 154294 259026 154350
rect 259094 154294 259150 154350
rect 259218 154294 259274 154350
rect 259342 154294 259398 154350
rect 258970 154170 259026 154226
rect 259094 154170 259150 154226
rect 259218 154170 259274 154226
rect 259342 154170 259398 154226
rect 258970 154046 259026 154102
rect 259094 154046 259150 154102
rect 259218 154046 259274 154102
rect 259342 154046 259398 154102
rect 258970 153922 259026 153978
rect 259094 153922 259150 153978
rect 259218 153922 259274 153978
rect 259342 153922 259398 153978
rect 273250 148366 273306 148422
rect 273374 148366 273430 148422
rect 273498 148366 273554 148422
rect 273622 148366 273678 148422
rect 276970 154294 277026 154350
rect 277094 154294 277150 154350
rect 277218 154294 277274 154350
rect 277342 154294 277398 154350
rect 276970 154170 277026 154226
rect 277094 154170 277150 154226
rect 277218 154170 277274 154226
rect 277342 154170 277398 154226
rect 276970 154046 277026 154102
rect 277094 154046 277150 154102
rect 277218 154046 277274 154102
rect 277342 154046 277398 154102
rect 276970 153922 277026 153978
rect 277094 153922 277150 153978
rect 277218 153922 277274 153978
rect 277342 153922 277398 153978
rect 291250 148366 291306 148422
rect 291374 148366 291430 148422
rect 291498 148366 291554 148422
rect 291622 148366 291678 148422
rect 294970 154294 295026 154350
rect 295094 154294 295150 154350
rect 295218 154294 295274 154350
rect 295342 154294 295398 154350
rect 294970 154170 295026 154226
rect 295094 154170 295150 154226
rect 295218 154170 295274 154226
rect 295342 154170 295398 154226
rect 294970 154046 295026 154102
rect 295094 154046 295150 154102
rect 295218 154046 295274 154102
rect 295342 154046 295398 154102
rect 294970 153922 295026 153978
rect 295094 153922 295150 153978
rect 295218 153922 295274 153978
rect 295342 153922 295398 153978
rect 309250 148366 309306 148422
rect 309374 148366 309430 148422
rect 309498 148366 309554 148422
rect 309622 148366 309678 148422
rect 312970 154294 313026 154350
rect 313094 154294 313150 154350
rect 313218 154294 313274 154350
rect 313342 154294 313398 154350
rect 312970 154170 313026 154226
rect 313094 154170 313150 154226
rect 313218 154170 313274 154226
rect 313342 154170 313398 154226
rect 312970 154046 313026 154102
rect 313094 154046 313150 154102
rect 313218 154046 313274 154102
rect 313342 154046 313398 154102
rect 312970 153922 313026 153978
rect 313094 153922 313150 153978
rect 313218 153922 313274 153978
rect 313342 153922 313398 153978
rect 327250 148366 327306 148422
rect 327374 148366 327430 148422
rect 327498 148366 327554 148422
rect 327622 148366 327678 148422
rect 330970 154294 331026 154350
rect 331094 154294 331150 154350
rect 331218 154294 331274 154350
rect 331342 154294 331398 154350
rect 330970 154170 331026 154226
rect 331094 154170 331150 154226
rect 331218 154170 331274 154226
rect 331342 154170 331398 154226
rect 330970 154046 331026 154102
rect 331094 154046 331150 154102
rect 331218 154046 331274 154102
rect 331342 154046 331398 154102
rect 330970 153922 331026 153978
rect 331094 153922 331150 153978
rect 331218 153922 331274 153978
rect 331342 153922 331398 153978
rect 345250 148366 345306 148422
rect 345374 148366 345430 148422
rect 345498 148366 345554 148422
rect 345622 148366 345678 148422
rect 348970 154294 349026 154350
rect 349094 154294 349150 154350
rect 349218 154294 349274 154350
rect 349342 154294 349398 154350
rect 348970 154170 349026 154226
rect 349094 154170 349150 154226
rect 349218 154170 349274 154226
rect 349342 154170 349398 154226
rect 348970 154046 349026 154102
rect 349094 154046 349150 154102
rect 349218 154046 349274 154102
rect 349342 154046 349398 154102
rect 348970 153922 349026 153978
rect 349094 153922 349150 153978
rect 349218 153922 349274 153978
rect 349342 153922 349398 153978
rect 363250 148366 363306 148422
rect 363374 148366 363430 148422
rect 363498 148366 363554 148422
rect 363622 148366 363678 148422
rect 366970 154294 367026 154350
rect 367094 154294 367150 154350
rect 367218 154294 367274 154350
rect 367342 154294 367398 154350
rect 366970 154170 367026 154226
rect 367094 154170 367150 154226
rect 367218 154170 367274 154226
rect 367342 154170 367398 154226
rect 366970 154046 367026 154102
rect 367094 154046 367150 154102
rect 367218 154046 367274 154102
rect 367342 154046 367398 154102
rect 366970 153922 367026 153978
rect 367094 153922 367150 153978
rect 367218 153922 367274 153978
rect 367342 153922 367398 153978
rect 381250 309922 381306 309978
rect 381374 309922 381430 309978
rect 381498 309922 381554 309978
rect 381622 309922 381678 309978
rect 381250 292294 381306 292350
rect 381374 292294 381430 292350
rect 381498 292294 381554 292350
rect 381622 292294 381678 292350
rect 381250 292170 381306 292226
rect 381374 292170 381430 292226
rect 381498 292170 381554 292226
rect 381622 292170 381678 292226
rect 381250 292046 381306 292102
rect 381374 292046 381430 292102
rect 381498 292046 381554 292102
rect 381622 292046 381678 292102
rect 381250 291922 381306 291978
rect 381374 291922 381430 291978
rect 381498 291922 381554 291978
rect 381622 291922 381678 291978
rect 381250 274294 381306 274350
rect 381374 274294 381430 274350
rect 381498 274294 381554 274350
rect 381622 274294 381678 274350
rect 381250 274170 381306 274226
rect 381374 274170 381430 274226
rect 381498 274170 381554 274226
rect 381622 274170 381678 274226
rect 381250 274046 381306 274102
rect 381374 274046 381430 274102
rect 381498 274046 381554 274102
rect 381622 274046 381678 274102
rect 381250 273922 381306 273978
rect 381374 273922 381430 273978
rect 381498 273922 381554 273978
rect 381622 273922 381678 273978
rect 381250 256294 381306 256350
rect 381374 256294 381430 256350
rect 381498 256294 381554 256350
rect 381622 256294 381678 256350
rect 381250 256170 381306 256226
rect 381374 256170 381430 256226
rect 381498 256170 381554 256226
rect 381622 256170 381678 256226
rect 381250 256046 381306 256102
rect 381374 256046 381430 256102
rect 381498 256046 381554 256102
rect 381622 256046 381678 256102
rect 381250 255922 381306 255978
rect 381374 255922 381430 255978
rect 381498 255922 381554 255978
rect 381622 255922 381678 255978
rect 381250 238294 381306 238350
rect 381374 238294 381430 238350
rect 381498 238294 381554 238350
rect 381622 238294 381678 238350
rect 381250 238170 381306 238226
rect 381374 238170 381430 238226
rect 381498 238170 381554 238226
rect 381622 238170 381678 238226
rect 381250 238046 381306 238102
rect 381374 238046 381430 238102
rect 381498 238046 381554 238102
rect 381622 238046 381678 238102
rect 381250 237922 381306 237978
rect 381374 237922 381430 237978
rect 381498 237922 381554 237978
rect 381622 237922 381678 237978
rect 381250 220294 381306 220350
rect 381374 220294 381430 220350
rect 381498 220294 381554 220350
rect 381622 220294 381678 220350
rect 381250 220170 381306 220226
rect 381374 220170 381430 220226
rect 381498 220170 381554 220226
rect 381622 220170 381678 220226
rect 381250 220046 381306 220102
rect 381374 220046 381430 220102
rect 381498 220046 381554 220102
rect 381622 220046 381678 220102
rect 381250 219922 381306 219978
rect 381374 219922 381430 219978
rect 381498 219922 381554 219978
rect 381622 219922 381678 219978
rect 381250 202294 381306 202350
rect 381374 202294 381430 202350
rect 381498 202294 381554 202350
rect 381622 202294 381678 202350
rect 381250 202170 381306 202226
rect 381374 202170 381430 202226
rect 381498 202170 381554 202226
rect 381622 202170 381678 202226
rect 381250 202046 381306 202102
rect 381374 202046 381430 202102
rect 381498 202046 381554 202102
rect 381622 202046 381678 202102
rect 381250 201922 381306 201978
rect 381374 201922 381430 201978
rect 381498 201922 381554 201978
rect 381622 201922 381678 201978
rect 381250 184294 381306 184350
rect 381374 184294 381430 184350
rect 381498 184294 381554 184350
rect 381622 184294 381678 184350
rect 381250 184170 381306 184226
rect 381374 184170 381430 184226
rect 381498 184170 381554 184226
rect 381622 184170 381678 184226
rect 381250 184046 381306 184102
rect 381374 184046 381430 184102
rect 381498 184046 381554 184102
rect 381622 184046 381678 184102
rect 381250 183922 381306 183978
rect 381374 183922 381430 183978
rect 381498 183922 381554 183978
rect 381622 183922 381678 183978
rect 381250 166294 381306 166350
rect 381374 166294 381430 166350
rect 381498 166294 381554 166350
rect 381622 166294 381678 166350
rect 381250 166170 381306 166226
rect 381374 166170 381430 166226
rect 381498 166170 381554 166226
rect 381622 166170 381678 166226
rect 381250 166046 381306 166102
rect 381374 166046 381430 166102
rect 381498 166046 381554 166102
rect 381622 166046 381678 166102
rect 381250 165922 381306 165978
rect 381374 165922 381430 165978
rect 381498 165922 381554 165978
rect 381622 165922 381678 165978
rect 204970 136294 205026 136350
rect 205094 136294 205150 136350
rect 205218 136294 205274 136350
rect 205342 136294 205398 136350
rect 204970 136170 205026 136226
rect 205094 136170 205150 136226
rect 205218 136170 205274 136226
rect 205342 136170 205398 136226
rect 204970 136046 205026 136102
rect 205094 136046 205150 136102
rect 205218 136046 205274 136102
rect 205342 136046 205398 136102
rect 204970 135922 205026 135978
rect 205094 135922 205150 135978
rect 205218 135922 205274 135978
rect 205342 135922 205398 135978
rect 204970 118294 205026 118350
rect 205094 118294 205150 118350
rect 205218 118294 205274 118350
rect 205342 118294 205398 118350
rect 204970 118170 205026 118226
rect 205094 118170 205150 118226
rect 205218 118170 205274 118226
rect 205342 118170 205398 118226
rect 204970 118046 205026 118102
rect 205094 118046 205150 118102
rect 205218 118046 205274 118102
rect 205342 118046 205398 118102
rect 204970 117922 205026 117978
rect 205094 117922 205150 117978
rect 205218 117922 205274 117978
rect 205342 117922 205398 117978
rect 204970 100294 205026 100350
rect 205094 100294 205150 100350
rect 205218 100294 205274 100350
rect 205342 100294 205398 100350
rect 204970 100170 205026 100226
rect 205094 100170 205150 100226
rect 205218 100170 205274 100226
rect 205342 100170 205398 100226
rect 204970 100046 205026 100102
rect 205094 100046 205150 100102
rect 205218 100046 205274 100102
rect 205342 100046 205398 100102
rect 204970 99922 205026 99978
rect 205094 99922 205150 99978
rect 205218 99922 205274 99978
rect 205342 99922 205398 99978
rect 204970 82294 205026 82350
rect 205094 82294 205150 82350
rect 205218 82294 205274 82350
rect 205342 82294 205398 82350
rect 204970 82170 205026 82226
rect 205094 82170 205150 82226
rect 205218 82170 205274 82226
rect 205342 82170 205398 82226
rect 204970 82046 205026 82102
rect 205094 82046 205150 82102
rect 205218 82046 205274 82102
rect 205342 82046 205398 82102
rect 204970 81922 205026 81978
rect 205094 81922 205150 81978
rect 205218 81922 205274 81978
rect 205342 81922 205398 81978
rect 204970 64294 205026 64350
rect 205094 64294 205150 64350
rect 205218 64294 205274 64350
rect 205342 64294 205398 64350
rect 204970 64170 205026 64226
rect 205094 64170 205150 64226
rect 205218 64170 205274 64226
rect 205342 64170 205398 64226
rect 204970 64046 205026 64102
rect 205094 64046 205150 64102
rect 205218 64046 205274 64102
rect 205342 64046 205398 64102
rect 204970 63922 205026 63978
rect 205094 63922 205150 63978
rect 205218 63922 205274 63978
rect 205342 63922 205398 63978
rect 204970 46294 205026 46350
rect 205094 46294 205150 46350
rect 205218 46294 205274 46350
rect 205342 46294 205398 46350
rect 204970 46170 205026 46226
rect 205094 46170 205150 46226
rect 205218 46170 205274 46226
rect 205342 46170 205398 46226
rect 204970 46046 205026 46102
rect 205094 46046 205150 46102
rect 205218 46046 205274 46102
rect 205342 46046 205398 46102
rect 204970 45922 205026 45978
rect 205094 45922 205150 45978
rect 205218 45922 205274 45978
rect 205342 45922 205398 45978
rect 204970 28294 205026 28350
rect 205094 28294 205150 28350
rect 205218 28294 205274 28350
rect 205342 28294 205398 28350
rect 204970 28170 205026 28226
rect 205094 28170 205150 28226
rect 205218 28170 205274 28226
rect 205342 28170 205398 28226
rect 204970 28046 205026 28102
rect 205094 28046 205150 28102
rect 205218 28046 205274 28102
rect 205342 28046 205398 28102
rect 204970 27922 205026 27978
rect 205094 27922 205150 27978
rect 205218 27922 205274 27978
rect 205342 27922 205398 27978
rect 204970 10294 205026 10350
rect 205094 10294 205150 10350
rect 205218 10294 205274 10350
rect 205342 10294 205398 10350
rect 204970 10170 205026 10226
rect 205094 10170 205150 10226
rect 205218 10170 205274 10226
rect 205342 10170 205398 10226
rect 204970 10046 205026 10102
rect 205094 10046 205150 10102
rect 205218 10046 205274 10102
rect 205342 10046 205398 10102
rect 204970 9922 205026 9978
rect 205094 9922 205150 9978
rect 205218 9922 205274 9978
rect 205342 9922 205398 9978
rect 204970 -1176 205026 -1120
rect 205094 -1176 205150 -1120
rect 205218 -1176 205274 -1120
rect 205342 -1176 205398 -1120
rect 204970 -1300 205026 -1244
rect 205094 -1300 205150 -1244
rect 205218 -1300 205274 -1244
rect 205342 -1300 205398 -1244
rect 204970 -1424 205026 -1368
rect 205094 -1424 205150 -1368
rect 205218 -1424 205274 -1368
rect 205342 -1424 205398 -1368
rect 204970 -1548 205026 -1492
rect 205094 -1548 205150 -1492
rect 205218 -1548 205274 -1492
rect 205342 -1548 205398 -1492
rect 219250 4294 219306 4350
rect 219374 4294 219430 4350
rect 219498 4294 219554 4350
rect 219622 4294 219678 4350
rect 219250 4170 219306 4226
rect 219374 4170 219430 4226
rect 219498 4170 219554 4226
rect 219622 4170 219678 4226
rect 219250 4046 219306 4102
rect 219374 4046 219430 4102
rect 219498 4046 219554 4102
rect 219622 4046 219678 4102
rect 219250 3922 219306 3978
rect 219374 3922 219430 3978
rect 219498 3922 219554 3978
rect 219622 3922 219678 3978
rect 219250 -216 219306 -160
rect 219374 -216 219430 -160
rect 219498 -216 219554 -160
rect 219622 -216 219678 -160
rect 219250 -340 219306 -284
rect 219374 -340 219430 -284
rect 219498 -340 219554 -284
rect 219622 -340 219678 -284
rect 219250 -464 219306 -408
rect 219374 -464 219430 -408
rect 219498 -464 219554 -408
rect 219622 -464 219678 -408
rect 219250 -588 219306 -532
rect 219374 -588 219430 -532
rect 219498 -588 219554 -532
rect 219622 -588 219678 -532
rect 237250 4294 237306 4350
rect 237374 4294 237430 4350
rect 237498 4294 237554 4350
rect 237622 4294 237678 4350
rect 237250 4170 237306 4226
rect 237374 4170 237430 4226
rect 237498 4170 237554 4226
rect 237622 4170 237678 4226
rect 237250 4046 237306 4102
rect 237374 4046 237430 4102
rect 237498 4046 237554 4102
rect 237622 4046 237678 4102
rect 237250 3922 237306 3978
rect 237374 3922 237430 3978
rect 237498 3922 237554 3978
rect 237622 3922 237678 3978
rect 237250 -216 237306 -160
rect 237374 -216 237430 -160
rect 237498 -216 237554 -160
rect 237622 -216 237678 -160
rect 237250 -340 237306 -284
rect 237374 -340 237430 -284
rect 237498 -340 237554 -284
rect 237622 -340 237678 -284
rect 237250 -464 237306 -408
rect 237374 -464 237430 -408
rect 237498 -464 237554 -408
rect 237622 -464 237678 -408
rect 237250 -588 237306 -532
rect 237374 -588 237430 -532
rect 237498 -588 237554 -532
rect 237622 -588 237678 -532
rect 255250 4294 255306 4350
rect 255374 4294 255430 4350
rect 255498 4294 255554 4350
rect 255622 4294 255678 4350
rect 255250 4170 255306 4226
rect 255374 4170 255430 4226
rect 255498 4170 255554 4226
rect 255622 4170 255678 4226
rect 255250 4046 255306 4102
rect 255374 4046 255430 4102
rect 255498 4046 255554 4102
rect 255622 4046 255678 4102
rect 255250 3922 255306 3978
rect 255374 3922 255430 3978
rect 255498 3922 255554 3978
rect 255622 3922 255678 3978
rect 255250 -216 255306 -160
rect 255374 -216 255430 -160
rect 255498 -216 255554 -160
rect 255622 -216 255678 -160
rect 255250 -340 255306 -284
rect 255374 -340 255430 -284
rect 255498 -340 255554 -284
rect 255622 -340 255678 -284
rect 255250 -464 255306 -408
rect 255374 -464 255430 -408
rect 255498 -464 255554 -408
rect 255622 -464 255678 -408
rect 255250 -588 255306 -532
rect 255374 -588 255430 -532
rect 255498 -588 255554 -532
rect 255622 -588 255678 -532
rect 273250 4294 273306 4350
rect 273374 4294 273430 4350
rect 273498 4294 273554 4350
rect 273622 4294 273678 4350
rect 273250 4170 273306 4226
rect 273374 4170 273430 4226
rect 273498 4170 273554 4226
rect 273622 4170 273678 4226
rect 273250 4046 273306 4102
rect 273374 4046 273430 4102
rect 273498 4046 273554 4102
rect 273622 4046 273678 4102
rect 273250 3922 273306 3978
rect 273374 3922 273430 3978
rect 273498 3922 273554 3978
rect 273622 3922 273678 3978
rect 273250 -216 273306 -160
rect 273374 -216 273430 -160
rect 273498 -216 273554 -160
rect 273622 -216 273678 -160
rect 273250 -340 273306 -284
rect 273374 -340 273430 -284
rect 273498 -340 273554 -284
rect 273622 -340 273678 -284
rect 273250 -464 273306 -408
rect 273374 -464 273430 -408
rect 273498 -464 273554 -408
rect 273622 -464 273678 -408
rect 273250 -588 273306 -532
rect 273374 -588 273430 -532
rect 273498 -588 273554 -532
rect 273622 -588 273678 -532
rect 291250 4294 291306 4350
rect 291374 4294 291430 4350
rect 291498 4294 291554 4350
rect 291622 4294 291678 4350
rect 291250 4170 291306 4226
rect 291374 4170 291430 4226
rect 291498 4170 291554 4226
rect 291622 4170 291678 4226
rect 291250 4046 291306 4102
rect 291374 4046 291430 4102
rect 291498 4046 291554 4102
rect 291622 4046 291678 4102
rect 291250 3922 291306 3978
rect 291374 3922 291430 3978
rect 291498 3922 291554 3978
rect 291622 3922 291678 3978
rect 291250 -216 291306 -160
rect 291374 -216 291430 -160
rect 291498 -216 291554 -160
rect 291622 -216 291678 -160
rect 291250 -340 291306 -284
rect 291374 -340 291430 -284
rect 291498 -340 291554 -284
rect 291622 -340 291678 -284
rect 291250 -464 291306 -408
rect 291374 -464 291430 -408
rect 291498 -464 291554 -408
rect 291622 -464 291678 -408
rect 291250 -588 291306 -532
rect 291374 -588 291430 -532
rect 291498 -588 291554 -532
rect 291622 -588 291678 -532
rect 309250 4294 309306 4350
rect 309374 4294 309430 4350
rect 309498 4294 309554 4350
rect 309622 4294 309678 4350
rect 309250 4170 309306 4226
rect 309374 4170 309430 4226
rect 309498 4170 309554 4226
rect 309622 4170 309678 4226
rect 309250 4046 309306 4102
rect 309374 4046 309430 4102
rect 309498 4046 309554 4102
rect 309622 4046 309678 4102
rect 309250 3922 309306 3978
rect 309374 3922 309430 3978
rect 309498 3922 309554 3978
rect 309622 3922 309678 3978
rect 309250 -216 309306 -160
rect 309374 -216 309430 -160
rect 309498 -216 309554 -160
rect 309622 -216 309678 -160
rect 309250 -340 309306 -284
rect 309374 -340 309430 -284
rect 309498 -340 309554 -284
rect 309622 -340 309678 -284
rect 309250 -464 309306 -408
rect 309374 -464 309430 -408
rect 309498 -464 309554 -408
rect 309622 -464 309678 -408
rect 309250 -588 309306 -532
rect 309374 -588 309430 -532
rect 309498 -588 309554 -532
rect 309622 -588 309678 -532
rect 327250 4294 327306 4350
rect 327374 4294 327430 4350
rect 327498 4294 327554 4350
rect 327622 4294 327678 4350
rect 327250 4170 327306 4226
rect 327374 4170 327430 4226
rect 327498 4170 327554 4226
rect 327622 4170 327678 4226
rect 327250 4046 327306 4102
rect 327374 4046 327430 4102
rect 327498 4046 327554 4102
rect 327622 4046 327678 4102
rect 327250 3922 327306 3978
rect 327374 3922 327430 3978
rect 327498 3922 327554 3978
rect 327622 3922 327678 3978
rect 327250 -216 327306 -160
rect 327374 -216 327430 -160
rect 327498 -216 327554 -160
rect 327622 -216 327678 -160
rect 327250 -340 327306 -284
rect 327374 -340 327430 -284
rect 327498 -340 327554 -284
rect 327622 -340 327678 -284
rect 327250 -464 327306 -408
rect 327374 -464 327430 -408
rect 327498 -464 327554 -408
rect 327622 -464 327678 -408
rect 327250 -588 327306 -532
rect 327374 -588 327430 -532
rect 327498 -588 327554 -532
rect 327622 -588 327678 -532
rect 345250 4294 345306 4350
rect 345374 4294 345430 4350
rect 345498 4294 345554 4350
rect 345622 4294 345678 4350
rect 345250 4170 345306 4226
rect 345374 4170 345430 4226
rect 345498 4170 345554 4226
rect 345622 4170 345678 4226
rect 345250 4046 345306 4102
rect 345374 4046 345430 4102
rect 345498 4046 345554 4102
rect 345622 4046 345678 4102
rect 345250 3922 345306 3978
rect 345374 3922 345430 3978
rect 345498 3922 345554 3978
rect 345622 3922 345678 3978
rect 345250 -216 345306 -160
rect 345374 -216 345430 -160
rect 345498 -216 345554 -160
rect 345622 -216 345678 -160
rect 345250 -340 345306 -284
rect 345374 -340 345430 -284
rect 345498 -340 345554 -284
rect 345622 -340 345678 -284
rect 345250 -464 345306 -408
rect 345374 -464 345430 -408
rect 345498 -464 345554 -408
rect 345622 -464 345678 -408
rect 345250 -588 345306 -532
rect 345374 -588 345430 -532
rect 345498 -588 345554 -532
rect 345622 -588 345678 -532
rect 363250 4294 363306 4350
rect 363374 4294 363430 4350
rect 363498 4294 363554 4350
rect 363622 4294 363678 4350
rect 363250 4170 363306 4226
rect 363374 4170 363430 4226
rect 363498 4170 363554 4226
rect 363622 4170 363678 4226
rect 363250 4046 363306 4102
rect 363374 4046 363430 4102
rect 363498 4046 363554 4102
rect 363622 4046 363678 4102
rect 363250 3922 363306 3978
rect 363374 3922 363430 3978
rect 363498 3922 363554 3978
rect 363622 3922 363678 3978
rect 381250 148294 381306 148350
rect 381374 148294 381430 148350
rect 381498 148294 381554 148350
rect 381622 148294 381678 148350
rect 381250 148170 381306 148226
rect 381374 148170 381430 148226
rect 381498 148170 381554 148226
rect 381622 148170 381678 148226
rect 381250 148046 381306 148102
rect 381374 148046 381430 148102
rect 381498 148046 381554 148102
rect 381622 148046 381678 148102
rect 381250 147922 381306 147978
rect 381374 147922 381430 147978
rect 381498 147922 381554 147978
rect 381622 147922 381678 147978
rect 381250 130294 381306 130350
rect 381374 130294 381430 130350
rect 381498 130294 381554 130350
rect 381622 130294 381678 130350
rect 381250 130170 381306 130226
rect 381374 130170 381430 130226
rect 381498 130170 381554 130226
rect 381622 130170 381678 130226
rect 381250 130046 381306 130102
rect 381374 130046 381430 130102
rect 381498 130046 381554 130102
rect 381622 130046 381678 130102
rect 381250 129922 381306 129978
rect 381374 129922 381430 129978
rect 381498 129922 381554 129978
rect 381622 129922 381678 129978
rect 381250 112294 381306 112350
rect 381374 112294 381430 112350
rect 381498 112294 381554 112350
rect 381622 112294 381678 112350
rect 381250 112170 381306 112226
rect 381374 112170 381430 112226
rect 381498 112170 381554 112226
rect 381622 112170 381678 112226
rect 381250 112046 381306 112102
rect 381374 112046 381430 112102
rect 381498 112046 381554 112102
rect 381622 112046 381678 112102
rect 381250 111922 381306 111978
rect 381374 111922 381430 111978
rect 381498 111922 381554 111978
rect 381622 111922 381678 111978
rect 381250 94294 381306 94350
rect 381374 94294 381430 94350
rect 381498 94294 381554 94350
rect 381622 94294 381678 94350
rect 381250 94170 381306 94226
rect 381374 94170 381430 94226
rect 381498 94170 381554 94226
rect 381622 94170 381678 94226
rect 381250 94046 381306 94102
rect 381374 94046 381430 94102
rect 381498 94046 381554 94102
rect 381622 94046 381678 94102
rect 381250 93922 381306 93978
rect 381374 93922 381430 93978
rect 381498 93922 381554 93978
rect 381622 93922 381678 93978
rect 381250 76294 381306 76350
rect 381374 76294 381430 76350
rect 381498 76294 381554 76350
rect 381622 76294 381678 76350
rect 381250 76170 381306 76226
rect 381374 76170 381430 76226
rect 381498 76170 381554 76226
rect 381622 76170 381678 76226
rect 381250 76046 381306 76102
rect 381374 76046 381430 76102
rect 381498 76046 381554 76102
rect 381622 76046 381678 76102
rect 381250 75922 381306 75978
rect 381374 75922 381430 75978
rect 381498 75922 381554 75978
rect 381622 75922 381678 75978
rect 381250 58294 381306 58350
rect 381374 58294 381430 58350
rect 381498 58294 381554 58350
rect 381622 58294 381678 58350
rect 381250 58170 381306 58226
rect 381374 58170 381430 58226
rect 381498 58170 381554 58226
rect 381622 58170 381678 58226
rect 381250 58046 381306 58102
rect 381374 58046 381430 58102
rect 381498 58046 381554 58102
rect 381622 58046 381678 58102
rect 381250 57922 381306 57978
rect 381374 57922 381430 57978
rect 381498 57922 381554 57978
rect 381622 57922 381678 57978
rect 381250 40294 381306 40350
rect 381374 40294 381430 40350
rect 381498 40294 381554 40350
rect 381622 40294 381678 40350
rect 381250 40170 381306 40226
rect 381374 40170 381430 40226
rect 381498 40170 381554 40226
rect 381622 40170 381678 40226
rect 381250 40046 381306 40102
rect 381374 40046 381430 40102
rect 381498 40046 381554 40102
rect 381622 40046 381678 40102
rect 381250 39922 381306 39978
rect 381374 39922 381430 39978
rect 381498 39922 381554 39978
rect 381622 39922 381678 39978
rect 381250 22294 381306 22350
rect 381374 22294 381430 22350
rect 381498 22294 381554 22350
rect 381622 22294 381678 22350
rect 381250 22170 381306 22226
rect 381374 22170 381430 22226
rect 381498 22170 381554 22226
rect 381622 22170 381678 22226
rect 381250 22046 381306 22102
rect 381374 22046 381430 22102
rect 381498 22046 381554 22102
rect 381622 22046 381678 22102
rect 381250 21922 381306 21978
rect 381374 21922 381430 21978
rect 381498 21922 381554 21978
rect 381622 21922 381678 21978
rect 381250 4294 381306 4350
rect 381374 4294 381430 4350
rect 381498 4294 381554 4350
rect 381622 4294 381678 4350
rect 381250 4170 381306 4226
rect 381374 4170 381430 4226
rect 381498 4170 381554 4226
rect 381622 4170 381678 4226
rect 381250 4046 381306 4102
rect 381374 4046 381430 4102
rect 381498 4046 381554 4102
rect 381622 4046 381678 4102
rect 381250 3922 381306 3978
rect 381374 3922 381430 3978
rect 381498 3922 381554 3978
rect 381622 3922 381678 3978
rect 363250 -216 363306 -160
rect 363374 -216 363430 -160
rect 363498 -216 363554 -160
rect 363622 -216 363678 -160
rect 363250 -340 363306 -284
rect 363374 -340 363430 -284
rect 363498 -340 363554 -284
rect 363622 -340 363678 -284
rect 363250 -464 363306 -408
rect 363374 -464 363430 -408
rect 363498 -464 363554 -408
rect 363622 -464 363678 -408
rect 363250 -588 363306 -532
rect 363374 -588 363430 -532
rect 363498 -588 363554 -532
rect 363622 -588 363678 -532
rect 381250 -216 381306 -160
rect 381374 -216 381430 -160
rect 381498 -216 381554 -160
rect 381622 -216 381678 -160
rect 381250 -340 381306 -284
rect 381374 -340 381430 -284
rect 381498 -340 381554 -284
rect 381622 -340 381678 -284
rect 381250 -464 381306 -408
rect 381374 -464 381430 -408
rect 381498 -464 381554 -408
rect 381622 -464 381678 -408
rect 381250 -588 381306 -532
rect 381374 -588 381430 -532
rect 381498 -588 381554 -532
rect 381622 -588 381678 -532
rect 384970 598116 385026 598172
rect 385094 598116 385150 598172
rect 385218 598116 385274 598172
rect 385342 598116 385398 598172
rect 384970 597992 385026 598048
rect 385094 597992 385150 598048
rect 385218 597992 385274 598048
rect 385342 597992 385398 598048
rect 384970 597868 385026 597924
rect 385094 597868 385150 597924
rect 385218 597868 385274 597924
rect 385342 597868 385398 597924
rect 384970 597744 385026 597800
rect 385094 597744 385150 597800
rect 385218 597744 385274 597800
rect 385342 597744 385398 597800
rect 384970 586294 385026 586350
rect 385094 586294 385150 586350
rect 385218 586294 385274 586350
rect 385342 586294 385398 586350
rect 384970 586170 385026 586226
rect 385094 586170 385150 586226
rect 385218 586170 385274 586226
rect 385342 586170 385398 586226
rect 384970 586046 385026 586102
rect 385094 586046 385150 586102
rect 385218 586046 385274 586102
rect 385342 586046 385398 586102
rect 384970 585922 385026 585978
rect 385094 585922 385150 585978
rect 385218 585922 385274 585978
rect 385342 585922 385398 585978
rect 384970 568294 385026 568350
rect 385094 568294 385150 568350
rect 385218 568294 385274 568350
rect 385342 568294 385398 568350
rect 384970 568170 385026 568226
rect 385094 568170 385150 568226
rect 385218 568170 385274 568226
rect 385342 568170 385398 568226
rect 384970 568046 385026 568102
rect 385094 568046 385150 568102
rect 385218 568046 385274 568102
rect 385342 568046 385398 568102
rect 384970 567922 385026 567978
rect 385094 567922 385150 567978
rect 385218 567922 385274 567978
rect 385342 567922 385398 567978
rect 384970 550294 385026 550350
rect 385094 550294 385150 550350
rect 385218 550294 385274 550350
rect 385342 550294 385398 550350
rect 384970 550170 385026 550226
rect 385094 550170 385150 550226
rect 385218 550170 385274 550226
rect 385342 550170 385398 550226
rect 384970 550046 385026 550102
rect 385094 550046 385150 550102
rect 385218 550046 385274 550102
rect 385342 550046 385398 550102
rect 384970 549922 385026 549978
rect 385094 549922 385150 549978
rect 385218 549922 385274 549978
rect 385342 549922 385398 549978
rect 384970 532294 385026 532350
rect 385094 532294 385150 532350
rect 385218 532294 385274 532350
rect 385342 532294 385398 532350
rect 384970 532170 385026 532226
rect 385094 532170 385150 532226
rect 385218 532170 385274 532226
rect 385342 532170 385398 532226
rect 384970 532046 385026 532102
rect 385094 532046 385150 532102
rect 385218 532046 385274 532102
rect 385342 532046 385398 532102
rect 384970 531922 385026 531978
rect 385094 531922 385150 531978
rect 385218 531922 385274 531978
rect 385342 531922 385398 531978
rect 384970 514294 385026 514350
rect 385094 514294 385150 514350
rect 385218 514294 385274 514350
rect 385342 514294 385398 514350
rect 384970 514170 385026 514226
rect 385094 514170 385150 514226
rect 385218 514170 385274 514226
rect 385342 514170 385398 514226
rect 384970 514046 385026 514102
rect 385094 514046 385150 514102
rect 385218 514046 385274 514102
rect 385342 514046 385398 514102
rect 384970 513922 385026 513978
rect 385094 513922 385150 513978
rect 385218 513922 385274 513978
rect 385342 513922 385398 513978
rect 384970 496294 385026 496350
rect 385094 496294 385150 496350
rect 385218 496294 385274 496350
rect 385342 496294 385398 496350
rect 384970 496170 385026 496226
rect 385094 496170 385150 496226
rect 385218 496170 385274 496226
rect 385342 496170 385398 496226
rect 384970 496046 385026 496102
rect 385094 496046 385150 496102
rect 385218 496046 385274 496102
rect 385342 496046 385398 496102
rect 384970 495922 385026 495978
rect 385094 495922 385150 495978
rect 385218 495922 385274 495978
rect 385342 495922 385398 495978
rect 384970 478294 385026 478350
rect 385094 478294 385150 478350
rect 385218 478294 385274 478350
rect 385342 478294 385398 478350
rect 384970 478170 385026 478226
rect 385094 478170 385150 478226
rect 385218 478170 385274 478226
rect 385342 478170 385398 478226
rect 384970 478046 385026 478102
rect 385094 478046 385150 478102
rect 385218 478046 385274 478102
rect 385342 478046 385398 478102
rect 384970 477922 385026 477978
rect 385094 477922 385150 477978
rect 385218 477922 385274 477978
rect 385342 477922 385398 477978
rect 384970 460294 385026 460350
rect 385094 460294 385150 460350
rect 385218 460294 385274 460350
rect 385342 460294 385398 460350
rect 384970 460170 385026 460226
rect 385094 460170 385150 460226
rect 385218 460170 385274 460226
rect 385342 460170 385398 460226
rect 384970 460046 385026 460102
rect 385094 460046 385150 460102
rect 385218 460046 385274 460102
rect 385342 460046 385398 460102
rect 384970 459922 385026 459978
rect 385094 459922 385150 459978
rect 385218 459922 385274 459978
rect 385342 459922 385398 459978
rect 384970 442294 385026 442350
rect 385094 442294 385150 442350
rect 385218 442294 385274 442350
rect 385342 442294 385398 442350
rect 384970 442170 385026 442226
rect 385094 442170 385150 442226
rect 385218 442170 385274 442226
rect 385342 442170 385398 442226
rect 384970 442046 385026 442102
rect 385094 442046 385150 442102
rect 385218 442046 385274 442102
rect 385342 442046 385398 442102
rect 384970 441922 385026 441978
rect 385094 441922 385150 441978
rect 385218 441922 385274 441978
rect 385342 441922 385398 441978
rect 384970 424294 385026 424350
rect 385094 424294 385150 424350
rect 385218 424294 385274 424350
rect 385342 424294 385398 424350
rect 384970 424170 385026 424226
rect 385094 424170 385150 424226
rect 385218 424170 385274 424226
rect 385342 424170 385398 424226
rect 384970 424046 385026 424102
rect 385094 424046 385150 424102
rect 385218 424046 385274 424102
rect 385342 424046 385398 424102
rect 384970 423922 385026 423978
rect 385094 423922 385150 423978
rect 385218 423922 385274 423978
rect 385342 423922 385398 423978
rect 384970 406294 385026 406350
rect 385094 406294 385150 406350
rect 385218 406294 385274 406350
rect 385342 406294 385398 406350
rect 384970 406170 385026 406226
rect 385094 406170 385150 406226
rect 385218 406170 385274 406226
rect 385342 406170 385398 406226
rect 384970 406046 385026 406102
rect 385094 406046 385150 406102
rect 385218 406046 385274 406102
rect 385342 406046 385398 406102
rect 384970 405922 385026 405978
rect 385094 405922 385150 405978
rect 385218 405922 385274 405978
rect 385342 405922 385398 405978
rect 384970 388294 385026 388350
rect 385094 388294 385150 388350
rect 385218 388294 385274 388350
rect 385342 388294 385398 388350
rect 384970 388170 385026 388226
rect 385094 388170 385150 388226
rect 385218 388170 385274 388226
rect 385342 388170 385398 388226
rect 384970 388046 385026 388102
rect 385094 388046 385150 388102
rect 385218 388046 385274 388102
rect 385342 388046 385398 388102
rect 384970 387922 385026 387978
rect 385094 387922 385150 387978
rect 385218 387922 385274 387978
rect 385342 387922 385398 387978
rect 384970 370294 385026 370350
rect 385094 370294 385150 370350
rect 385218 370294 385274 370350
rect 385342 370294 385398 370350
rect 384970 370170 385026 370226
rect 385094 370170 385150 370226
rect 385218 370170 385274 370226
rect 385342 370170 385398 370226
rect 384970 370046 385026 370102
rect 385094 370046 385150 370102
rect 385218 370046 385274 370102
rect 385342 370046 385398 370102
rect 384970 369922 385026 369978
rect 385094 369922 385150 369978
rect 385218 369922 385274 369978
rect 385342 369922 385398 369978
rect 384970 352294 385026 352350
rect 385094 352294 385150 352350
rect 385218 352294 385274 352350
rect 385342 352294 385398 352350
rect 384970 352170 385026 352226
rect 385094 352170 385150 352226
rect 385218 352170 385274 352226
rect 385342 352170 385398 352226
rect 384970 352046 385026 352102
rect 385094 352046 385150 352102
rect 385218 352046 385274 352102
rect 385342 352046 385398 352102
rect 384970 351922 385026 351978
rect 385094 351922 385150 351978
rect 385218 351922 385274 351978
rect 385342 351922 385398 351978
rect 384970 334294 385026 334350
rect 385094 334294 385150 334350
rect 385218 334294 385274 334350
rect 385342 334294 385398 334350
rect 384970 334170 385026 334226
rect 385094 334170 385150 334226
rect 385218 334170 385274 334226
rect 385342 334170 385398 334226
rect 384970 334046 385026 334102
rect 385094 334046 385150 334102
rect 385218 334046 385274 334102
rect 385342 334046 385398 334102
rect 384970 333922 385026 333978
rect 385094 333922 385150 333978
rect 385218 333922 385274 333978
rect 385342 333922 385398 333978
rect 384970 316294 385026 316350
rect 385094 316294 385150 316350
rect 385218 316294 385274 316350
rect 385342 316294 385398 316350
rect 384970 316170 385026 316226
rect 385094 316170 385150 316226
rect 385218 316170 385274 316226
rect 385342 316170 385398 316226
rect 384970 316046 385026 316102
rect 385094 316046 385150 316102
rect 385218 316046 385274 316102
rect 385342 316046 385398 316102
rect 384970 315922 385026 315978
rect 385094 315922 385150 315978
rect 385218 315922 385274 315978
rect 385342 315922 385398 315978
rect 399250 597156 399306 597212
rect 399374 597156 399430 597212
rect 399498 597156 399554 597212
rect 399622 597156 399678 597212
rect 399250 597032 399306 597088
rect 399374 597032 399430 597088
rect 399498 597032 399554 597088
rect 399622 597032 399678 597088
rect 399250 596908 399306 596964
rect 399374 596908 399430 596964
rect 399498 596908 399554 596964
rect 399622 596908 399678 596964
rect 399250 596784 399306 596840
rect 399374 596784 399430 596840
rect 399498 596784 399554 596840
rect 399622 596784 399678 596840
rect 399250 580294 399306 580350
rect 399374 580294 399430 580350
rect 399498 580294 399554 580350
rect 399622 580294 399678 580350
rect 399250 580170 399306 580226
rect 399374 580170 399430 580226
rect 399498 580170 399554 580226
rect 399622 580170 399678 580226
rect 399250 580046 399306 580102
rect 399374 580046 399430 580102
rect 399498 580046 399554 580102
rect 399622 580046 399678 580102
rect 399250 579922 399306 579978
rect 399374 579922 399430 579978
rect 399498 579922 399554 579978
rect 399622 579922 399678 579978
rect 399250 562294 399306 562350
rect 399374 562294 399430 562350
rect 399498 562294 399554 562350
rect 399622 562294 399678 562350
rect 399250 562170 399306 562226
rect 399374 562170 399430 562226
rect 399498 562170 399554 562226
rect 399622 562170 399678 562226
rect 399250 562046 399306 562102
rect 399374 562046 399430 562102
rect 399498 562046 399554 562102
rect 399622 562046 399678 562102
rect 399250 561922 399306 561978
rect 399374 561922 399430 561978
rect 399498 561922 399554 561978
rect 399622 561922 399678 561978
rect 399250 544294 399306 544350
rect 399374 544294 399430 544350
rect 399498 544294 399554 544350
rect 399622 544294 399678 544350
rect 399250 544170 399306 544226
rect 399374 544170 399430 544226
rect 399498 544170 399554 544226
rect 399622 544170 399678 544226
rect 399250 544046 399306 544102
rect 399374 544046 399430 544102
rect 399498 544046 399554 544102
rect 399622 544046 399678 544102
rect 399250 543922 399306 543978
rect 399374 543922 399430 543978
rect 399498 543922 399554 543978
rect 399622 543922 399678 543978
rect 399250 526294 399306 526350
rect 399374 526294 399430 526350
rect 399498 526294 399554 526350
rect 399622 526294 399678 526350
rect 399250 526170 399306 526226
rect 399374 526170 399430 526226
rect 399498 526170 399554 526226
rect 399622 526170 399678 526226
rect 399250 526046 399306 526102
rect 399374 526046 399430 526102
rect 399498 526046 399554 526102
rect 399622 526046 399678 526102
rect 399250 525922 399306 525978
rect 399374 525922 399430 525978
rect 399498 525922 399554 525978
rect 399622 525922 399678 525978
rect 399250 508294 399306 508350
rect 399374 508294 399430 508350
rect 399498 508294 399554 508350
rect 399622 508294 399678 508350
rect 399250 508170 399306 508226
rect 399374 508170 399430 508226
rect 399498 508170 399554 508226
rect 399622 508170 399678 508226
rect 399250 508046 399306 508102
rect 399374 508046 399430 508102
rect 399498 508046 399554 508102
rect 399622 508046 399678 508102
rect 399250 507922 399306 507978
rect 399374 507922 399430 507978
rect 399498 507922 399554 507978
rect 399622 507922 399678 507978
rect 399250 490294 399306 490350
rect 399374 490294 399430 490350
rect 399498 490294 399554 490350
rect 399622 490294 399678 490350
rect 399250 490170 399306 490226
rect 399374 490170 399430 490226
rect 399498 490170 399554 490226
rect 399622 490170 399678 490226
rect 399250 490046 399306 490102
rect 399374 490046 399430 490102
rect 399498 490046 399554 490102
rect 399622 490046 399678 490102
rect 399250 489922 399306 489978
rect 399374 489922 399430 489978
rect 399498 489922 399554 489978
rect 399622 489922 399678 489978
rect 399250 472294 399306 472350
rect 399374 472294 399430 472350
rect 399498 472294 399554 472350
rect 399622 472294 399678 472350
rect 399250 472170 399306 472226
rect 399374 472170 399430 472226
rect 399498 472170 399554 472226
rect 399622 472170 399678 472226
rect 399250 472046 399306 472102
rect 399374 472046 399430 472102
rect 399498 472046 399554 472102
rect 399622 472046 399678 472102
rect 399250 471922 399306 471978
rect 399374 471922 399430 471978
rect 399498 471922 399554 471978
rect 399622 471922 399678 471978
rect 399250 454294 399306 454350
rect 399374 454294 399430 454350
rect 399498 454294 399554 454350
rect 399622 454294 399678 454350
rect 399250 454170 399306 454226
rect 399374 454170 399430 454226
rect 399498 454170 399554 454226
rect 399622 454170 399678 454226
rect 399250 454046 399306 454102
rect 399374 454046 399430 454102
rect 399498 454046 399554 454102
rect 399622 454046 399678 454102
rect 399250 453922 399306 453978
rect 399374 453922 399430 453978
rect 399498 453922 399554 453978
rect 399622 453922 399678 453978
rect 399250 436294 399306 436350
rect 399374 436294 399430 436350
rect 399498 436294 399554 436350
rect 399622 436294 399678 436350
rect 399250 436170 399306 436226
rect 399374 436170 399430 436226
rect 399498 436170 399554 436226
rect 399622 436170 399678 436226
rect 399250 436046 399306 436102
rect 399374 436046 399430 436102
rect 399498 436046 399554 436102
rect 399622 436046 399678 436102
rect 399250 435922 399306 435978
rect 399374 435922 399430 435978
rect 399498 435922 399554 435978
rect 399622 435922 399678 435978
rect 399250 418294 399306 418350
rect 399374 418294 399430 418350
rect 399498 418294 399554 418350
rect 399622 418294 399678 418350
rect 399250 418170 399306 418226
rect 399374 418170 399430 418226
rect 399498 418170 399554 418226
rect 399622 418170 399678 418226
rect 399250 418046 399306 418102
rect 399374 418046 399430 418102
rect 399498 418046 399554 418102
rect 399622 418046 399678 418102
rect 399250 417922 399306 417978
rect 399374 417922 399430 417978
rect 399498 417922 399554 417978
rect 399622 417922 399678 417978
rect 399250 400294 399306 400350
rect 399374 400294 399430 400350
rect 399498 400294 399554 400350
rect 399622 400294 399678 400350
rect 399250 400170 399306 400226
rect 399374 400170 399430 400226
rect 399498 400170 399554 400226
rect 399622 400170 399678 400226
rect 399250 400046 399306 400102
rect 399374 400046 399430 400102
rect 399498 400046 399554 400102
rect 399622 400046 399678 400102
rect 399250 399922 399306 399978
rect 399374 399922 399430 399978
rect 399498 399922 399554 399978
rect 399622 399922 399678 399978
rect 399250 382294 399306 382350
rect 399374 382294 399430 382350
rect 399498 382294 399554 382350
rect 399622 382294 399678 382350
rect 399250 382170 399306 382226
rect 399374 382170 399430 382226
rect 399498 382170 399554 382226
rect 399622 382170 399678 382226
rect 399250 382046 399306 382102
rect 399374 382046 399430 382102
rect 399498 382046 399554 382102
rect 399622 382046 399678 382102
rect 399250 381922 399306 381978
rect 399374 381922 399430 381978
rect 399498 381922 399554 381978
rect 399622 381922 399678 381978
rect 399250 364294 399306 364350
rect 399374 364294 399430 364350
rect 399498 364294 399554 364350
rect 399622 364294 399678 364350
rect 399250 364170 399306 364226
rect 399374 364170 399430 364226
rect 399498 364170 399554 364226
rect 399622 364170 399678 364226
rect 399250 364046 399306 364102
rect 399374 364046 399430 364102
rect 399498 364046 399554 364102
rect 399622 364046 399678 364102
rect 399250 363922 399306 363978
rect 399374 363922 399430 363978
rect 399498 363922 399554 363978
rect 399622 363922 399678 363978
rect 399250 346294 399306 346350
rect 399374 346294 399430 346350
rect 399498 346294 399554 346350
rect 399622 346294 399678 346350
rect 399250 346170 399306 346226
rect 399374 346170 399430 346226
rect 399498 346170 399554 346226
rect 399622 346170 399678 346226
rect 399250 346046 399306 346102
rect 399374 346046 399430 346102
rect 399498 346046 399554 346102
rect 399622 346046 399678 346102
rect 399250 345922 399306 345978
rect 399374 345922 399430 345978
rect 399498 345922 399554 345978
rect 399622 345922 399678 345978
rect 399250 328294 399306 328350
rect 399374 328294 399430 328350
rect 399498 328294 399554 328350
rect 399622 328294 399678 328350
rect 399250 328170 399306 328226
rect 399374 328170 399430 328226
rect 399498 328170 399554 328226
rect 399622 328170 399678 328226
rect 399250 328046 399306 328102
rect 399374 328046 399430 328102
rect 399498 328046 399554 328102
rect 399622 328046 399678 328102
rect 399250 327922 399306 327978
rect 399374 327922 399430 327978
rect 399498 327922 399554 327978
rect 399622 327922 399678 327978
rect 399250 310294 399306 310350
rect 399374 310294 399430 310350
rect 399498 310294 399554 310350
rect 399622 310294 399678 310350
rect 399250 310170 399306 310226
rect 399374 310170 399430 310226
rect 399498 310170 399554 310226
rect 399622 310170 399678 310226
rect 399250 310046 399306 310102
rect 399374 310046 399430 310102
rect 399498 310046 399554 310102
rect 399622 310046 399678 310102
rect 399250 309922 399306 309978
rect 399374 309922 399430 309978
rect 399498 309922 399554 309978
rect 399622 309922 399678 309978
rect 384970 298294 385026 298350
rect 385094 298294 385150 298350
rect 385218 298294 385274 298350
rect 385342 298294 385398 298350
rect 384970 298170 385026 298226
rect 385094 298170 385150 298226
rect 385218 298170 385274 298226
rect 385342 298170 385398 298226
rect 384970 298046 385026 298102
rect 385094 298046 385150 298102
rect 385218 298046 385274 298102
rect 385342 298046 385398 298102
rect 384970 297922 385026 297978
rect 385094 297922 385150 297978
rect 385218 297922 385274 297978
rect 385342 297922 385398 297978
rect 384970 280294 385026 280350
rect 385094 280294 385150 280350
rect 385218 280294 385274 280350
rect 385342 280294 385398 280350
rect 384970 280170 385026 280226
rect 385094 280170 385150 280226
rect 385218 280170 385274 280226
rect 385342 280170 385398 280226
rect 384970 280046 385026 280102
rect 385094 280046 385150 280102
rect 385218 280046 385274 280102
rect 385342 280046 385398 280102
rect 384970 279922 385026 279978
rect 385094 279922 385150 279978
rect 385218 279922 385274 279978
rect 385342 279922 385398 279978
rect 384970 262294 385026 262350
rect 385094 262294 385150 262350
rect 385218 262294 385274 262350
rect 385342 262294 385398 262350
rect 384970 262170 385026 262226
rect 385094 262170 385150 262226
rect 385218 262170 385274 262226
rect 385342 262170 385398 262226
rect 384970 262046 385026 262102
rect 385094 262046 385150 262102
rect 385218 262046 385274 262102
rect 385342 262046 385398 262102
rect 384970 261922 385026 261978
rect 385094 261922 385150 261978
rect 385218 261922 385274 261978
rect 385342 261922 385398 261978
rect 384970 244294 385026 244350
rect 385094 244294 385150 244350
rect 385218 244294 385274 244350
rect 385342 244294 385398 244350
rect 384970 244170 385026 244226
rect 385094 244170 385150 244226
rect 385218 244170 385274 244226
rect 385342 244170 385398 244226
rect 384970 244046 385026 244102
rect 385094 244046 385150 244102
rect 385218 244046 385274 244102
rect 385342 244046 385398 244102
rect 384970 243922 385026 243978
rect 385094 243922 385150 243978
rect 385218 243922 385274 243978
rect 385342 243922 385398 243978
rect 384970 226294 385026 226350
rect 385094 226294 385150 226350
rect 385218 226294 385274 226350
rect 385342 226294 385398 226350
rect 384970 226170 385026 226226
rect 385094 226170 385150 226226
rect 385218 226170 385274 226226
rect 385342 226170 385398 226226
rect 384970 226046 385026 226102
rect 385094 226046 385150 226102
rect 385218 226046 385274 226102
rect 385342 226046 385398 226102
rect 384970 225922 385026 225978
rect 385094 225922 385150 225978
rect 385218 225922 385274 225978
rect 385342 225922 385398 225978
rect 384970 208294 385026 208350
rect 385094 208294 385150 208350
rect 385218 208294 385274 208350
rect 385342 208294 385398 208350
rect 384970 208170 385026 208226
rect 385094 208170 385150 208226
rect 385218 208170 385274 208226
rect 385342 208170 385398 208226
rect 384970 208046 385026 208102
rect 385094 208046 385150 208102
rect 385218 208046 385274 208102
rect 385342 208046 385398 208102
rect 384970 207922 385026 207978
rect 385094 207922 385150 207978
rect 385218 207922 385274 207978
rect 385342 207922 385398 207978
rect 384970 190294 385026 190350
rect 385094 190294 385150 190350
rect 385218 190294 385274 190350
rect 385342 190294 385398 190350
rect 384970 190170 385026 190226
rect 385094 190170 385150 190226
rect 385218 190170 385274 190226
rect 385342 190170 385398 190226
rect 384970 190046 385026 190102
rect 385094 190046 385150 190102
rect 385218 190046 385274 190102
rect 385342 190046 385398 190102
rect 384970 189922 385026 189978
rect 385094 189922 385150 189978
rect 385218 189922 385274 189978
rect 385342 189922 385398 189978
rect 384970 172294 385026 172350
rect 385094 172294 385150 172350
rect 385218 172294 385274 172350
rect 385342 172294 385398 172350
rect 384970 172170 385026 172226
rect 385094 172170 385150 172226
rect 385218 172170 385274 172226
rect 385342 172170 385398 172226
rect 384970 172046 385026 172102
rect 385094 172046 385150 172102
rect 385218 172046 385274 172102
rect 385342 172046 385398 172102
rect 384970 171922 385026 171978
rect 385094 171922 385150 171978
rect 385218 171922 385274 171978
rect 385342 171922 385398 171978
rect 399250 292294 399306 292350
rect 399374 292294 399430 292350
rect 399498 292294 399554 292350
rect 399622 292294 399678 292350
rect 399250 292170 399306 292226
rect 399374 292170 399430 292226
rect 399498 292170 399554 292226
rect 399622 292170 399678 292226
rect 399250 292046 399306 292102
rect 399374 292046 399430 292102
rect 399498 292046 399554 292102
rect 399622 292046 399678 292102
rect 399250 291922 399306 291978
rect 399374 291922 399430 291978
rect 399498 291922 399554 291978
rect 399622 291922 399678 291978
rect 399250 274294 399306 274350
rect 399374 274294 399430 274350
rect 399498 274294 399554 274350
rect 399622 274294 399678 274350
rect 399250 274170 399306 274226
rect 399374 274170 399430 274226
rect 399498 274170 399554 274226
rect 399622 274170 399678 274226
rect 399250 274046 399306 274102
rect 399374 274046 399430 274102
rect 399498 274046 399554 274102
rect 399622 274046 399678 274102
rect 399250 273922 399306 273978
rect 399374 273922 399430 273978
rect 399498 273922 399554 273978
rect 399622 273922 399678 273978
rect 399250 256294 399306 256350
rect 399374 256294 399430 256350
rect 399498 256294 399554 256350
rect 399622 256294 399678 256350
rect 399250 256170 399306 256226
rect 399374 256170 399430 256226
rect 399498 256170 399554 256226
rect 399622 256170 399678 256226
rect 399250 256046 399306 256102
rect 399374 256046 399430 256102
rect 399498 256046 399554 256102
rect 399622 256046 399678 256102
rect 399250 255922 399306 255978
rect 399374 255922 399430 255978
rect 399498 255922 399554 255978
rect 399622 255922 399678 255978
rect 399250 238294 399306 238350
rect 399374 238294 399430 238350
rect 399498 238294 399554 238350
rect 399622 238294 399678 238350
rect 399250 238170 399306 238226
rect 399374 238170 399430 238226
rect 399498 238170 399554 238226
rect 399622 238170 399678 238226
rect 399250 238046 399306 238102
rect 399374 238046 399430 238102
rect 399498 238046 399554 238102
rect 399622 238046 399678 238102
rect 399250 237922 399306 237978
rect 399374 237922 399430 237978
rect 399498 237922 399554 237978
rect 399622 237922 399678 237978
rect 399250 220294 399306 220350
rect 399374 220294 399430 220350
rect 399498 220294 399554 220350
rect 399622 220294 399678 220350
rect 399250 220170 399306 220226
rect 399374 220170 399430 220226
rect 399498 220170 399554 220226
rect 399622 220170 399678 220226
rect 399250 220046 399306 220102
rect 399374 220046 399430 220102
rect 399498 220046 399554 220102
rect 399622 220046 399678 220102
rect 399250 219922 399306 219978
rect 399374 219922 399430 219978
rect 399498 219922 399554 219978
rect 399622 219922 399678 219978
rect 399250 202294 399306 202350
rect 399374 202294 399430 202350
rect 399498 202294 399554 202350
rect 399622 202294 399678 202350
rect 399250 202170 399306 202226
rect 399374 202170 399430 202226
rect 399498 202170 399554 202226
rect 399622 202170 399678 202226
rect 399250 202046 399306 202102
rect 399374 202046 399430 202102
rect 399498 202046 399554 202102
rect 399622 202046 399678 202102
rect 399250 201922 399306 201978
rect 399374 201922 399430 201978
rect 399498 201922 399554 201978
rect 399622 201922 399678 201978
rect 399250 184294 399306 184350
rect 399374 184294 399430 184350
rect 399498 184294 399554 184350
rect 399622 184294 399678 184350
rect 399250 184170 399306 184226
rect 399374 184170 399430 184226
rect 399498 184170 399554 184226
rect 399622 184170 399678 184226
rect 399250 184046 399306 184102
rect 399374 184046 399430 184102
rect 399498 184046 399554 184102
rect 399622 184046 399678 184102
rect 399250 183922 399306 183978
rect 399374 183922 399430 183978
rect 399498 183922 399554 183978
rect 399622 183922 399678 183978
rect 399250 166294 399306 166350
rect 399374 166294 399430 166350
rect 399498 166294 399554 166350
rect 399622 166294 399678 166350
rect 399250 166170 399306 166226
rect 399374 166170 399430 166226
rect 399498 166170 399554 166226
rect 399622 166170 399678 166226
rect 399250 166046 399306 166102
rect 399374 166046 399430 166102
rect 399498 166046 399554 166102
rect 399622 166046 399678 166102
rect 399250 165922 399306 165978
rect 399374 165922 399430 165978
rect 399498 165922 399554 165978
rect 399622 165922 399678 165978
rect 384970 154294 385026 154350
rect 385094 154294 385150 154350
rect 385218 154294 385274 154350
rect 385342 154294 385398 154350
rect 384970 154170 385026 154226
rect 385094 154170 385150 154226
rect 385218 154170 385274 154226
rect 385342 154170 385398 154226
rect 384970 154046 385026 154102
rect 385094 154046 385150 154102
rect 385218 154046 385274 154102
rect 385342 154046 385398 154102
rect 384970 153922 385026 153978
rect 385094 153922 385150 153978
rect 385218 153922 385274 153978
rect 385342 153922 385398 153978
rect 384970 136294 385026 136350
rect 385094 136294 385150 136350
rect 385218 136294 385274 136350
rect 385342 136294 385398 136350
rect 384970 136170 385026 136226
rect 385094 136170 385150 136226
rect 385218 136170 385274 136226
rect 385342 136170 385398 136226
rect 384970 136046 385026 136102
rect 385094 136046 385150 136102
rect 385218 136046 385274 136102
rect 385342 136046 385398 136102
rect 384970 135922 385026 135978
rect 385094 135922 385150 135978
rect 385218 135922 385274 135978
rect 385342 135922 385398 135978
rect 384970 118294 385026 118350
rect 385094 118294 385150 118350
rect 385218 118294 385274 118350
rect 385342 118294 385398 118350
rect 384970 118170 385026 118226
rect 385094 118170 385150 118226
rect 385218 118170 385274 118226
rect 385342 118170 385398 118226
rect 384970 118046 385026 118102
rect 385094 118046 385150 118102
rect 385218 118046 385274 118102
rect 385342 118046 385398 118102
rect 384970 117922 385026 117978
rect 385094 117922 385150 117978
rect 385218 117922 385274 117978
rect 385342 117922 385398 117978
rect 384970 100294 385026 100350
rect 385094 100294 385150 100350
rect 385218 100294 385274 100350
rect 385342 100294 385398 100350
rect 384970 100170 385026 100226
rect 385094 100170 385150 100226
rect 385218 100170 385274 100226
rect 385342 100170 385398 100226
rect 384970 100046 385026 100102
rect 385094 100046 385150 100102
rect 385218 100046 385274 100102
rect 385342 100046 385398 100102
rect 384970 99922 385026 99978
rect 385094 99922 385150 99978
rect 385218 99922 385274 99978
rect 385342 99922 385398 99978
rect 384970 82294 385026 82350
rect 385094 82294 385150 82350
rect 385218 82294 385274 82350
rect 385342 82294 385398 82350
rect 384970 82170 385026 82226
rect 385094 82170 385150 82226
rect 385218 82170 385274 82226
rect 385342 82170 385398 82226
rect 384970 82046 385026 82102
rect 385094 82046 385150 82102
rect 385218 82046 385274 82102
rect 385342 82046 385398 82102
rect 384970 81922 385026 81978
rect 385094 81922 385150 81978
rect 385218 81922 385274 81978
rect 385342 81922 385398 81978
rect 384970 64294 385026 64350
rect 385094 64294 385150 64350
rect 385218 64294 385274 64350
rect 385342 64294 385398 64350
rect 384970 64170 385026 64226
rect 385094 64170 385150 64226
rect 385218 64170 385274 64226
rect 385342 64170 385398 64226
rect 384970 64046 385026 64102
rect 385094 64046 385150 64102
rect 385218 64046 385274 64102
rect 385342 64046 385398 64102
rect 384970 63922 385026 63978
rect 385094 63922 385150 63978
rect 385218 63922 385274 63978
rect 385342 63922 385398 63978
rect 384970 46294 385026 46350
rect 385094 46294 385150 46350
rect 385218 46294 385274 46350
rect 385342 46294 385398 46350
rect 384970 46170 385026 46226
rect 385094 46170 385150 46226
rect 385218 46170 385274 46226
rect 385342 46170 385398 46226
rect 384970 46046 385026 46102
rect 385094 46046 385150 46102
rect 385218 46046 385274 46102
rect 385342 46046 385398 46102
rect 384970 45922 385026 45978
rect 385094 45922 385150 45978
rect 385218 45922 385274 45978
rect 385342 45922 385398 45978
rect 384970 28294 385026 28350
rect 385094 28294 385150 28350
rect 385218 28294 385274 28350
rect 385342 28294 385398 28350
rect 384970 28170 385026 28226
rect 385094 28170 385150 28226
rect 385218 28170 385274 28226
rect 385342 28170 385398 28226
rect 384970 28046 385026 28102
rect 385094 28046 385150 28102
rect 385218 28046 385274 28102
rect 385342 28046 385398 28102
rect 384970 27922 385026 27978
rect 385094 27922 385150 27978
rect 385218 27922 385274 27978
rect 385342 27922 385398 27978
rect 384970 10294 385026 10350
rect 385094 10294 385150 10350
rect 385218 10294 385274 10350
rect 385342 10294 385398 10350
rect 384970 10170 385026 10226
rect 385094 10170 385150 10226
rect 385218 10170 385274 10226
rect 385342 10170 385398 10226
rect 384970 10046 385026 10102
rect 385094 10046 385150 10102
rect 385218 10046 385274 10102
rect 385342 10046 385398 10102
rect 384970 9922 385026 9978
rect 385094 9922 385150 9978
rect 385218 9922 385274 9978
rect 385342 9922 385398 9978
rect 384970 -1176 385026 -1120
rect 385094 -1176 385150 -1120
rect 385218 -1176 385274 -1120
rect 385342 -1176 385398 -1120
rect 384970 -1300 385026 -1244
rect 385094 -1300 385150 -1244
rect 385218 -1300 385274 -1244
rect 385342 -1300 385398 -1244
rect 384970 -1424 385026 -1368
rect 385094 -1424 385150 -1368
rect 385218 -1424 385274 -1368
rect 385342 -1424 385398 -1368
rect 384970 -1548 385026 -1492
rect 385094 -1548 385150 -1492
rect 385218 -1548 385274 -1492
rect 385342 -1548 385398 -1492
rect 399250 148294 399306 148350
rect 399374 148294 399430 148350
rect 399498 148294 399554 148350
rect 399622 148294 399678 148350
rect 399250 148170 399306 148226
rect 399374 148170 399430 148226
rect 399498 148170 399554 148226
rect 399622 148170 399678 148226
rect 399250 148046 399306 148102
rect 399374 148046 399430 148102
rect 399498 148046 399554 148102
rect 399622 148046 399678 148102
rect 399250 147922 399306 147978
rect 399374 147922 399430 147978
rect 399498 147922 399554 147978
rect 399622 147922 399678 147978
rect 399250 130294 399306 130350
rect 399374 130294 399430 130350
rect 399498 130294 399554 130350
rect 399622 130294 399678 130350
rect 399250 130170 399306 130226
rect 399374 130170 399430 130226
rect 399498 130170 399554 130226
rect 399622 130170 399678 130226
rect 399250 130046 399306 130102
rect 399374 130046 399430 130102
rect 399498 130046 399554 130102
rect 399622 130046 399678 130102
rect 399250 129922 399306 129978
rect 399374 129922 399430 129978
rect 399498 129922 399554 129978
rect 399622 129922 399678 129978
rect 399250 112294 399306 112350
rect 399374 112294 399430 112350
rect 399498 112294 399554 112350
rect 399622 112294 399678 112350
rect 399250 112170 399306 112226
rect 399374 112170 399430 112226
rect 399498 112170 399554 112226
rect 399622 112170 399678 112226
rect 399250 112046 399306 112102
rect 399374 112046 399430 112102
rect 399498 112046 399554 112102
rect 399622 112046 399678 112102
rect 399250 111922 399306 111978
rect 399374 111922 399430 111978
rect 399498 111922 399554 111978
rect 399622 111922 399678 111978
rect 399250 94294 399306 94350
rect 399374 94294 399430 94350
rect 399498 94294 399554 94350
rect 399622 94294 399678 94350
rect 399250 94170 399306 94226
rect 399374 94170 399430 94226
rect 399498 94170 399554 94226
rect 399622 94170 399678 94226
rect 399250 94046 399306 94102
rect 399374 94046 399430 94102
rect 399498 94046 399554 94102
rect 399622 94046 399678 94102
rect 399250 93922 399306 93978
rect 399374 93922 399430 93978
rect 399498 93922 399554 93978
rect 399622 93922 399678 93978
rect 399250 76294 399306 76350
rect 399374 76294 399430 76350
rect 399498 76294 399554 76350
rect 399622 76294 399678 76350
rect 399250 76170 399306 76226
rect 399374 76170 399430 76226
rect 399498 76170 399554 76226
rect 399622 76170 399678 76226
rect 399250 76046 399306 76102
rect 399374 76046 399430 76102
rect 399498 76046 399554 76102
rect 399622 76046 399678 76102
rect 399250 75922 399306 75978
rect 399374 75922 399430 75978
rect 399498 75922 399554 75978
rect 399622 75922 399678 75978
rect 399250 58294 399306 58350
rect 399374 58294 399430 58350
rect 399498 58294 399554 58350
rect 399622 58294 399678 58350
rect 399250 58170 399306 58226
rect 399374 58170 399430 58226
rect 399498 58170 399554 58226
rect 399622 58170 399678 58226
rect 399250 58046 399306 58102
rect 399374 58046 399430 58102
rect 399498 58046 399554 58102
rect 399622 58046 399678 58102
rect 399250 57922 399306 57978
rect 399374 57922 399430 57978
rect 399498 57922 399554 57978
rect 399622 57922 399678 57978
rect 399250 40294 399306 40350
rect 399374 40294 399430 40350
rect 399498 40294 399554 40350
rect 399622 40294 399678 40350
rect 399250 40170 399306 40226
rect 399374 40170 399430 40226
rect 399498 40170 399554 40226
rect 399622 40170 399678 40226
rect 399250 40046 399306 40102
rect 399374 40046 399430 40102
rect 399498 40046 399554 40102
rect 399622 40046 399678 40102
rect 399250 39922 399306 39978
rect 399374 39922 399430 39978
rect 399498 39922 399554 39978
rect 399622 39922 399678 39978
rect 399250 22294 399306 22350
rect 399374 22294 399430 22350
rect 399498 22294 399554 22350
rect 399622 22294 399678 22350
rect 399250 22170 399306 22226
rect 399374 22170 399430 22226
rect 399498 22170 399554 22226
rect 399622 22170 399678 22226
rect 399250 22046 399306 22102
rect 399374 22046 399430 22102
rect 399498 22046 399554 22102
rect 399622 22046 399678 22102
rect 399250 21922 399306 21978
rect 399374 21922 399430 21978
rect 399498 21922 399554 21978
rect 399622 21922 399678 21978
rect 399250 4294 399306 4350
rect 399374 4294 399430 4350
rect 399498 4294 399554 4350
rect 399622 4294 399678 4350
rect 399250 4170 399306 4226
rect 399374 4170 399430 4226
rect 399498 4170 399554 4226
rect 399622 4170 399678 4226
rect 399250 4046 399306 4102
rect 399374 4046 399430 4102
rect 399498 4046 399554 4102
rect 399622 4046 399678 4102
rect 399250 3922 399306 3978
rect 399374 3922 399430 3978
rect 399498 3922 399554 3978
rect 399622 3922 399678 3978
rect 399250 -216 399306 -160
rect 399374 -216 399430 -160
rect 399498 -216 399554 -160
rect 399622 -216 399678 -160
rect 399250 -340 399306 -284
rect 399374 -340 399430 -284
rect 399498 -340 399554 -284
rect 399622 -340 399678 -284
rect 399250 -464 399306 -408
rect 399374 -464 399430 -408
rect 399498 -464 399554 -408
rect 399622 -464 399678 -408
rect 399250 -588 399306 -532
rect 399374 -588 399430 -532
rect 399498 -588 399554 -532
rect 399622 -588 399678 -532
rect 402970 598116 403026 598172
rect 403094 598116 403150 598172
rect 403218 598116 403274 598172
rect 403342 598116 403398 598172
rect 402970 597992 403026 598048
rect 403094 597992 403150 598048
rect 403218 597992 403274 598048
rect 403342 597992 403398 598048
rect 402970 597868 403026 597924
rect 403094 597868 403150 597924
rect 403218 597868 403274 597924
rect 403342 597868 403398 597924
rect 402970 597744 403026 597800
rect 403094 597744 403150 597800
rect 403218 597744 403274 597800
rect 403342 597744 403398 597800
rect 402970 586294 403026 586350
rect 403094 586294 403150 586350
rect 403218 586294 403274 586350
rect 403342 586294 403398 586350
rect 402970 586170 403026 586226
rect 403094 586170 403150 586226
rect 403218 586170 403274 586226
rect 403342 586170 403398 586226
rect 402970 586046 403026 586102
rect 403094 586046 403150 586102
rect 403218 586046 403274 586102
rect 403342 586046 403398 586102
rect 402970 585922 403026 585978
rect 403094 585922 403150 585978
rect 403218 585922 403274 585978
rect 403342 585922 403398 585978
rect 402970 568294 403026 568350
rect 403094 568294 403150 568350
rect 403218 568294 403274 568350
rect 403342 568294 403398 568350
rect 402970 568170 403026 568226
rect 403094 568170 403150 568226
rect 403218 568170 403274 568226
rect 403342 568170 403398 568226
rect 402970 568046 403026 568102
rect 403094 568046 403150 568102
rect 403218 568046 403274 568102
rect 403342 568046 403398 568102
rect 402970 567922 403026 567978
rect 403094 567922 403150 567978
rect 403218 567922 403274 567978
rect 403342 567922 403398 567978
rect 402970 550294 403026 550350
rect 403094 550294 403150 550350
rect 403218 550294 403274 550350
rect 403342 550294 403398 550350
rect 402970 550170 403026 550226
rect 403094 550170 403150 550226
rect 403218 550170 403274 550226
rect 403342 550170 403398 550226
rect 402970 550046 403026 550102
rect 403094 550046 403150 550102
rect 403218 550046 403274 550102
rect 403342 550046 403398 550102
rect 402970 549922 403026 549978
rect 403094 549922 403150 549978
rect 403218 549922 403274 549978
rect 403342 549922 403398 549978
rect 402970 532294 403026 532350
rect 403094 532294 403150 532350
rect 403218 532294 403274 532350
rect 403342 532294 403398 532350
rect 402970 532170 403026 532226
rect 403094 532170 403150 532226
rect 403218 532170 403274 532226
rect 403342 532170 403398 532226
rect 402970 532046 403026 532102
rect 403094 532046 403150 532102
rect 403218 532046 403274 532102
rect 403342 532046 403398 532102
rect 402970 531922 403026 531978
rect 403094 531922 403150 531978
rect 403218 531922 403274 531978
rect 403342 531922 403398 531978
rect 402970 514294 403026 514350
rect 403094 514294 403150 514350
rect 403218 514294 403274 514350
rect 403342 514294 403398 514350
rect 402970 514170 403026 514226
rect 403094 514170 403150 514226
rect 403218 514170 403274 514226
rect 403342 514170 403398 514226
rect 402970 514046 403026 514102
rect 403094 514046 403150 514102
rect 403218 514046 403274 514102
rect 403342 514046 403398 514102
rect 402970 513922 403026 513978
rect 403094 513922 403150 513978
rect 403218 513922 403274 513978
rect 403342 513922 403398 513978
rect 402970 496294 403026 496350
rect 403094 496294 403150 496350
rect 403218 496294 403274 496350
rect 403342 496294 403398 496350
rect 402970 496170 403026 496226
rect 403094 496170 403150 496226
rect 403218 496170 403274 496226
rect 403342 496170 403398 496226
rect 402970 496046 403026 496102
rect 403094 496046 403150 496102
rect 403218 496046 403274 496102
rect 403342 496046 403398 496102
rect 402970 495922 403026 495978
rect 403094 495922 403150 495978
rect 403218 495922 403274 495978
rect 403342 495922 403398 495978
rect 402970 478294 403026 478350
rect 403094 478294 403150 478350
rect 403218 478294 403274 478350
rect 403342 478294 403398 478350
rect 402970 478170 403026 478226
rect 403094 478170 403150 478226
rect 403218 478170 403274 478226
rect 403342 478170 403398 478226
rect 402970 478046 403026 478102
rect 403094 478046 403150 478102
rect 403218 478046 403274 478102
rect 403342 478046 403398 478102
rect 402970 477922 403026 477978
rect 403094 477922 403150 477978
rect 403218 477922 403274 477978
rect 403342 477922 403398 477978
rect 402970 460294 403026 460350
rect 403094 460294 403150 460350
rect 403218 460294 403274 460350
rect 403342 460294 403398 460350
rect 402970 460170 403026 460226
rect 403094 460170 403150 460226
rect 403218 460170 403274 460226
rect 403342 460170 403398 460226
rect 402970 460046 403026 460102
rect 403094 460046 403150 460102
rect 403218 460046 403274 460102
rect 403342 460046 403398 460102
rect 402970 459922 403026 459978
rect 403094 459922 403150 459978
rect 403218 459922 403274 459978
rect 403342 459922 403398 459978
rect 417250 597156 417306 597212
rect 417374 597156 417430 597212
rect 417498 597156 417554 597212
rect 417622 597156 417678 597212
rect 417250 597032 417306 597088
rect 417374 597032 417430 597088
rect 417498 597032 417554 597088
rect 417622 597032 417678 597088
rect 417250 596908 417306 596964
rect 417374 596908 417430 596964
rect 417498 596908 417554 596964
rect 417622 596908 417678 596964
rect 417250 596784 417306 596840
rect 417374 596784 417430 596840
rect 417498 596784 417554 596840
rect 417622 596784 417678 596840
rect 417250 580294 417306 580350
rect 417374 580294 417430 580350
rect 417498 580294 417554 580350
rect 417622 580294 417678 580350
rect 417250 580170 417306 580226
rect 417374 580170 417430 580226
rect 417498 580170 417554 580226
rect 417622 580170 417678 580226
rect 417250 580046 417306 580102
rect 417374 580046 417430 580102
rect 417498 580046 417554 580102
rect 417622 580046 417678 580102
rect 417250 579922 417306 579978
rect 417374 579922 417430 579978
rect 417498 579922 417554 579978
rect 417622 579922 417678 579978
rect 417250 562294 417306 562350
rect 417374 562294 417430 562350
rect 417498 562294 417554 562350
rect 417622 562294 417678 562350
rect 417250 562170 417306 562226
rect 417374 562170 417430 562226
rect 417498 562170 417554 562226
rect 417622 562170 417678 562226
rect 417250 562046 417306 562102
rect 417374 562046 417430 562102
rect 417498 562046 417554 562102
rect 417622 562046 417678 562102
rect 417250 561922 417306 561978
rect 417374 561922 417430 561978
rect 417498 561922 417554 561978
rect 417622 561922 417678 561978
rect 417250 544294 417306 544350
rect 417374 544294 417430 544350
rect 417498 544294 417554 544350
rect 417622 544294 417678 544350
rect 417250 544170 417306 544226
rect 417374 544170 417430 544226
rect 417498 544170 417554 544226
rect 417622 544170 417678 544226
rect 417250 544046 417306 544102
rect 417374 544046 417430 544102
rect 417498 544046 417554 544102
rect 417622 544046 417678 544102
rect 417250 543922 417306 543978
rect 417374 543922 417430 543978
rect 417498 543922 417554 543978
rect 417622 543922 417678 543978
rect 417250 526294 417306 526350
rect 417374 526294 417430 526350
rect 417498 526294 417554 526350
rect 417622 526294 417678 526350
rect 417250 526170 417306 526226
rect 417374 526170 417430 526226
rect 417498 526170 417554 526226
rect 417622 526170 417678 526226
rect 417250 526046 417306 526102
rect 417374 526046 417430 526102
rect 417498 526046 417554 526102
rect 417622 526046 417678 526102
rect 417250 525922 417306 525978
rect 417374 525922 417430 525978
rect 417498 525922 417554 525978
rect 417622 525922 417678 525978
rect 417250 508294 417306 508350
rect 417374 508294 417430 508350
rect 417498 508294 417554 508350
rect 417622 508294 417678 508350
rect 417250 508170 417306 508226
rect 417374 508170 417430 508226
rect 417498 508170 417554 508226
rect 417622 508170 417678 508226
rect 417250 508046 417306 508102
rect 417374 508046 417430 508102
rect 417498 508046 417554 508102
rect 417622 508046 417678 508102
rect 417250 507922 417306 507978
rect 417374 507922 417430 507978
rect 417498 507922 417554 507978
rect 417622 507922 417678 507978
rect 417250 490294 417306 490350
rect 417374 490294 417430 490350
rect 417498 490294 417554 490350
rect 417622 490294 417678 490350
rect 417250 490170 417306 490226
rect 417374 490170 417430 490226
rect 417498 490170 417554 490226
rect 417622 490170 417678 490226
rect 417250 490046 417306 490102
rect 417374 490046 417430 490102
rect 417498 490046 417554 490102
rect 417622 490046 417678 490102
rect 417250 489922 417306 489978
rect 417374 489922 417430 489978
rect 417498 489922 417554 489978
rect 417622 489922 417678 489978
rect 417250 472294 417306 472350
rect 417374 472294 417430 472350
rect 417498 472294 417554 472350
rect 417622 472294 417678 472350
rect 417250 472170 417306 472226
rect 417374 472170 417430 472226
rect 417498 472170 417554 472226
rect 417622 472170 417678 472226
rect 417250 472046 417306 472102
rect 417374 472046 417430 472102
rect 417498 472046 417554 472102
rect 417622 472046 417678 472102
rect 417250 471922 417306 471978
rect 417374 471922 417430 471978
rect 417498 471922 417554 471978
rect 417622 471922 417678 471978
rect 420970 598116 421026 598172
rect 421094 598116 421150 598172
rect 421218 598116 421274 598172
rect 421342 598116 421398 598172
rect 420970 597992 421026 598048
rect 421094 597992 421150 598048
rect 421218 597992 421274 598048
rect 421342 597992 421398 598048
rect 420970 597868 421026 597924
rect 421094 597868 421150 597924
rect 421218 597868 421274 597924
rect 421342 597868 421398 597924
rect 420970 597744 421026 597800
rect 421094 597744 421150 597800
rect 421218 597744 421274 597800
rect 421342 597744 421398 597800
rect 420970 586294 421026 586350
rect 421094 586294 421150 586350
rect 421218 586294 421274 586350
rect 421342 586294 421398 586350
rect 420970 586170 421026 586226
rect 421094 586170 421150 586226
rect 421218 586170 421274 586226
rect 421342 586170 421398 586226
rect 420970 586046 421026 586102
rect 421094 586046 421150 586102
rect 421218 586046 421274 586102
rect 421342 586046 421398 586102
rect 420970 585922 421026 585978
rect 421094 585922 421150 585978
rect 421218 585922 421274 585978
rect 421342 585922 421398 585978
rect 420970 568294 421026 568350
rect 421094 568294 421150 568350
rect 421218 568294 421274 568350
rect 421342 568294 421398 568350
rect 420970 568170 421026 568226
rect 421094 568170 421150 568226
rect 421218 568170 421274 568226
rect 421342 568170 421398 568226
rect 420970 568046 421026 568102
rect 421094 568046 421150 568102
rect 421218 568046 421274 568102
rect 421342 568046 421398 568102
rect 420970 567922 421026 567978
rect 421094 567922 421150 567978
rect 421218 567922 421274 567978
rect 421342 567922 421398 567978
rect 420970 550294 421026 550350
rect 421094 550294 421150 550350
rect 421218 550294 421274 550350
rect 421342 550294 421398 550350
rect 420970 550170 421026 550226
rect 421094 550170 421150 550226
rect 421218 550170 421274 550226
rect 421342 550170 421398 550226
rect 420970 550046 421026 550102
rect 421094 550046 421150 550102
rect 421218 550046 421274 550102
rect 421342 550046 421398 550102
rect 420970 549922 421026 549978
rect 421094 549922 421150 549978
rect 421218 549922 421274 549978
rect 421342 549922 421398 549978
rect 420970 532294 421026 532350
rect 421094 532294 421150 532350
rect 421218 532294 421274 532350
rect 421342 532294 421398 532350
rect 420970 532170 421026 532226
rect 421094 532170 421150 532226
rect 421218 532170 421274 532226
rect 421342 532170 421398 532226
rect 420970 532046 421026 532102
rect 421094 532046 421150 532102
rect 421218 532046 421274 532102
rect 421342 532046 421398 532102
rect 420970 531922 421026 531978
rect 421094 531922 421150 531978
rect 421218 531922 421274 531978
rect 421342 531922 421398 531978
rect 420970 514294 421026 514350
rect 421094 514294 421150 514350
rect 421218 514294 421274 514350
rect 421342 514294 421398 514350
rect 420970 514170 421026 514226
rect 421094 514170 421150 514226
rect 421218 514170 421274 514226
rect 421342 514170 421398 514226
rect 420970 514046 421026 514102
rect 421094 514046 421150 514102
rect 421218 514046 421274 514102
rect 421342 514046 421398 514102
rect 420970 513922 421026 513978
rect 421094 513922 421150 513978
rect 421218 513922 421274 513978
rect 421342 513922 421398 513978
rect 420970 496294 421026 496350
rect 421094 496294 421150 496350
rect 421218 496294 421274 496350
rect 421342 496294 421398 496350
rect 420970 496170 421026 496226
rect 421094 496170 421150 496226
rect 421218 496170 421274 496226
rect 421342 496170 421398 496226
rect 420970 496046 421026 496102
rect 421094 496046 421150 496102
rect 421218 496046 421274 496102
rect 421342 496046 421398 496102
rect 420970 495922 421026 495978
rect 421094 495922 421150 495978
rect 421218 495922 421274 495978
rect 421342 495922 421398 495978
rect 420970 478294 421026 478350
rect 421094 478294 421150 478350
rect 421218 478294 421274 478350
rect 421342 478294 421398 478350
rect 420970 478170 421026 478226
rect 421094 478170 421150 478226
rect 421218 478170 421274 478226
rect 421342 478170 421398 478226
rect 420970 478046 421026 478102
rect 421094 478046 421150 478102
rect 421218 478046 421274 478102
rect 421342 478046 421398 478102
rect 420970 477922 421026 477978
rect 421094 477922 421150 477978
rect 421218 477922 421274 477978
rect 421342 477922 421398 477978
rect 420970 460294 421026 460350
rect 421094 460294 421150 460350
rect 421218 460294 421274 460350
rect 421342 460294 421398 460350
rect 420970 460170 421026 460226
rect 421094 460170 421150 460226
rect 421218 460170 421274 460226
rect 421342 460170 421398 460226
rect 420970 460046 421026 460102
rect 421094 460046 421150 460102
rect 421218 460046 421274 460102
rect 421342 460046 421398 460102
rect 420970 459922 421026 459978
rect 421094 459922 421150 459978
rect 421218 459922 421274 459978
rect 421342 459922 421398 459978
rect 435250 597156 435306 597212
rect 435374 597156 435430 597212
rect 435498 597156 435554 597212
rect 435622 597156 435678 597212
rect 435250 597032 435306 597088
rect 435374 597032 435430 597088
rect 435498 597032 435554 597088
rect 435622 597032 435678 597088
rect 435250 596908 435306 596964
rect 435374 596908 435430 596964
rect 435498 596908 435554 596964
rect 435622 596908 435678 596964
rect 435250 596784 435306 596840
rect 435374 596784 435430 596840
rect 435498 596784 435554 596840
rect 435622 596784 435678 596840
rect 435250 580294 435306 580350
rect 435374 580294 435430 580350
rect 435498 580294 435554 580350
rect 435622 580294 435678 580350
rect 435250 580170 435306 580226
rect 435374 580170 435430 580226
rect 435498 580170 435554 580226
rect 435622 580170 435678 580226
rect 435250 580046 435306 580102
rect 435374 580046 435430 580102
rect 435498 580046 435554 580102
rect 435622 580046 435678 580102
rect 435250 579922 435306 579978
rect 435374 579922 435430 579978
rect 435498 579922 435554 579978
rect 435622 579922 435678 579978
rect 435250 562294 435306 562350
rect 435374 562294 435430 562350
rect 435498 562294 435554 562350
rect 435622 562294 435678 562350
rect 435250 562170 435306 562226
rect 435374 562170 435430 562226
rect 435498 562170 435554 562226
rect 435622 562170 435678 562226
rect 435250 562046 435306 562102
rect 435374 562046 435430 562102
rect 435498 562046 435554 562102
rect 435622 562046 435678 562102
rect 435250 561922 435306 561978
rect 435374 561922 435430 561978
rect 435498 561922 435554 561978
rect 435622 561922 435678 561978
rect 435250 544294 435306 544350
rect 435374 544294 435430 544350
rect 435498 544294 435554 544350
rect 435622 544294 435678 544350
rect 435250 544170 435306 544226
rect 435374 544170 435430 544226
rect 435498 544170 435554 544226
rect 435622 544170 435678 544226
rect 435250 544046 435306 544102
rect 435374 544046 435430 544102
rect 435498 544046 435554 544102
rect 435622 544046 435678 544102
rect 435250 543922 435306 543978
rect 435374 543922 435430 543978
rect 435498 543922 435554 543978
rect 435622 543922 435678 543978
rect 435250 526294 435306 526350
rect 435374 526294 435430 526350
rect 435498 526294 435554 526350
rect 435622 526294 435678 526350
rect 435250 526170 435306 526226
rect 435374 526170 435430 526226
rect 435498 526170 435554 526226
rect 435622 526170 435678 526226
rect 435250 526046 435306 526102
rect 435374 526046 435430 526102
rect 435498 526046 435554 526102
rect 435622 526046 435678 526102
rect 435250 525922 435306 525978
rect 435374 525922 435430 525978
rect 435498 525922 435554 525978
rect 435622 525922 435678 525978
rect 435250 508294 435306 508350
rect 435374 508294 435430 508350
rect 435498 508294 435554 508350
rect 435622 508294 435678 508350
rect 435250 508170 435306 508226
rect 435374 508170 435430 508226
rect 435498 508170 435554 508226
rect 435622 508170 435678 508226
rect 435250 508046 435306 508102
rect 435374 508046 435430 508102
rect 435498 508046 435554 508102
rect 435622 508046 435678 508102
rect 435250 507922 435306 507978
rect 435374 507922 435430 507978
rect 435498 507922 435554 507978
rect 435622 507922 435678 507978
rect 435250 490294 435306 490350
rect 435374 490294 435430 490350
rect 435498 490294 435554 490350
rect 435622 490294 435678 490350
rect 435250 490170 435306 490226
rect 435374 490170 435430 490226
rect 435498 490170 435554 490226
rect 435622 490170 435678 490226
rect 435250 490046 435306 490102
rect 435374 490046 435430 490102
rect 435498 490046 435554 490102
rect 435622 490046 435678 490102
rect 435250 489922 435306 489978
rect 435374 489922 435430 489978
rect 435498 489922 435554 489978
rect 435622 489922 435678 489978
rect 435250 472294 435306 472350
rect 435374 472294 435430 472350
rect 435498 472294 435554 472350
rect 435622 472294 435678 472350
rect 435250 472170 435306 472226
rect 435374 472170 435430 472226
rect 435498 472170 435554 472226
rect 435622 472170 435678 472226
rect 435250 472046 435306 472102
rect 435374 472046 435430 472102
rect 435498 472046 435554 472102
rect 435622 472046 435678 472102
rect 435250 471922 435306 471978
rect 435374 471922 435430 471978
rect 435498 471922 435554 471978
rect 435622 471922 435678 471978
rect 438970 598116 439026 598172
rect 439094 598116 439150 598172
rect 439218 598116 439274 598172
rect 439342 598116 439398 598172
rect 438970 597992 439026 598048
rect 439094 597992 439150 598048
rect 439218 597992 439274 598048
rect 439342 597992 439398 598048
rect 438970 597868 439026 597924
rect 439094 597868 439150 597924
rect 439218 597868 439274 597924
rect 439342 597868 439398 597924
rect 438970 597744 439026 597800
rect 439094 597744 439150 597800
rect 439218 597744 439274 597800
rect 439342 597744 439398 597800
rect 438970 586294 439026 586350
rect 439094 586294 439150 586350
rect 439218 586294 439274 586350
rect 439342 586294 439398 586350
rect 438970 586170 439026 586226
rect 439094 586170 439150 586226
rect 439218 586170 439274 586226
rect 439342 586170 439398 586226
rect 438970 586046 439026 586102
rect 439094 586046 439150 586102
rect 439218 586046 439274 586102
rect 439342 586046 439398 586102
rect 438970 585922 439026 585978
rect 439094 585922 439150 585978
rect 439218 585922 439274 585978
rect 439342 585922 439398 585978
rect 438970 568294 439026 568350
rect 439094 568294 439150 568350
rect 439218 568294 439274 568350
rect 439342 568294 439398 568350
rect 438970 568170 439026 568226
rect 439094 568170 439150 568226
rect 439218 568170 439274 568226
rect 439342 568170 439398 568226
rect 438970 568046 439026 568102
rect 439094 568046 439150 568102
rect 439218 568046 439274 568102
rect 439342 568046 439398 568102
rect 438970 567922 439026 567978
rect 439094 567922 439150 567978
rect 439218 567922 439274 567978
rect 439342 567922 439398 567978
rect 438970 550294 439026 550350
rect 439094 550294 439150 550350
rect 439218 550294 439274 550350
rect 439342 550294 439398 550350
rect 438970 550170 439026 550226
rect 439094 550170 439150 550226
rect 439218 550170 439274 550226
rect 439342 550170 439398 550226
rect 438970 550046 439026 550102
rect 439094 550046 439150 550102
rect 439218 550046 439274 550102
rect 439342 550046 439398 550102
rect 438970 549922 439026 549978
rect 439094 549922 439150 549978
rect 439218 549922 439274 549978
rect 439342 549922 439398 549978
rect 438970 532294 439026 532350
rect 439094 532294 439150 532350
rect 439218 532294 439274 532350
rect 439342 532294 439398 532350
rect 438970 532170 439026 532226
rect 439094 532170 439150 532226
rect 439218 532170 439274 532226
rect 439342 532170 439398 532226
rect 438970 532046 439026 532102
rect 439094 532046 439150 532102
rect 439218 532046 439274 532102
rect 439342 532046 439398 532102
rect 438970 531922 439026 531978
rect 439094 531922 439150 531978
rect 439218 531922 439274 531978
rect 439342 531922 439398 531978
rect 438970 514294 439026 514350
rect 439094 514294 439150 514350
rect 439218 514294 439274 514350
rect 439342 514294 439398 514350
rect 438970 514170 439026 514226
rect 439094 514170 439150 514226
rect 439218 514170 439274 514226
rect 439342 514170 439398 514226
rect 438970 514046 439026 514102
rect 439094 514046 439150 514102
rect 439218 514046 439274 514102
rect 439342 514046 439398 514102
rect 438970 513922 439026 513978
rect 439094 513922 439150 513978
rect 439218 513922 439274 513978
rect 439342 513922 439398 513978
rect 438970 496294 439026 496350
rect 439094 496294 439150 496350
rect 439218 496294 439274 496350
rect 439342 496294 439398 496350
rect 438970 496170 439026 496226
rect 439094 496170 439150 496226
rect 439218 496170 439274 496226
rect 439342 496170 439398 496226
rect 438970 496046 439026 496102
rect 439094 496046 439150 496102
rect 439218 496046 439274 496102
rect 439342 496046 439398 496102
rect 438970 495922 439026 495978
rect 439094 495922 439150 495978
rect 439218 495922 439274 495978
rect 439342 495922 439398 495978
rect 438970 478294 439026 478350
rect 439094 478294 439150 478350
rect 439218 478294 439274 478350
rect 439342 478294 439398 478350
rect 438970 478170 439026 478226
rect 439094 478170 439150 478226
rect 439218 478170 439274 478226
rect 439342 478170 439398 478226
rect 438970 478046 439026 478102
rect 439094 478046 439150 478102
rect 439218 478046 439274 478102
rect 439342 478046 439398 478102
rect 438970 477922 439026 477978
rect 439094 477922 439150 477978
rect 439218 477922 439274 477978
rect 439342 477922 439398 477978
rect 438970 460294 439026 460350
rect 439094 460294 439150 460350
rect 439218 460294 439274 460350
rect 439342 460294 439398 460350
rect 438970 460170 439026 460226
rect 439094 460170 439150 460226
rect 439218 460170 439274 460226
rect 439342 460170 439398 460226
rect 438970 460046 439026 460102
rect 439094 460046 439150 460102
rect 439218 460046 439274 460102
rect 439342 460046 439398 460102
rect 438970 459922 439026 459978
rect 439094 459922 439150 459978
rect 439218 459922 439274 459978
rect 439342 459922 439398 459978
rect 453250 597156 453306 597212
rect 453374 597156 453430 597212
rect 453498 597156 453554 597212
rect 453622 597156 453678 597212
rect 453250 597032 453306 597088
rect 453374 597032 453430 597088
rect 453498 597032 453554 597088
rect 453622 597032 453678 597088
rect 453250 596908 453306 596964
rect 453374 596908 453430 596964
rect 453498 596908 453554 596964
rect 453622 596908 453678 596964
rect 453250 596784 453306 596840
rect 453374 596784 453430 596840
rect 453498 596784 453554 596840
rect 453622 596784 453678 596840
rect 453250 580294 453306 580350
rect 453374 580294 453430 580350
rect 453498 580294 453554 580350
rect 453622 580294 453678 580350
rect 453250 580170 453306 580226
rect 453374 580170 453430 580226
rect 453498 580170 453554 580226
rect 453622 580170 453678 580226
rect 453250 580046 453306 580102
rect 453374 580046 453430 580102
rect 453498 580046 453554 580102
rect 453622 580046 453678 580102
rect 453250 579922 453306 579978
rect 453374 579922 453430 579978
rect 453498 579922 453554 579978
rect 453622 579922 453678 579978
rect 453250 562294 453306 562350
rect 453374 562294 453430 562350
rect 453498 562294 453554 562350
rect 453622 562294 453678 562350
rect 453250 562170 453306 562226
rect 453374 562170 453430 562226
rect 453498 562170 453554 562226
rect 453622 562170 453678 562226
rect 453250 562046 453306 562102
rect 453374 562046 453430 562102
rect 453498 562046 453554 562102
rect 453622 562046 453678 562102
rect 453250 561922 453306 561978
rect 453374 561922 453430 561978
rect 453498 561922 453554 561978
rect 453622 561922 453678 561978
rect 453250 544294 453306 544350
rect 453374 544294 453430 544350
rect 453498 544294 453554 544350
rect 453622 544294 453678 544350
rect 453250 544170 453306 544226
rect 453374 544170 453430 544226
rect 453498 544170 453554 544226
rect 453622 544170 453678 544226
rect 453250 544046 453306 544102
rect 453374 544046 453430 544102
rect 453498 544046 453554 544102
rect 453622 544046 453678 544102
rect 453250 543922 453306 543978
rect 453374 543922 453430 543978
rect 453498 543922 453554 543978
rect 453622 543922 453678 543978
rect 453250 526294 453306 526350
rect 453374 526294 453430 526350
rect 453498 526294 453554 526350
rect 453622 526294 453678 526350
rect 453250 526170 453306 526226
rect 453374 526170 453430 526226
rect 453498 526170 453554 526226
rect 453622 526170 453678 526226
rect 453250 526046 453306 526102
rect 453374 526046 453430 526102
rect 453498 526046 453554 526102
rect 453622 526046 453678 526102
rect 453250 525922 453306 525978
rect 453374 525922 453430 525978
rect 453498 525922 453554 525978
rect 453622 525922 453678 525978
rect 453250 508294 453306 508350
rect 453374 508294 453430 508350
rect 453498 508294 453554 508350
rect 453622 508294 453678 508350
rect 453250 508170 453306 508226
rect 453374 508170 453430 508226
rect 453498 508170 453554 508226
rect 453622 508170 453678 508226
rect 453250 508046 453306 508102
rect 453374 508046 453430 508102
rect 453498 508046 453554 508102
rect 453622 508046 453678 508102
rect 453250 507922 453306 507978
rect 453374 507922 453430 507978
rect 453498 507922 453554 507978
rect 453622 507922 453678 507978
rect 453250 490294 453306 490350
rect 453374 490294 453430 490350
rect 453498 490294 453554 490350
rect 453622 490294 453678 490350
rect 453250 490170 453306 490226
rect 453374 490170 453430 490226
rect 453498 490170 453554 490226
rect 453622 490170 453678 490226
rect 453250 490046 453306 490102
rect 453374 490046 453430 490102
rect 453498 490046 453554 490102
rect 453622 490046 453678 490102
rect 453250 489922 453306 489978
rect 453374 489922 453430 489978
rect 453498 489922 453554 489978
rect 453622 489922 453678 489978
rect 453250 472294 453306 472350
rect 453374 472294 453430 472350
rect 453498 472294 453554 472350
rect 453622 472294 453678 472350
rect 453250 472170 453306 472226
rect 453374 472170 453430 472226
rect 453498 472170 453554 472226
rect 453622 472170 453678 472226
rect 453250 472046 453306 472102
rect 453374 472046 453430 472102
rect 453498 472046 453554 472102
rect 453622 472046 453678 472102
rect 453250 471922 453306 471978
rect 453374 471922 453430 471978
rect 453498 471922 453554 471978
rect 453622 471922 453678 471978
rect 456970 598116 457026 598172
rect 457094 598116 457150 598172
rect 457218 598116 457274 598172
rect 457342 598116 457398 598172
rect 456970 597992 457026 598048
rect 457094 597992 457150 598048
rect 457218 597992 457274 598048
rect 457342 597992 457398 598048
rect 456970 597868 457026 597924
rect 457094 597868 457150 597924
rect 457218 597868 457274 597924
rect 457342 597868 457398 597924
rect 456970 597744 457026 597800
rect 457094 597744 457150 597800
rect 457218 597744 457274 597800
rect 457342 597744 457398 597800
rect 456970 586294 457026 586350
rect 457094 586294 457150 586350
rect 457218 586294 457274 586350
rect 457342 586294 457398 586350
rect 456970 586170 457026 586226
rect 457094 586170 457150 586226
rect 457218 586170 457274 586226
rect 457342 586170 457398 586226
rect 456970 586046 457026 586102
rect 457094 586046 457150 586102
rect 457218 586046 457274 586102
rect 457342 586046 457398 586102
rect 456970 585922 457026 585978
rect 457094 585922 457150 585978
rect 457218 585922 457274 585978
rect 457342 585922 457398 585978
rect 456970 568294 457026 568350
rect 457094 568294 457150 568350
rect 457218 568294 457274 568350
rect 457342 568294 457398 568350
rect 456970 568170 457026 568226
rect 457094 568170 457150 568226
rect 457218 568170 457274 568226
rect 457342 568170 457398 568226
rect 456970 568046 457026 568102
rect 457094 568046 457150 568102
rect 457218 568046 457274 568102
rect 457342 568046 457398 568102
rect 456970 567922 457026 567978
rect 457094 567922 457150 567978
rect 457218 567922 457274 567978
rect 457342 567922 457398 567978
rect 456970 550294 457026 550350
rect 457094 550294 457150 550350
rect 457218 550294 457274 550350
rect 457342 550294 457398 550350
rect 456970 550170 457026 550226
rect 457094 550170 457150 550226
rect 457218 550170 457274 550226
rect 457342 550170 457398 550226
rect 456970 550046 457026 550102
rect 457094 550046 457150 550102
rect 457218 550046 457274 550102
rect 457342 550046 457398 550102
rect 456970 549922 457026 549978
rect 457094 549922 457150 549978
rect 457218 549922 457274 549978
rect 457342 549922 457398 549978
rect 456970 532294 457026 532350
rect 457094 532294 457150 532350
rect 457218 532294 457274 532350
rect 457342 532294 457398 532350
rect 456970 532170 457026 532226
rect 457094 532170 457150 532226
rect 457218 532170 457274 532226
rect 457342 532170 457398 532226
rect 456970 532046 457026 532102
rect 457094 532046 457150 532102
rect 457218 532046 457274 532102
rect 457342 532046 457398 532102
rect 456970 531922 457026 531978
rect 457094 531922 457150 531978
rect 457218 531922 457274 531978
rect 457342 531922 457398 531978
rect 456970 514294 457026 514350
rect 457094 514294 457150 514350
rect 457218 514294 457274 514350
rect 457342 514294 457398 514350
rect 456970 514170 457026 514226
rect 457094 514170 457150 514226
rect 457218 514170 457274 514226
rect 457342 514170 457398 514226
rect 456970 514046 457026 514102
rect 457094 514046 457150 514102
rect 457218 514046 457274 514102
rect 457342 514046 457398 514102
rect 456970 513922 457026 513978
rect 457094 513922 457150 513978
rect 457218 513922 457274 513978
rect 457342 513922 457398 513978
rect 456970 496294 457026 496350
rect 457094 496294 457150 496350
rect 457218 496294 457274 496350
rect 457342 496294 457398 496350
rect 456970 496170 457026 496226
rect 457094 496170 457150 496226
rect 457218 496170 457274 496226
rect 457342 496170 457398 496226
rect 456970 496046 457026 496102
rect 457094 496046 457150 496102
rect 457218 496046 457274 496102
rect 457342 496046 457398 496102
rect 456970 495922 457026 495978
rect 457094 495922 457150 495978
rect 457218 495922 457274 495978
rect 457342 495922 457398 495978
rect 456970 478294 457026 478350
rect 457094 478294 457150 478350
rect 457218 478294 457274 478350
rect 457342 478294 457398 478350
rect 456970 478170 457026 478226
rect 457094 478170 457150 478226
rect 457218 478170 457274 478226
rect 457342 478170 457398 478226
rect 456970 478046 457026 478102
rect 457094 478046 457150 478102
rect 457218 478046 457274 478102
rect 457342 478046 457398 478102
rect 456970 477922 457026 477978
rect 457094 477922 457150 477978
rect 457218 477922 457274 477978
rect 457342 477922 457398 477978
rect 456970 460294 457026 460350
rect 457094 460294 457150 460350
rect 457218 460294 457274 460350
rect 457342 460294 457398 460350
rect 456970 460170 457026 460226
rect 457094 460170 457150 460226
rect 457218 460170 457274 460226
rect 457342 460170 457398 460226
rect 456970 460046 457026 460102
rect 457094 460046 457150 460102
rect 457218 460046 457274 460102
rect 457342 460046 457398 460102
rect 456970 459922 457026 459978
rect 457094 459922 457150 459978
rect 457218 459922 457274 459978
rect 457342 459922 457398 459978
rect 471250 597156 471306 597212
rect 471374 597156 471430 597212
rect 471498 597156 471554 597212
rect 471622 597156 471678 597212
rect 471250 597032 471306 597088
rect 471374 597032 471430 597088
rect 471498 597032 471554 597088
rect 471622 597032 471678 597088
rect 471250 596908 471306 596964
rect 471374 596908 471430 596964
rect 471498 596908 471554 596964
rect 471622 596908 471678 596964
rect 471250 596784 471306 596840
rect 471374 596784 471430 596840
rect 471498 596784 471554 596840
rect 471622 596784 471678 596840
rect 471250 580294 471306 580350
rect 471374 580294 471430 580350
rect 471498 580294 471554 580350
rect 471622 580294 471678 580350
rect 471250 580170 471306 580226
rect 471374 580170 471430 580226
rect 471498 580170 471554 580226
rect 471622 580170 471678 580226
rect 471250 580046 471306 580102
rect 471374 580046 471430 580102
rect 471498 580046 471554 580102
rect 471622 580046 471678 580102
rect 471250 579922 471306 579978
rect 471374 579922 471430 579978
rect 471498 579922 471554 579978
rect 471622 579922 471678 579978
rect 471250 562294 471306 562350
rect 471374 562294 471430 562350
rect 471498 562294 471554 562350
rect 471622 562294 471678 562350
rect 471250 562170 471306 562226
rect 471374 562170 471430 562226
rect 471498 562170 471554 562226
rect 471622 562170 471678 562226
rect 471250 562046 471306 562102
rect 471374 562046 471430 562102
rect 471498 562046 471554 562102
rect 471622 562046 471678 562102
rect 471250 561922 471306 561978
rect 471374 561922 471430 561978
rect 471498 561922 471554 561978
rect 471622 561922 471678 561978
rect 471250 544294 471306 544350
rect 471374 544294 471430 544350
rect 471498 544294 471554 544350
rect 471622 544294 471678 544350
rect 471250 544170 471306 544226
rect 471374 544170 471430 544226
rect 471498 544170 471554 544226
rect 471622 544170 471678 544226
rect 471250 544046 471306 544102
rect 471374 544046 471430 544102
rect 471498 544046 471554 544102
rect 471622 544046 471678 544102
rect 471250 543922 471306 543978
rect 471374 543922 471430 543978
rect 471498 543922 471554 543978
rect 471622 543922 471678 543978
rect 471250 526294 471306 526350
rect 471374 526294 471430 526350
rect 471498 526294 471554 526350
rect 471622 526294 471678 526350
rect 471250 526170 471306 526226
rect 471374 526170 471430 526226
rect 471498 526170 471554 526226
rect 471622 526170 471678 526226
rect 471250 526046 471306 526102
rect 471374 526046 471430 526102
rect 471498 526046 471554 526102
rect 471622 526046 471678 526102
rect 471250 525922 471306 525978
rect 471374 525922 471430 525978
rect 471498 525922 471554 525978
rect 471622 525922 471678 525978
rect 471250 508294 471306 508350
rect 471374 508294 471430 508350
rect 471498 508294 471554 508350
rect 471622 508294 471678 508350
rect 471250 508170 471306 508226
rect 471374 508170 471430 508226
rect 471498 508170 471554 508226
rect 471622 508170 471678 508226
rect 471250 508046 471306 508102
rect 471374 508046 471430 508102
rect 471498 508046 471554 508102
rect 471622 508046 471678 508102
rect 471250 507922 471306 507978
rect 471374 507922 471430 507978
rect 471498 507922 471554 507978
rect 471622 507922 471678 507978
rect 471250 490294 471306 490350
rect 471374 490294 471430 490350
rect 471498 490294 471554 490350
rect 471622 490294 471678 490350
rect 471250 490170 471306 490226
rect 471374 490170 471430 490226
rect 471498 490170 471554 490226
rect 471622 490170 471678 490226
rect 471250 490046 471306 490102
rect 471374 490046 471430 490102
rect 471498 490046 471554 490102
rect 471622 490046 471678 490102
rect 471250 489922 471306 489978
rect 471374 489922 471430 489978
rect 471498 489922 471554 489978
rect 471622 489922 471678 489978
rect 471250 472294 471306 472350
rect 471374 472294 471430 472350
rect 471498 472294 471554 472350
rect 471622 472294 471678 472350
rect 471250 472170 471306 472226
rect 471374 472170 471430 472226
rect 471498 472170 471554 472226
rect 471622 472170 471678 472226
rect 471250 472046 471306 472102
rect 471374 472046 471430 472102
rect 471498 472046 471554 472102
rect 471622 472046 471678 472102
rect 471250 471922 471306 471978
rect 471374 471922 471430 471978
rect 471498 471922 471554 471978
rect 471622 471922 471678 471978
rect 474970 598116 475026 598172
rect 475094 598116 475150 598172
rect 475218 598116 475274 598172
rect 475342 598116 475398 598172
rect 474970 597992 475026 598048
rect 475094 597992 475150 598048
rect 475218 597992 475274 598048
rect 475342 597992 475398 598048
rect 474970 597868 475026 597924
rect 475094 597868 475150 597924
rect 475218 597868 475274 597924
rect 475342 597868 475398 597924
rect 474970 597744 475026 597800
rect 475094 597744 475150 597800
rect 475218 597744 475274 597800
rect 475342 597744 475398 597800
rect 474970 586294 475026 586350
rect 475094 586294 475150 586350
rect 475218 586294 475274 586350
rect 475342 586294 475398 586350
rect 474970 586170 475026 586226
rect 475094 586170 475150 586226
rect 475218 586170 475274 586226
rect 475342 586170 475398 586226
rect 474970 586046 475026 586102
rect 475094 586046 475150 586102
rect 475218 586046 475274 586102
rect 475342 586046 475398 586102
rect 474970 585922 475026 585978
rect 475094 585922 475150 585978
rect 475218 585922 475274 585978
rect 475342 585922 475398 585978
rect 474970 568294 475026 568350
rect 475094 568294 475150 568350
rect 475218 568294 475274 568350
rect 475342 568294 475398 568350
rect 474970 568170 475026 568226
rect 475094 568170 475150 568226
rect 475218 568170 475274 568226
rect 475342 568170 475398 568226
rect 474970 568046 475026 568102
rect 475094 568046 475150 568102
rect 475218 568046 475274 568102
rect 475342 568046 475398 568102
rect 474970 567922 475026 567978
rect 475094 567922 475150 567978
rect 475218 567922 475274 567978
rect 475342 567922 475398 567978
rect 474970 550294 475026 550350
rect 475094 550294 475150 550350
rect 475218 550294 475274 550350
rect 475342 550294 475398 550350
rect 474970 550170 475026 550226
rect 475094 550170 475150 550226
rect 475218 550170 475274 550226
rect 475342 550170 475398 550226
rect 474970 550046 475026 550102
rect 475094 550046 475150 550102
rect 475218 550046 475274 550102
rect 475342 550046 475398 550102
rect 474970 549922 475026 549978
rect 475094 549922 475150 549978
rect 475218 549922 475274 549978
rect 475342 549922 475398 549978
rect 474970 532294 475026 532350
rect 475094 532294 475150 532350
rect 475218 532294 475274 532350
rect 475342 532294 475398 532350
rect 474970 532170 475026 532226
rect 475094 532170 475150 532226
rect 475218 532170 475274 532226
rect 475342 532170 475398 532226
rect 474970 532046 475026 532102
rect 475094 532046 475150 532102
rect 475218 532046 475274 532102
rect 475342 532046 475398 532102
rect 474970 531922 475026 531978
rect 475094 531922 475150 531978
rect 475218 531922 475274 531978
rect 475342 531922 475398 531978
rect 474970 514294 475026 514350
rect 475094 514294 475150 514350
rect 475218 514294 475274 514350
rect 475342 514294 475398 514350
rect 474970 514170 475026 514226
rect 475094 514170 475150 514226
rect 475218 514170 475274 514226
rect 475342 514170 475398 514226
rect 474970 514046 475026 514102
rect 475094 514046 475150 514102
rect 475218 514046 475274 514102
rect 475342 514046 475398 514102
rect 474970 513922 475026 513978
rect 475094 513922 475150 513978
rect 475218 513922 475274 513978
rect 475342 513922 475398 513978
rect 474970 496294 475026 496350
rect 475094 496294 475150 496350
rect 475218 496294 475274 496350
rect 475342 496294 475398 496350
rect 474970 496170 475026 496226
rect 475094 496170 475150 496226
rect 475218 496170 475274 496226
rect 475342 496170 475398 496226
rect 474970 496046 475026 496102
rect 475094 496046 475150 496102
rect 475218 496046 475274 496102
rect 475342 496046 475398 496102
rect 474970 495922 475026 495978
rect 475094 495922 475150 495978
rect 475218 495922 475274 495978
rect 475342 495922 475398 495978
rect 474970 478294 475026 478350
rect 475094 478294 475150 478350
rect 475218 478294 475274 478350
rect 475342 478294 475398 478350
rect 474970 478170 475026 478226
rect 475094 478170 475150 478226
rect 475218 478170 475274 478226
rect 475342 478170 475398 478226
rect 474970 478046 475026 478102
rect 475094 478046 475150 478102
rect 475218 478046 475274 478102
rect 475342 478046 475398 478102
rect 474970 477922 475026 477978
rect 475094 477922 475150 477978
rect 475218 477922 475274 477978
rect 475342 477922 475398 477978
rect 474970 460294 475026 460350
rect 475094 460294 475150 460350
rect 475218 460294 475274 460350
rect 475342 460294 475398 460350
rect 474970 460170 475026 460226
rect 475094 460170 475150 460226
rect 475218 460170 475274 460226
rect 475342 460170 475398 460226
rect 474970 460046 475026 460102
rect 475094 460046 475150 460102
rect 475218 460046 475274 460102
rect 475342 460046 475398 460102
rect 474970 459922 475026 459978
rect 475094 459922 475150 459978
rect 475218 459922 475274 459978
rect 475342 459922 475398 459978
rect 489250 597156 489306 597212
rect 489374 597156 489430 597212
rect 489498 597156 489554 597212
rect 489622 597156 489678 597212
rect 489250 597032 489306 597088
rect 489374 597032 489430 597088
rect 489498 597032 489554 597088
rect 489622 597032 489678 597088
rect 489250 596908 489306 596964
rect 489374 596908 489430 596964
rect 489498 596908 489554 596964
rect 489622 596908 489678 596964
rect 489250 596784 489306 596840
rect 489374 596784 489430 596840
rect 489498 596784 489554 596840
rect 489622 596784 489678 596840
rect 489250 580294 489306 580350
rect 489374 580294 489430 580350
rect 489498 580294 489554 580350
rect 489622 580294 489678 580350
rect 489250 580170 489306 580226
rect 489374 580170 489430 580226
rect 489498 580170 489554 580226
rect 489622 580170 489678 580226
rect 489250 580046 489306 580102
rect 489374 580046 489430 580102
rect 489498 580046 489554 580102
rect 489622 580046 489678 580102
rect 489250 579922 489306 579978
rect 489374 579922 489430 579978
rect 489498 579922 489554 579978
rect 489622 579922 489678 579978
rect 489250 562294 489306 562350
rect 489374 562294 489430 562350
rect 489498 562294 489554 562350
rect 489622 562294 489678 562350
rect 489250 562170 489306 562226
rect 489374 562170 489430 562226
rect 489498 562170 489554 562226
rect 489622 562170 489678 562226
rect 489250 562046 489306 562102
rect 489374 562046 489430 562102
rect 489498 562046 489554 562102
rect 489622 562046 489678 562102
rect 489250 561922 489306 561978
rect 489374 561922 489430 561978
rect 489498 561922 489554 561978
rect 489622 561922 489678 561978
rect 489250 544294 489306 544350
rect 489374 544294 489430 544350
rect 489498 544294 489554 544350
rect 489622 544294 489678 544350
rect 489250 544170 489306 544226
rect 489374 544170 489430 544226
rect 489498 544170 489554 544226
rect 489622 544170 489678 544226
rect 489250 544046 489306 544102
rect 489374 544046 489430 544102
rect 489498 544046 489554 544102
rect 489622 544046 489678 544102
rect 489250 543922 489306 543978
rect 489374 543922 489430 543978
rect 489498 543922 489554 543978
rect 489622 543922 489678 543978
rect 489250 526294 489306 526350
rect 489374 526294 489430 526350
rect 489498 526294 489554 526350
rect 489622 526294 489678 526350
rect 489250 526170 489306 526226
rect 489374 526170 489430 526226
rect 489498 526170 489554 526226
rect 489622 526170 489678 526226
rect 489250 526046 489306 526102
rect 489374 526046 489430 526102
rect 489498 526046 489554 526102
rect 489622 526046 489678 526102
rect 489250 525922 489306 525978
rect 489374 525922 489430 525978
rect 489498 525922 489554 525978
rect 489622 525922 489678 525978
rect 489250 508294 489306 508350
rect 489374 508294 489430 508350
rect 489498 508294 489554 508350
rect 489622 508294 489678 508350
rect 489250 508170 489306 508226
rect 489374 508170 489430 508226
rect 489498 508170 489554 508226
rect 489622 508170 489678 508226
rect 489250 508046 489306 508102
rect 489374 508046 489430 508102
rect 489498 508046 489554 508102
rect 489622 508046 489678 508102
rect 489250 507922 489306 507978
rect 489374 507922 489430 507978
rect 489498 507922 489554 507978
rect 489622 507922 489678 507978
rect 489250 490294 489306 490350
rect 489374 490294 489430 490350
rect 489498 490294 489554 490350
rect 489622 490294 489678 490350
rect 489250 490170 489306 490226
rect 489374 490170 489430 490226
rect 489498 490170 489554 490226
rect 489622 490170 489678 490226
rect 489250 490046 489306 490102
rect 489374 490046 489430 490102
rect 489498 490046 489554 490102
rect 489622 490046 489678 490102
rect 489250 489922 489306 489978
rect 489374 489922 489430 489978
rect 489498 489922 489554 489978
rect 489622 489922 489678 489978
rect 489250 472294 489306 472350
rect 489374 472294 489430 472350
rect 489498 472294 489554 472350
rect 489622 472294 489678 472350
rect 489250 472170 489306 472226
rect 489374 472170 489430 472226
rect 489498 472170 489554 472226
rect 489622 472170 489678 472226
rect 489250 472046 489306 472102
rect 489374 472046 489430 472102
rect 489498 472046 489554 472102
rect 489622 472046 489678 472102
rect 489250 471922 489306 471978
rect 489374 471922 489430 471978
rect 489498 471922 489554 471978
rect 489622 471922 489678 471978
rect 492970 598116 493026 598172
rect 493094 598116 493150 598172
rect 493218 598116 493274 598172
rect 493342 598116 493398 598172
rect 492970 597992 493026 598048
rect 493094 597992 493150 598048
rect 493218 597992 493274 598048
rect 493342 597992 493398 598048
rect 492970 597868 493026 597924
rect 493094 597868 493150 597924
rect 493218 597868 493274 597924
rect 493342 597868 493398 597924
rect 492970 597744 493026 597800
rect 493094 597744 493150 597800
rect 493218 597744 493274 597800
rect 493342 597744 493398 597800
rect 492970 586294 493026 586350
rect 493094 586294 493150 586350
rect 493218 586294 493274 586350
rect 493342 586294 493398 586350
rect 492970 586170 493026 586226
rect 493094 586170 493150 586226
rect 493218 586170 493274 586226
rect 493342 586170 493398 586226
rect 492970 586046 493026 586102
rect 493094 586046 493150 586102
rect 493218 586046 493274 586102
rect 493342 586046 493398 586102
rect 492970 585922 493026 585978
rect 493094 585922 493150 585978
rect 493218 585922 493274 585978
rect 493342 585922 493398 585978
rect 492970 568294 493026 568350
rect 493094 568294 493150 568350
rect 493218 568294 493274 568350
rect 493342 568294 493398 568350
rect 492970 568170 493026 568226
rect 493094 568170 493150 568226
rect 493218 568170 493274 568226
rect 493342 568170 493398 568226
rect 492970 568046 493026 568102
rect 493094 568046 493150 568102
rect 493218 568046 493274 568102
rect 493342 568046 493398 568102
rect 492970 567922 493026 567978
rect 493094 567922 493150 567978
rect 493218 567922 493274 567978
rect 493342 567922 493398 567978
rect 492970 550294 493026 550350
rect 493094 550294 493150 550350
rect 493218 550294 493274 550350
rect 493342 550294 493398 550350
rect 492970 550170 493026 550226
rect 493094 550170 493150 550226
rect 493218 550170 493274 550226
rect 493342 550170 493398 550226
rect 492970 550046 493026 550102
rect 493094 550046 493150 550102
rect 493218 550046 493274 550102
rect 493342 550046 493398 550102
rect 492970 549922 493026 549978
rect 493094 549922 493150 549978
rect 493218 549922 493274 549978
rect 493342 549922 493398 549978
rect 492970 532294 493026 532350
rect 493094 532294 493150 532350
rect 493218 532294 493274 532350
rect 493342 532294 493398 532350
rect 492970 532170 493026 532226
rect 493094 532170 493150 532226
rect 493218 532170 493274 532226
rect 493342 532170 493398 532226
rect 492970 532046 493026 532102
rect 493094 532046 493150 532102
rect 493218 532046 493274 532102
rect 493342 532046 493398 532102
rect 492970 531922 493026 531978
rect 493094 531922 493150 531978
rect 493218 531922 493274 531978
rect 493342 531922 493398 531978
rect 492970 514294 493026 514350
rect 493094 514294 493150 514350
rect 493218 514294 493274 514350
rect 493342 514294 493398 514350
rect 492970 514170 493026 514226
rect 493094 514170 493150 514226
rect 493218 514170 493274 514226
rect 493342 514170 493398 514226
rect 492970 514046 493026 514102
rect 493094 514046 493150 514102
rect 493218 514046 493274 514102
rect 493342 514046 493398 514102
rect 492970 513922 493026 513978
rect 493094 513922 493150 513978
rect 493218 513922 493274 513978
rect 493342 513922 493398 513978
rect 492970 496294 493026 496350
rect 493094 496294 493150 496350
rect 493218 496294 493274 496350
rect 493342 496294 493398 496350
rect 492970 496170 493026 496226
rect 493094 496170 493150 496226
rect 493218 496170 493274 496226
rect 493342 496170 493398 496226
rect 492970 496046 493026 496102
rect 493094 496046 493150 496102
rect 493218 496046 493274 496102
rect 493342 496046 493398 496102
rect 492970 495922 493026 495978
rect 493094 495922 493150 495978
rect 493218 495922 493274 495978
rect 493342 495922 493398 495978
rect 492970 478294 493026 478350
rect 493094 478294 493150 478350
rect 493218 478294 493274 478350
rect 493342 478294 493398 478350
rect 492970 478170 493026 478226
rect 493094 478170 493150 478226
rect 493218 478170 493274 478226
rect 493342 478170 493398 478226
rect 492970 478046 493026 478102
rect 493094 478046 493150 478102
rect 493218 478046 493274 478102
rect 493342 478046 493398 478102
rect 492970 477922 493026 477978
rect 493094 477922 493150 477978
rect 493218 477922 493274 477978
rect 493342 477922 493398 477978
rect 492970 460294 493026 460350
rect 493094 460294 493150 460350
rect 493218 460294 493274 460350
rect 493342 460294 493398 460350
rect 492970 460170 493026 460226
rect 493094 460170 493150 460226
rect 493218 460170 493274 460226
rect 493342 460170 493398 460226
rect 492970 460046 493026 460102
rect 493094 460046 493150 460102
rect 493218 460046 493274 460102
rect 493342 460046 493398 460102
rect 492970 459922 493026 459978
rect 493094 459922 493150 459978
rect 493218 459922 493274 459978
rect 493342 459922 493398 459978
rect 507250 597156 507306 597212
rect 507374 597156 507430 597212
rect 507498 597156 507554 597212
rect 507622 597156 507678 597212
rect 507250 597032 507306 597088
rect 507374 597032 507430 597088
rect 507498 597032 507554 597088
rect 507622 597032 507678 597088
rect 507250 596908 507306 596964
rect 507374 596908 507430 596964
rect 507498 596908 507554 596964
rect 507622 596908 507678 596964
rect 507250 596784 507306 596840
rect 507374 596784 507430 596840
rect 507498 596784 507554 596840
rect 507622 596784 507678 596840
rect 507250 580294 507306 580350
rect 507374 580294 507430 580350
rect 507498 580294 507554 580350
rect 507622 580294 507678 580350
rect 507250 580170 507306 580226
rect 507374 580170 507430 580226
rect 507498 580170 507554 580226
rect 507622 580170 507678 580226
rect 507250 580046 507306 580102
rect 507374 580046 507430 580102
rect 507498 580046 507554 580102
rect 507622 580046 507678 580102
rect 507250 579922 507306 579978
rect 507374 579922 507430 579978
rect 507498 579922 507554 579978
rect 507622 579922 507678 579978
rect 507250 562294 507306 562350
rect 507374 562294 507430 562350
rect 507498 562294 507554 562350
rect 507622 562294 507678 562350
rect 507250 562170 507306 562226
rect 507374 562170 507430 562226
rect 507498 562170 507554 562226
rect 507622 562170 507678 562226
rect 507250 562046 507306 562102
rect 507374 562046 507430 562102
rect 507498 562046 507554 562102
rect 507622 562046 507678 562102
rect 507250 561922 507306 561978
rect 507374 561922 507430 561978
rect 507498 561922 507554 561978
rect 507622 561922 507678 561978
rect 507250 544294 507306 544350
rect 507374 544294 507430 544350
rect 507498 544294 507554 544350
rect 507622 544294 507678 544350
rect 507250 544170 507306 544226
rect 507374 544170 507430 544226
rect 507498 544170 507554 544226
rect 507622 544170 507678 544226
rect 507250 544046 507306 544102
rect 507374 544046 507430 544102
rect 507498 544046 507554 544102
rect 507622 544046 507678 544102
rect 507250 543922 507306 543978
rect 507374 543922 507430 543978
rect 507498 543922 507554 543978
rect 507622 543922 507678 543978
rect 507250 526294 507306 526350
rect 507374 526294 507430 526350
rect 507498 526294 507554 526350
rect 507622 526294 507678 526350
rect 507250 526170 507306 526226
rect 507374 526170 507430 526226
rect 507498 526170 507554 526226
rect 507622 526170 507678 526226
rect 507250 526046 507306 526102
rect 507374 526046 507430 526102
rect 507498 526046 507554 526102
rect 507622 526046 507678 526102
rect 507250 525922 507306 525978
rect 507374 525922 507430 525978
rect 507498 525922 507554 525978
rect 507622 525922 507678 525978
rect 507250 508294 507306 508350
rect 507374 508294 507430 508350
rect 507498 508294 507554 508350
rect 507622 508294 507678 508350
rect 507250 508170 507306 508226
rect 507374 508170 507430 508226
rect 507498 508170 507554 508226
rect 507622 508170 507678 508226
rect 507250 508046 507306 508102
rect 507374 508046 507430 508102
rect 507498 508046 507554 508102
rect 507622 508046 507678 508102
rect 507250 507922 507306 507978
rect 507374 507922 507430 507978
rect 507498 507922 507554 507978
rect 507622 507922 507678 507978
rect 507250 490294 507306 490350
rect 507374 490294 507430 490350
rect 507498 490294 507554 490350
rect 507622 490294 507678 490350
rect 507250 490170 507306 490226
rect 507374 490170 507430 490226
rect 507498 490170 507554 490226
rect 507622 490170 507678 490226
rect 507250 490046 507306 490102
rect 507374 490046 507430 490102
rect 507498 490046 507554 490102
rect 507622 490046 507678 490102
rect 507250 489922 507306 489978
rect 507374 489922 507430 489978
rect 507498 489922 507554 489978
rect 507622 489922 507678 489978
rect 507250 472294 507306 472350
rect 507374 472294 507430 472350
rect 507498 472294 507554 472350
rect 507622 472294 507678 472350
rect 507250 472170 507306 472226
rect 507374 472170 507430 472226
rect 507498 472170 507554 472226
rect 507622 472170 507678 472226
rect 507250 472046 507306 472102
rect 507374 472046 507430 472102
rect 507498 472046 507554 472102
rect 507622 472046 507678 472102
rect 507250 471922 507306 471978
rect 507374 471922 507430 471978
rect 507498 471922 507554 471978
rect 507622 471922 507678 471978
rect 510970 598116 511026 598172
rect 511094 598116 511150 598172
rect 511218 598116 511274 598172
rect 511342 598116 511398 598172
rect 510970 597992 511026 598048
rect 511094 597992 511150 598048
rect 511218 597992 511274 598048
rect 511342 597992 511398 598048
rect 510970 597868 511026 597924
rect 511094 597868 511150 597924
rect 511218 597868 511274 597924
rect 511342 597868 511398 597924
rect 510970 597744 511026 597800
rect 511094 597744 511150 597800
rect 511218 597744 511274 597800
rect 511342 597744 511398 597800
rect 510970 586294 511026 586350
rect 511094 586294 511150 586350
rect 511218 586294 511274 586350
rect 511342 586294 511398 586350
rect 510970 586170 511026 586226
rect 511094 586170 511150 586226
rect 511218 586170 511274 586226
rect 511342 586170 511398 586226
rect 510970 586046 511026 586102
rect 511094 586046 511150 586102
rect 511218 586046 511274 586102
rect 511342 586046 511398 586102
rect 510970 585922 511026 585978
rect 511094 585922 511150 585978
rect 511218 585922 511274 585978
rect 511342 585922 511398 585978
rect 510970 568294 511026 568350
rect 511094 568294 511150 568350
rect 511218 568294 511274 568350
rect 511342 568294 511398 568350
rect 510970 568170 511026 568226
rect 511094 568170 511150 568226
rect 511218 568170 511274 568226
rect 511342 568170 511398 568226
rect 510970 568046 511026 568102
rect 511094 568046 511150 568102
rect 511218 568046 511274 568102
rect 511342 568046 511398 568102
rect 510970 567922 511026 567978
rect 511094 567922 511150 567978
rect 511218 567922 511274 567978
rect 511342 567922 511398 567978
rect 510970 550294 511026 550350
rect 511094 550294 511150 550350
rect 511218 550294 511274 550350
rect 511342 550294 511398 550350
rect 510970 550170 511026 550226
rect 511094 550170 511150 550226
rect 511218 550170 511274 550226
rect 511342 550170 511398 550226
rect 510970 550046 511026 550102
rect 511094 550046 511150 550102
rect 511218 550046 511274 550102
rect 511342 550046 511398 550102
rect 510970 549922 511026 549978
rect 511094 549922 511150 549978
rect 511218 549922 511274 549978
rect 511342 549922 511398 549978
rect 510970 532294 511026 532350
rect 511094 532294 511150 532350
rect 511218 532294 511274 532350
rect 511342 532294 511398 532350
rect 510970 532170 511026 532226
rect 511094 532170 511150 532226
rect 511218 532170 511274 532226
rect 511342 532170 511398 532226
rect 510970 532046 511026 532102
rect 511094 532046 511150 532102
rect 511218 532046 511274 532102
rect 511342 532046 511398 532102
rect 510970 531922 511026 531978
rect 511094 531922 511150 531978
rect 511218 531922 511274 531978
rect 511342 531922 511398 531978
rect 510970 514294 511026 514350
rect 511094 514294 511150 514350
rect 511218 514294 511274 514350
rect 511342 514294 511398 514350
rect 510970 514170 511026 514226
rect 511094 514170 511150 514226
rect 511218 514170 511274 514226
rect 511342 514170 511398 514226
rect 510970 514046 511026 514102
rect 511094 514046 511150 514102
rect 511218 514046 511274 514102
rect 511342 514046 511398 514102
rect 510970 513922 511026 513978
rect 511094 513922 511150 513978
rect 511218 513922 511274 513978
rect 511342 513922 511398 513978
rect 510970 496294 511026 496350
rect 511094 496294 511150 496350
rect 511218 496294 511274 496350
rect 511342 496294 511398 496350
rect 510970 496170 511026 496226
rect 511094 496170 511150 496226
rect 511218 496170 511274 496226
rect 511342 496170 511398 496226
rect 510970 496046 511026 496102
rect 511094 496046 511150 496102
rect 511218 496046 511274 496102
rect 511342 496046 511398 496102
rect 510970 495922 511026 495978
rect 511094 495922 511150 495978
rect 511218 495922 511274 495978
rect 511342 495922 511398 495978
rect 510970 478294 511026 478350
rect 511094 478294 511150 478350
rect 511218 478294 511274 478350
rect 511342 478294 511398 478350
rect 510970 478170 511026 478226
rect 511094 478170 511150 478226
rect 511218 478170 511274 478226
rect 511342 478170 511398 478226
rect 510970 478046 511026 478102
rect 511094 478046 511150 478102
rect 511218 478046 511274 478102
rect 511342 478046 511398 478102
rect 510970 477922 511026 477978
rect 511094 477922 511150 477978
rect 511218 477922 511274 477978
rect 511342 477922 511398 477978
rect 510970 460294 511026 460350
rect 511094 460294 511150 460350
rect 511218 460294 511274 460350
rect 511342 460294 511398 460350
rect 510970 460170 511026 460226
rect 511094 460170 511150 460226
rect 511218 460170 511274 460226
rect 511342 460170 511398 460226
rect 510970 460046 511026 460102
rect 511094 460046 511150 460102
rect 511218 460046 511274 460102
rect 511342 460046 511398 460102
rect 510970 459922 511026 459978
rect 511094 459922 511150 459978
rect 511218 459922 511274 459978
rect 511342 459922 511398 459978
rect 525250 597156 525306 597212
rect 525374 597156 525430 597212
rect 525498 597156 525554 597212
rect 525622 597156 525678 597212
rect 525250 597032 525306 597088
rect 525374 597032 525430 597088
rect 525498 597032 525554 597088
rect 525622 597032 525678 597088
rect 525250 596908 525306 596964
rect 525374 596908 525430 596964
rect 525498 596908 525554 596964
rect 525622 596908 525678 596964
rect 525250 596784 525306 596840
rect 525374 596784 525430 596840
rect 525498 596784 525554 596840
rect 525622 596784 525678 596840
rect 525250 580294 525306 580350
rect 525374 580294 525430 580350
rect 525498 580294 525554 580350
rect 525622 580294 525678 580350
rect 525250 580170 525306 580226
rect 525374 580170 525430 580226
rect 525498 580170 525554 580226
rect 525622 580170 525678 580226
rect 525250 580046 525306 580102
rect 525374 580046 525430 580102
rect 525498 580046 525554 580102
rect 525622 580046 525678 580102
rect 525250 579922 525306 579978
rect 525374 579922 525430 579978
rect 525498 579922 525554 579978
rect 525622 579922 525678 579978
rect 525250 562294 525306 562350
rect 525374 562294 525430 562350
rect 525498 562294 525554 562350
rect 525622 562294 525678 562350
rect 525250 562170 525306 562226
rect 525374 562170 525430 562226
rect 525498 562170 525554 562226
rect 525622 562170 525678 562226
rect 525250 562046 525306 562102
rect 525374 562046 525430 562102
rect 525498 562046 525554 562102
rect 525622 562046 525678 562102
rect 525250 561922 525306 561978
rect 525374 561922 525430 561978
rect 525498 561922 525554 561978
rect 525622 561922 525678 561978
rect 525250 544294 525306 544350
rect 525374 544294 525430 544350
rect 525498 544294 525554 544350
rect 525622 544294 525678 544350
rect 525250 544170 525306 544226
rect 525374 544170 525430 544226
rect 525498 544170 525554 544226
rect 525622 544170 525678 544226
rect 525250 544046 525306 544102
rect 525374 544046 525430 544102
rect 525498 544046 525554 544102
rect 525622 544046 525678 544102
rect 525250 543922 525306 543978
rect 525374 543922 525430 543978
rect 525498 543922 525554 543978
rect 525622 543922 525678 543978
rect 525250 526294 525306 526350
rect 525374 526294 525430 526350
rect 525498 526294 525554 526350
rect 525622 526294 525678 526350
rect 525250 526170 525306 526226
rect 525374 526170 525430 526226
rect 525498 526170 525554 526226
rect 525622 526170 525678 526226
rect 525250 526046 525306 526102
rect 525374 526046 525430 526102
rect 525498 526046 525554 526102
rect 525622 526046 525678 526102
rect 525250 525922 525306 525978
rect 525374 525922 525430 525978
rect 525498 525922 525554 525978
rect 525622 525922 525678 525978
rect 525250 508294 525306 508350
rect 525374 508294 525430 508350
rect 525498 508294 525554 508350
rect 525622 508294 525678 508350
rect 525250 508170 525306 508226
rect 525374 508170 525430 508226
rect 525498 508170 525554 508226
rect 525622 508170 525678 508226
rect 525250 508046 525306 508102
rect 525374 508046 525430 508102
rect 525498 508046 525554 508102
rect 525622 508046 525678 508102
rect 525250 507922 525306 507978
rect 525374 507922 525430 507978
rect 525498 507922 525554 507978
rect 525622 507922 525678 507978
rect 525250 490294 525306 490350
rect 525374 490294 525430 490350
rect 525498 490294 525554 490350
rect 525622 490294 525678 490350
rect 525250 490170 525306 490226
rect 525374 490170 525430 490226
rect 525498 490170 525554 490226
rect 525622 490170 525678 490226
rect 525250 490046 525306 490102
rect 525374 490046 525430 490102
rect 525498 490046 525554 490102
rect 525622 490046 525678 490102
rect 525250 489922 525306 489978
rect 525374 489922 525430 489978
rect 525498 489922 525554 489978
rect 525622 489922 525678 489978
rect 525250 472294 525306 472350
rect 525374 472294 525430 472350
rect 525498 472294 525554 472350
rect 525622 472294 525678 472350
rect 525250 472170 525306 472226
rect 525374 472170 525430 472226
rect 525498 472170 525554 472226
rect 525622 472170 525678 472226
rect 525250 472046 525306 472102
rect 525374 472046 525430 472102
rect 525498 472046 525554 472102
rect 525622 472046 525678 472102
rect 525250 471922 525306 471978
rect 525374 471922 525430 471978
rect 525498 471922 525554 471978
rect 525622 471922 525678 471978
rect 528970 598116 529026 598172
rect 529094 598116 529150 598172
rect 529218 598116 529274 598172
rect 529342 598116 529398 598172
rect 528970 597992 529026 598048
rect 529094 597992 529150 598048
rect 529218 597992 529274 598048
rect 529342 597992 529398 598048
rect 528970 597868 529026 597924
rect 529094 597868 529150 597924
rect 529218 597868 529274 597924
rect 529342 597868 529398 597924
rect 528970 597744 529026 597800
rect 529094 597744 529150 597800
rect 529218 597744 529274 597800
rect 529342 597744 529398 597800
rect 528970 586294 529026 586350
rect 529094 586294 529150 586350
rect 529218 586294 529274 586350
rect 529342 586294 529398 586350
rect 528970 586170 529026 586226
rect 529094 586170 529150 586226
rect 529218 586170 529274 586226
rect 529342 586170 529398 586226
rect 528970 586046 529026 586102
rect 529094 586046 529150 586102
rect 529218 586046 529274 586102
rect 529342 586046 529398 586102
rect 528970 585922 529026 585978
rect 529094 585922 529150 585978
rect 529218 585922 529274 585978
rect 529342 585922 529398 585978
rect 528970 568294 529026 568350
rect 529094 568294 529150 568350
rect 529218 568294 529274 568350
rect 529342 568294 529398 568350
rect 528970 568170 529026 568226
rect 529094 568170 529150 568226
rect 529218 568170 529274 568226
rect 529342 568170 529398 568226
rect 528970 568046 529026 568102
rect 529094 568046 529150 568102
rect 529218 568046 529274 568102
rect 529342 568046 529398 568102
rect 528970 567922 529026 567978
rect 529094 567922 529150 567978
rect 529218 567922 529274 567978
rect 529342 567922 529398 567978
rect 528970 550294 529026 550350
rect 529094 550294 529150 550350
rect 529218 550294 529274 550350
rect 529342 550294 529398 550350
rect 528970 550170 529026 550226
rect 529094 550170 529150 550226
rect 529218 550170 529274 550226
rect 529342 550170 529398 550226
rect 528970 550046 529026 550102
rect 529094 550046 529150 550102
rect 529218 550046 529274 550102
rect 529342 550046 529398 550102
rect 528970 549922 529026 549978
rect 529094 549922 529150 549978
rect 529218 549922 529274 549978
rect 529342 549922 529398 549978
rect 528970 532294 529026 532350
rect 529094 532294 529150 532350
rect 529218 532294 529274 532350
rect 529342 532294 529398 532350
rect 528970 532170 529026 532226
rect 529094 532170 529150 532226
rect 529218 532170 529274 532226
rect 529342 532170 529398 532226
rect 528970 532046 529026 532102
rect 529094 532046 529150 532102
rect 529218 532046 529274 532102
rect 529342 532046 529398 532102
rect 528970 531922 529026 531978
rect 529094 531922 529150 531978
rect 529218 531922 529274 531978
rect 529342 531922 529398 531978
rect 528970 514294 529026 514350
rect 529094 514294 529150 514350
rect 529218 514294 529274 514350
rect 529342 514294 529398 514350
rect 528970 514170 529026 514226
rect 529094 514170 529150 514226
rect 529218 514170 529274 514226
rect 529342 514170 529398 514226
rect 528970 514046 529026 514102
rect 529094 514046 529150 514102
rect 529218 514046 529274 514102
rect 529342 514046 529398 514102
rect 528970 513922 529026 513978
rect 529094 513922 529150 513978
rect 529218 513922 529274 513978
rect 529342 513922 529398 513978
rect 528970 496294 529026 496350
rect 529094 496294 529150 496350
rect 529218 496294 529274 496350
rect 529342 496294 529398 496350
rect 528970 496170 529026 496226
rect 529094 496170 529150 496226
rect 529218 496170 529274 496226
rect 529342 496170 529398 496226
rect 528970 496046 529026 496102
rect 529094 496046 529150 496102
rect 529218 496046 529274 496102
rect 529342 496046 529398 496102
rect 528970 495922 529026 495978
rect 529094 495922 529150 495978
rect 529218 495922 529274 495978
rect 529342 495922 529398 495978
rect 528970 478294 529026 478350
rect 529094 478294 529150 478350
rect 529218 478294 529274 478350
rect 529342 478294 529398 478350
rect 528970 478170 529026 478226
rect 529094 478170 529150 478226
rect 529218 478170 529274 478226
rect 529342 478170 529398 478226
rect 528970 478046 529026 478102
rect 529094 478046 529150 478102
rect 529218 478046 529274 478102
rect 529342 478046 529398 478102
rect 528970 477922 529026 477978
rect 529094 477922 529150 477978
rect 529218 477922 529274 477978
rect 529342 477922 529398 477978
rect 528970 460294 529026 460350
rect 529094 460294 529150 460350
rect 529218 460294 529274 460350
rect 529342 460294 529398 460350
rect 528970 460170 529026 460226
rect 529094 460170 529150 460226
rect 529218 460170 529274 460226
rect 529342 460170 529398 460226
rect 528970 460046 529026 460102
rect 529094 460046 529150 460102
rect 529218 460046 529274 460102
rect 529342 460046 529398 460102
rect 528970 459922 529026 459978
rect 529094 459922 529150 459978
rect 529218 459922 529274 459978
rect 529342 459922 529398 459978
rect 543250 597156 543306 597212
rect 543374 597156 543430 597212
rect 543498 597156 543554 597212
rect 543622 597156 543678 597212
rect 543250 597032 543306 597088
rect 543374 597032 543430 597088
rect 543498 597032 543554 597088
rect 543622 597032 543678 597088
rect 543250 596908 543306 596964
rect 543374 596908 543430 596964
rect 543498 596908 543554 596964
rect 543622 596908 543678 596964
rect 543250 596784 543306 596840
rect 543374 596784 543430 596840
rect 543498 596784 543554 596840
rect 543622 596784 543678 596840
rect 543250 580294 543306 580350
rect 543374 580294 543430 580350
rect 543498 580294 543554 580350
rect 543622 580294 543678 580350
rect 543250 580170 543306 580226
rect 543374 580170 543430 580226
rect 543498 580170 543554 580226
rect 543622 580170 543678 580226
rect 543250 580046 543306 580102
rect 543374 580046 543430 580102
rect 543498 580046 543554 580102
rect 543622 580046 543678 580102
rect 543250 579922 543306 579978
rect 543374 579922 543430 579978
rect 543498 579922 543554 579978
rect 543622 579922 543678 579978
rect 543250 562294 543306 562350
rect 543374 562294 543430 562350
rect 543498 562294 543554 562350
rect 543622 562294 543678 562350
rect 543250 562170 543306 562226
rect 543374 562170 543430 562226
rect 543498 562170 543554 562226
rect 543622 562170 543678 562226
rect 543250 562046 543306 562102
rect 543374 562046 543430 562102
rect 543498 562046 543554 562102
rect 543622 562046 543678 562102
rect 543250 561922 543306 561978
rect 543374 561922 543430 561978
rect 543498 561922 543554 561978
rect 543622 561922 543678 561978
rect 543250 544294 543306 544350
rect 543374 544294 543430 544350
rect 543498 544294 543554 544350
rect 543622 544294 543678 544350
rect 543250 544170 543306 544226
rect 543374 544170 543430 544226
rect 543498 544170 543554 544226
rect 543622 544170 543678 544226
rect 543250 544046 543306 544102
rect 543374 544046 543430 544102
rect 543498 544046 543554 544102
rect 543622 544046 543678 544102
rect 543250 543922 543306 543978
rect 543374 543922 543430 543978
rect 543498 543922 543554 543978
rect 543622 543922 543678 543978
rect 543250 526294 543306 526350
rect 543374 526294 543430 526350
rect 543498 526294 543554 526350
rect 543622 526294 543678 526350
rect 543250 526170 543306 526226
rect 543374 526170 543430 526226
rect 543498 526170 543554 526226
rect 543622 526170 543678 526226
rect 543250 526046 543306 526102
rect 543374 526046 543430 526102
rect 543498 526046 543554 526102
rect 543622 526046 543678 526102
rect 543250 525922 543306 525978
rect 543374 525922 543430 525978
rect 543498 525922 543554 525978
rect 543622 525922 543678 525978
rect 543250 508294 543306 508350
rect 543374 508294 543430 508350
rect 543498 508294 543554 508350
rect 543622 508294 543678 508350
rect 543250 508170 543306 508226
rect 543374 508170 543430 508226
rect 543498 508170 543554 508226
rect 543622 508170 543678 508226
rect 543250 508046 543306 508102
rect 543374 508046 543430 508102
rect 543498 508046 543554 508102
rect 543622 508046 543678 508102
rect 543250 507922 543306 507978
rect 543374 507922 543430 507978
rect 543498 507922 543554 507978
rect 543622 507922 543678 507978
rect 543250 490294 543306 490350
rect 543374 490294 543430 490350
rect 543498 490294 543554 490350
rect 543622 490294 543678 490350
rect 543250 490170 543306 490226
rect 543374 490170 543430 490226
rect 543498 490170 543554 490226
rect 543622 490170 543678 490226
rect 543250 490046 543306 490102
rect 543374 490046 543430 490102
rect 543498 490046 543554 490102
rect 543622 490046 543678 490102
rect 543250 489922 543306 489978
rect 543374 489922 543430 489978
rect 543498 489922 543554 489978
rect 543622 489922 543678 489978
rect 543250 472294 543306 472350
rect 543374 472294 543430 472350
rect 543498 472294 543554 472350
rect 543622 472294 543678 472350
rect 543250 472170 543306 472226
rect 543374 472170 543430 472226
rect 543498 472170 543554 472226
rect 543622 472170 543678 472226
rect 543250 472046 543306 472102
rect 543374 472046 543430 472102
rect 543498 472046 543554 472102
rect 543622 472046 543678 472102
rect 543250 471922 543306 471978
rect 543374 471922 543430 471978
rect 543498 471922 543554 471978
rect 543622 471922 543678 471978
rect 546970 598116 547026 598172
rect 547094 598116 547150 598172
rect 547218 598116 547274 598172
rect 547342 598116 547398 598172
rect 546970 597992 547026 598048
rect 547094 597992 547150 598048
rect 547218 597992 547274 598048
rect 547342 597992 547398 598048
rect 546970 597868 547026 597924
rect 547094 597868 547150 597924
rect 547218 597868 547274 597924
rect 547342 597868 547398 597924
rect 546970 597744 547026 597800
rect 547094 597744 547150 597800
rect 547218 597744 547274 597800
rect 547342 597744 547398 597800
rect 546970 586294 547026 586350
rect 547094 586294 547150 586350
rect 547218 586294 547274 586350
rect 547342 586294 547398 586350
rect 546970 586170 547026 586226
rect 547094 586170 547150 586226
rect 547218 586170 547274 586226
rect 547342 586170 547398 586226
rect 546970 586046 547026 586102
rect 547094 586046 547150 586102
rect 547218 586046 547274 586102
rect 547342 586046 547398 586102
rect 546970 585922 547026 585978
rect 547094 585922 547150 585978
rect 547218 585922 547274 585978
rect 547342 585922 547398 585978
rect 546970 568294 547026 568350
rect 547094 568294 547150 568350
rect 547218 568294 547274 568350
rect 547342 568294 547398 568350
rect 546970 568170 547026 568226
rect 547094 568170 547150 568226
rect 547218 568170 547274 568226
rect 547342 568170 547398 568226
rect 546970 568046 547026 568102
rect 547094 568046 547150 568102
rect 547218 568046 547274 568102
rect 547342 568046 547398 568102
rect 546970 567922 547026 567978
rect 547094 567922 547150 567978
rect 547218 567922 547274 567978
rect 547342 567922 547398 567978
rect 546970 550294 547026 550350
rect 547094 550294 547150 550350
rect 547218 550294 547274 550350
rect 547342 550294 547398 550350
rect 546970 550170 547026 550226
rect 547094 550170 547150 550226
rect 547218 550170 547274 550226
rect 547342 550170 547398 550226
rect 546970 550046 547026 550102
rect 547094 550046 547150 550102
rect 547218 550046 547274 550102
rect 547342 550046 547398 550102
rect 546970 549922 547026 549978
rect 547094 549922 547150 549978
rect 547218 549922 547274 549978
rect 547342 549922 547398 549978
rect 546970 532294 547026 532350
rect 547094 532294 547150 532350
rect 547218 532294 547274 532350
rect 547342 532294 547398 532350
rect 546970 532170 547026 532226
rect 547094 532170 547150 532226
rect 547218 532170 547274 532226
rect 547342 532170 547398 532226
rect 546970 532046 547026 532102
rect 547094 532046 547150 532102
rect 547218 532046 547274 532102
rect 547342 532046 547398 532102
rect 546970 531922 547026 531978
rect 547094 531922 547150 531978
rect 547218 531922 547274 531978
rect 547342 531922 547398 531978
rect 546970 514294 547026 514350
rect 547094 514294 547150 514350
rect 547218 514294 547274 514350
rect 547342 514294 547398 514350
rect 546970 514170 547026 514226
rect 547094 514170 547150 514226
rect 547218 514170 547274 514226
rect 547342 514170 547398 514226
rect 546970 514046 547026 514102
rect 547094 514046 547150 514102
rect 547218 514046 547274 514102
rect 547342 514046 547398 514102
rect 546970 513922 547026 513978
rect 547094 513922 547150 513978
rect 547218 513922 547274 513978
rect 547342 513922 547398 513978
rect 546970 496294 547026 496350
rect 547094 496294 547150 496350
rect 547218 496294 547274 496350
rect 547342 496294 547398 496350
rect 546970 496170 547026 496226
rect 547094 496170 547150 496226
rect 547218 496170 547274 496226
rect 547342 496170 547398 496226
rect 546970 496046 547026 496102
rect 547094 496046 547150 496102
rect 547218 496046 547274 496102
rect 547342 496046 547398 496102
rect 546970 495922 547026 495978
rect 547094 495922 547150 495978
rect 547218 495922 547274 495978
rect 547342 495922 547398 495978
rect 546970 478294 547026 478350
rect 547094 478294 547150 478350
rect 547218 478294 547274 478350
rect 547342 478294 547398 478350
rect 546970 478170 547026 478226
rect 547094 478170 547150 478226
rect 547218 478170 547274 478226
rect 547342 478170 547398 478226
rect 546970 478046 547026 478102
rect 547094 478046 547150 478102
rect 547218 478046 547274 478102
rect 547342 478046 547398 478102
rect 546970 477922 547026 477978
rect 547094 477922 547150 477978
rect 547218 477922 547274 477978
rect 547342 477922 547398 477978
rect 546970 460294 547026 460350
rect 547094 460294 547150 460350
rect 547218 460294 547274 460350
rect 547342 460294 547398 460350
rect 546970 460170 547026 460226
rect 547094 460170 547150 460226
rect 547218 460170 547274 460226
rect 547342 460170 547398 460226
rect 546970 460046 547026 460102
rect 547094 460046 547150 460102
rect 547218 460046 547274 460102
rect 547342 460046 547398 460102
rect 546970 459922 547026 459978
rect 547094 459922 547150 459978
rect 547218 459922 547274 459978
rect 547342 459922 547398 459978
rect 561250 597156 561306 597212
rect 561374 597156 561430 597212
rect 561498 597156 561554 597212
rect 561622 597156 561678 597212
rect 561250 597032 561306 597088
rect 561374 597032 561430 597088
rect 561498 597032 561554 597088
rect 561622 597032 561678 597088
rect 561250 596908 561306 596964
rect 561374 596908 561430 596964
rect 561498 596908 561554 596964
rect 561622 596908 561678 596964
rect 561250 596784 561306 596840
rect 561374 596784 561430 596840
rect 561498 596784 561554 596840
rect 561622 596784 561678 596840
rect 561250 580294 561306 580350
rect 561374 580294 561430 580350
rect 561498 580294 561554 580350
rect 561622 580294 561678 580350
rect 561250 580170 561306 580226
rect 561374 580170 561430 580226
rect 561498 580170 561554 580226
rect 561622 580170 561678 580226
rect 561250 580046 561306 580102
rect 561374 580046 561430 580102
rect 561498 580046 561554 580102
rect 561622 580046 561678 580102
rect 561250 579922 561306 579978
rect 561374 579922 561430 579978
rect 561498 579922 561554 579978
rect 561622 579922 561678 579978
rect 561250 562294 561306 562350
rect 561374 562294 561430 562350
rect 561498 562294 561554 562350
rect 561622 562294 561678 562350
rect 561250 562170 561306 562226
rect 561374 562170 561430 562226
rect 561498 562170 561554 562226
rect 561622 562170 561678 562226
rect 561250 562046 561306 562102
rect 561374 562046 561430 562102
rect 561498 562046 561554 562102
rect 561622 562046 561678 562102
rect 561250 561922 561306 561978
rect 561374 561922 561430 561978
rect 561498 561922 561554 561978
rect 561622 561922 561678 561978
rect 561250 544294 561306 544350
rect 561374 544294 561430 544350
rect 561498 544294 561554 544350
rect 561622 544294 561678 544350
rect 561250 544170 561306 544226
rect 561374 544170 561430 544226
rect 561498 544170 561554 544226
rect 561622 544170 561678 544226
rect 561250 544046 561306 544102
rect 561374 544046 561430 544102
rect 561498 544046 561554 544102
rect 561622 544046 561678 544102
rect 561250 543922 561306 543978
rect 561374 543922 561430 543978
rect 561498 543922 561554 543978
rect 561622 543922 561678 543978
rect 561250 526294 561306 526350
rect 561374 526294 561430 526350
rect 561498 526294 561554 526350
rect 561622 526294 561678 526350
rect 561250 526170 561306 526226
rect 561374 526170 561430 526226
rect 561498 526170 561554 526226
rect 561622 526170 561678 526226
rect 561250 526046 561306 526102
rect 561374 526046 561430 526102
rect 561498 526046 561554 526102
rect 561622 526046 561678 526102
rect 561250 525922 561306 525978
rect 561374 525922 561430 525978
rect 561498 525922 561554 525978
rect 561622 525922 561678 525978
rect 561250 508294 561306 508350
rect 561374 508294 561430 508350
rect 561498 508294 561554 508350
rect 561622 508294 561678 508350
rect 561250 508170 561306 508226
rect 561374 508170 561430 508226
rect 561498 508170 561554 508226
rect 561622 508170 561678 508226
rect 561250 508046 561306 508102
rect 561374 508046 561430 508102
rect 561498 508046 561554 508102
rect 561622 508046 561678 508102
rect 561250 507922 561306 507978
rect 561374 507922 561430 507978
rect 561498 507922 561554 507978
rect 561622 507922 561678 507978
rect 561250 490294 561306 490350
rect 561374 490294 561430 490350
rect 561498 490294 561554 490350
rect 561622 490294 561678 490350
rect 561250 490170 561306 490226
rect 561374 490170 561430 490226
rect 561498 490170 561554 490226
rect 561622 490170 561678 490226
rect 561250 490046 561306 490102
rect 561374 490046 561430 490102
rect 561498 490046 561554 490102
rect 561622 490046 561678 490102
rect 561250 489922 561306 489978
rect 561374 489922 561430 489978
rect 561498 489922 561554 489978
rect 561622 489922 561678 489978
rect 561250 472294 561306 472350
rect 561374 472294 561430 472350
rect 561498 472294 561554 472350
rect 561622 472294 561678 472350
rect 561250 472170 561306 472226
rect 561374 472170 561430 472226
rect 561498 472170 561554 472226
rect 561622 472170 561678 472226
rect 561250 472046 561306 472102
rect 561374 472046 561430 472102
rect 561498 472046 561554 472102
rect 561622 472046 561678 472102
rect 561250 471922 561306 471978
rect 561374 471922 561430 471978
rect 561498 471922 561554 471978
rect 561622 471922 561678 471978
rect 564970 598116 565026 598172
rect 565094 598116 565150 598172
rect 565218 598116 565274 598172
rect 565342 598116 565398 598172
rect 564970 597992 565026 598048
rect 565094 597992 565150 598048
rect 565218 597992 565274 598048
rect 565342 597992 565398 598048
rect 564970 597868 565026 597924
rect 565094 597868 565150 597924
rect 565218 597868 565274 597924
rect 565342 597868 565398 597924
rect 564970 597744 565026 597800
rect 565094 597744 565150 597800
rect 565218 597744 565274 597800
rect 565342 597744 565398 597800
rect 564970 586294 565026 586350
rect 565094 586294 565150 586350
rect 565218 586294 565274 586350
rect 565342 586294 565398 586350
rect 564970 586170 565026 586226
rect 565094 586170 565150 586226
rect 565218 586170 565274 586226
rect 565342 586170 565398 586226
rect 564970 586046 565026 586102
rect 565094 586046 565150 586102
rect 565218 586046 565274 586102
rect 565342 586046 565398 586102
rect 564970 585922 565026 585978
rect 565094 585922 565150 585978
rect 565218 585922 565274 585978
rect 565342 585922 565398 585978
rect 564970 568294 565026 568350
rect 565094 568294 565150 568350
rect 565218 568294 565274 568350
rect 565342 568294 565398 568350
rect 564970 568170 565026 568226
rect 565094 568170 565150 568226
rect 565218 568170 565274 568226
rect 565342 568170 565398 568226
rect 564970 568046 565026 568102
rect 565094 568046 565150 568102
rect 565218 568046 565274 568102
rect 565342 568046 565398 568102
rect 564970 567922 565026 567978
rect 565094 567922 565150 567978
rect 565218 567922 565274 567978
rect 565342 567922 565398 567978
rect 564970 550294 565026 550350
rect 565094 550294 565150 550350
rect 565218 550294 565274 550350
rect 565342 550294 565398 550350
rect 564970 550170 565026 550226
rect 565094 550170 565150 550226
rect 565218 550170 565274 550226
rect 565342 550170 565398 550226
rect 564970 550046 565026 550102
rect 565094 550046 565150 550102
rect 565218 550046 565274 550102
rect 565342 550046 565398 550102
rect 564970 549922 565026 549978
rect 565094 549922 565150 549978
rect 565218 549922 565274 549978
rect 565342 549922 565398 549978
rect 564970 532294 565026 532350
rect 565094 532294 565150 532350
rect 565218 532294 565274 532350
rect 565342 532294 565398 532350
rect 564970 532170 565026 532226
rect 565094 532170 565150 532226
rect 565218 532170 565274 532226
rect 565342 532170 565398 532226
rect 564970 532046 565026 532102
rect 565094 532046 565150 532102
rect 565218 532046 565274 532102
rect 565342 532046 565398 532102
rect 564970 531922 565026 531978
rect 565094 531922 565150 531978
rect 565218 531922 565274 531978
rect 565342 531922 565398 531978
rect 564970 514294 565026 514350
rect 565094 514294 565150 514350
rect 565218 514294 565274 514350
rect 565342 514294 565398 514350
rect 564970 514170 565026 514226
rect 565094 514170 565150 514226
rect 565218 514170 565274 514226
rect 565342 514170 565398 514226
rect 564970 514046 565026 514102
rect 565094 514046 565150 514102
rect 565218 514046 565274 514102
rect 565342 514046 565398 514102
rect 564970 513922 565026 513978
rect 565094 513922 565150 513978
rect 565218 513922 565274 513978
rect 565342 513922 565398 513978
rect 564970 496294 565026 496350
rect 565094 496294 565150 496350
rect 565218 496294 565274 496350
rect 565342 496294 565398 496350
rect 564970 496170 565026 496226
rect 565094 496170 565150 496226
rect 565218 496170 565274 496226
rect 565342 496170 565398 496226
rect 564970 496046 565026 496102
rect 565094 496046 565150 496102
rect 565218 496046 565274 496102
rect 565342 496046 565398 496102
rect 564970 495922 565026 495978
rect 565094 495922 565150 495978
rect 565218 495922 565274 495978
rect 565342 495922 565398 495978
rect 564970 478294 565026 478350
rect 565094 478294 565150 478350
rect 565218 478294 565274 478350
rect 565342 478294 565398 478350
rect 564970 478170 565026 478226
rect 565094 478170 565150 478226
rect 565218 478170 565274 478226
rect 565342 478170 565398 478226
rect 564970 478046 565026 478102
rect 565094 478046 565150 478102
rect 565218 478046 565274 478102
rect 565342 478046 565398 478102
rect 564970 477922 565026 477978
rect 565094 477922 565150 477978
rect 565218 477922 565274 477978
rect 565342 477922 565398 477978
rect 564970 460294 565026 460350
rect 565094 460294 565150 460350
rect 565218 460294 565274 460350
rect 565342 460294 565398 460350
rect 564970 460170 565026 460226
rect 565094 460170 565150 460226
rect 565218 460170 565274 460226
rect 565342 460170 565398 460226
rect 564970 460046 565026 460102
rect 565094 460046 565150 460102
rect 565218 460046 565274 460102
rect 565342 460046 565398 460102
rect 564970 459922 565026 459978
rect 565094 459922 565150 459978
rect 565218 459922 565274 459978
rect 565342 459922 565398 459978
rect 579250 597156 579306 597212
rect 579374 597156 579430 597212
rect 579498 597156 579554 597212
rect 579622 597156 579678 597212
rect 579250 597032 579306 597088
rect 579374 597032 579430 597088
rect 579498 597032 579554 597088
rect 579622 597032 579678 597088
rect 579250 596908 579306 596964
rect 579374 596908 579430 596964
rect 579498 596908 579554 596964
rect 579622 596908 579678 596964
rect 579250 596784 579306 596840
rect 579374 596784 579430 596840
rect 579498 596784 579554 596840
rect 579622 596784 579678 596840
rect 579250 580294 579306 580350
rect 579374 580294 579430 580350
rect 579498 580294 579554 580350
rect 579622 580294 579678 580350
rect 579250 580170 579306 580226
rect 579374 580170 579430 580226
rect 579498 580170 579554 580226
rect 579622 580170 579678 580226
rect 579250 580046 579306 580102
rect 579374 580046 579430 580102
rect 579498 580046 579554 580102
rect 579622 580046 579678 580102
rect 579250 579922 579306 579978
rect 579374 579922 579430 579978
rect 579498 579922 579554 579978
rect 579622 579922 579678 579978
rect 579250 562294 579306 562350
rect 579374 562294 579430 562350
rect 579498 562294 579554 562350
rect 579622 562294 579678 562350
rect 579250 562170 579306 562226
rect 579374 562170 579430 562226
rect 579498 562170 579554 562226
rect 579622 562170 579678 562226
rect 579250 562046 579306 562102
rect 579374 562046 579430 562102
rect 579498 562046 579554 562102
rect 579622 562046 579678 562102
rect 579250 561922 579306 561978
rect 579374 561922 579430 561978
rect 579498 561922 579554 561978
rect 579622 561922 579678 561978
rect 579250 544294 579306 544350
rect 579374 544294 579430 544350
rect 579498 544294 579554 544350
rect 579622 544294 579678 544350
rect 579250 544170 579306 544226
rect 579374 544170 579430 544226
rect 579498 544170 579554 544226
rect 579622 544170 579678 544226
rect 579250 544046 579306 544102
rect 579374 544046 579430 544102
rect 579498 544046 579554 544102
rect 579622 544046 579678 544102
rect 579250 543922 579306 543978
rect 579374 543922 579430 543978
rect 579498 543922 579554 543978
rect 579622 543922 579678 543978
rect 579250 526294 579306 526350
rect 579374 526294 579430 526350
rect 579498 526294 579554 526350
rect 579622 526294 579678 526350
rect 579250 526170 579306 526226
rect 579374 526170 579430 526226
rect 579498 526170 579554 526226
rect 579622 526170 579678 526226
rect 579250 526046 579306 526102
rect 579374 526046 579430 526102
rect 579498 526046 579554 526102
rect 579622 526046 579678 526102
rect 579250 525922 579306 525978
rect 579374 525922 579430 525978
rect 579498 525922 579554 525978
rect 579622 525922 579678 525978
rect 579250 508294 579306 508350
rect 579374 508294 579430 508350
rect 579498 508294 579554 508350
rect 579622 508294 579678 508350
rect 579250 508170 579306 508226
rect 579374 508170 579430 508226
rect 579498 508170 579554 508226
rect 579622 508170 579678 508226
rect 579250 508046 579306 508102
rect 579374 508046 579430 508102
rect 579498 508046 579554 508102
rect 579622 508046 579678 508102
rect 579250 507922 579306 507978
rect 579374 507922 579430 507978
rect 579498 507922 579554 507978
rect 579622 507922 579678 507978
rect 579250 490294 579306 490350
rect 579374 490294 579430 490350
rect 579498 490294 579554 490350
rect 579622 490294 579678 490350
rect 579250 490170 579306 490226
rect 579374 490170 579430 490226
rect 579498 490170 579554 490226
rect 579622 490170 579678 490226
rect 579250 490046 579306 490102
rect 579374 490046 579430 490102
rect 579498 490046 579554 490102
rect 579622 490046 579678 490102
rect 579250 489922 579306 489978
rect 579374 489922 579430 489978
rect 579498 489922 579554 489978
rect 579622 489922 579678 489978
rect 579250 472294 579306 472350
rect 579374 472294 579430 472350
rect 579498 472294 579554 472350
rect 579622 472294 579678 472350
rect 579250 472170 579306 472226
rect 579374 472170 579430 472226
rect 579498 472170 579554 472226
rect 579622 472170 579678 472226
rect 579250 472046 579306 472102
rect 579374 472046 579430 472102
rect 579498 472046 579554 472102
rect 579622 472046 579678 472102
rect 579250 471922 579306 471978
rect 579374 471922 579430 471978
rect 579498 471922 579554 471978
rect 579622 471922 579678 471978
rect 402970 442294 403026 442350
rect 403094 442294 403150 442350
rect 403218 442294 403274 442350
rect 403342 442294 403398 442350
rect 402970 442170 403026 442226
rect 403094 442170 403150 442226
rect 403218 442170 403274 442226
rect 403342 442170 403398 442226
rect 402970 442046 403026 442102
rect 403094 442046 403150 442102
rect 403218 442046 403274 442102
rect 403342 442046 403398 442102
rect 402970 441922 403026 441978
rect 403094 441922 403150 441978
rect 403218 441922 403274 441978
rect 403342 441922 403398 441978
rect 402970 424294 403026 424350
rect 403094 424294 403150 424350
rect 403218 424294 403274 424350
rect 403342 424294 403398 424350
rect 402970 424170 403026 424226
rect 403094 424170 403150 424226
rect 403218 424170 403274 424226
rect 403342 424170 403398 424226
rect 402970 424046 403026 424102
rect 403094 424046 403150 424102
rect 403218 424046 403274 424102
rect 403342 424046 403398 424102
rect 402970 423922 403026 423978
rect 403094 423922 403150 423978
rect 403218 423922 403274 423978
rect 403342 423922 403398 423978
rect 402970 406294 403026 406350
rect 403094 406294 403150 406350
rect 403218 406294 403274 406350
rect 403342 406294 403398 406350
rect 402970 406170 403026 406226
rect 403094 406170 403150 406226
rect 403218 406170 403274 406226
rect 403342 406170 403398 406226
rect 402970 406046 403026 406102
rect 403094 406046 403150 406102
rect 403218 406046 403274 406102
rect 403342 406046 403398 406102
rect 402970 405922 403026 405978
rect 403094 405922 403150 405978
rect 403218 405922 403274 405978
rect 403342 405922 403398 405978
rect 402970 388294 403026 388350
rect 403094 388294 403150 388350
rect 403218 388294 403274 388350
rect 403342 388294 403398 388350
rect 402970 388170 403026 388226
rect 403094 388170 403150 388226
rect 403218 388170 403274 388226
rect 403342 388170 403398 388226
rect 402970 388046 403026 388102
rect 403094 388046 403150 388102
rect 403218 388046 403274 388102
rect 403342 388046 403398 388102
rect 402970 387922 403026 387978
rect 403094 387922 403150 387978
rect 403218 387922 403274 387978
rect 403342 387922 403398 387978
rect 402970 370294 403026 370350
rect 403094 370294 403150 370350
rect 403218 370294 403274 370350
rect 403342 370294 403398 370350
rect 402970 370170 403026 370226
rect 403094 370170 403150 370226
rect 403218 370170 403274 370226
rect 403342 370170 403398 370226
rect 402970 370046 403026 370102
rect 403094 370046 403150 370102
rect 403218 370046 403274 370102
rect 403342 370046 403398 370102
rect 402970 369922 403026 369978
rect 403094 369922 403150 369978
rect 403218 369922 403274 369978
rect 403342 369922 403398 369978
rect 402970 352294 403026 352350
rect 403094 352294 403150 352350
rect 403218 352294 403274 352350
rect 403342 352294 403398 352350
rect 402970 352170 403026 352226
rect 403094 352170 403150 352226
rect 403218 352170 403274 352226
rect 403342 352170 403398 352226
rect 402970 352046 403026 352102
rect 403094 352046 403150 352102
rect 403218 352046 403274 352102
rect 403342 352046 403398 352102
rect 402970 351922 403026 351978
rect 403094 351922 403150 351978
rect 403218 351922 403274 351978
rect 403342 351922 403398 351978
rect 402970 334294 403026 334350
rect 403094 334294 403150 334350
rect 403218 334294 403274 334350
rect 403342 334294 403398 334350
rect 402970 334170 403026 334226
rect 403094 334170 403150 334226
rect 403218 334170 403274 334226
rect 403342 334170 403398 334226
rect 402970 334046 403026 334102
rect 403094 334046 403150 334102
rect 403218 334046 403274 334102
rect 403342 334046 403398 334102
rect 402970 333922 403026 333978
rect 403094 333922 403150 333978
rect 403218 333922 403274 333978
rect 403342 333922 403398 333978
rect 579250 454294 579306 454350
rect 579374 454294 579430 454350
rect 579498 454294 579554 454350
rect 579622 454294 579678 454350
rect 579250 454170 579306 454226
rect 579374 454170 579430 454226
rect 579498 454170 579554 454226
rect 579622 454170 579678 454226
rect 579250 454046 579306 454102
rect 579374 454046 579430 454102
rect 579498 454046 579554 454102
rect 579622 454046 579678 454102
rect 579250 453922 579306 453978
rect 579374 453922 579430 453978
rect 579498 453922 579554 453978
rect 579622 453922 579678 453978
rect 579250 436294 579306 436350
rect 579374 436294 579430 436350
rect 579498 436294 579554 436350
rect 579622 436294 579678 436350
rect 579250 436170 579306 436226
rect 579374 436170 579430 436226
rect 579498 436170 579554 436226
rect 579622 436170 579678 436226
rect 579250 436046 579306 436102
rect 579374 436046 579430 436102
rect 579498 436046 579554 436102
rect 579622 436046 579678 436102
rect 579250 435922 579306 435978
rect 579374 435922 579430 435978
rect 579498 435922 579554 435978
rect 579622 435922 579678 435978
rect 579250 418294 579306 418350
rect 579374 418294 579430 418350
rect 579498 418294 579554 418350
rect 579622 418294 579678 418350
rect 579250 418170 579306 418226
rect 579374 418170 579430 418226
rect 579498 418170 579554 418226
rect 579622 418170 579678 418226
rect 579250 418046 579306 418102
rect 579374 418046 579430 418102
rect 579498 418046 579554 418102
rect 579622 418046 579678 418102
rect 579250 417922 579306 417978
rect 579374 417922 579430 417978
rect 579498 417922 579554 417978
rect 579622 417922 579678 417978
rect 579250 400294 579306 400350
rect 579374 400294 579430 400350
rect 579498 400294 579554 400350
rect 579622 400294 579678 400350
rect 579250 400170 579306 400226
rect 579374 400170 579430 400226
rect 579498 400170 579554 400226
rect 579622 400170 579678 400226
rect 579250 400046 579306 400102
rect 579374 400046 579430 400102
rect 579498 400046 579554 400102
rect 579622 400046 579678 400102
rect 579250 399922 579306 399978
rect 579374 399922 579430 399978
rect 579498 399922 579554 399978
rect 579622 399922 579678 399978
rect 579250 382294 579306 382350
rect 579374 382294 579430 382350
rect 579498 382294 579554 382350
rect 579622 382294 579678 382350
rect 579250 382170 579306 382226
rect 579374 382170 579430 382226
rect 579498 382170 579554 382226
rect 579622 382170 579678 382226
rect 579250 382046 579306 382102
rect 579374 382046 579430 382102
rect 579498 382046 579554 382102
rect 579622 382046 579678 382102
rect 579250 381922 579306 381978
rect 579374 381922 579430 381978
rect 579498 381922 579554 381978
rect 579622 381922 579678 381978
rect 579250 364294 579306 364350
rect 579374 364294 579430 364350
rect 579498 364294 579554 364350
rect 579622 364294 579678 364350
rect 579250 364170 579306 364226
rect 579374 364170 579430 364226
rect 579498 364170 579554 364226
rect 579622 364170 579678 364226
rect 579250 364046 579306 364102
rect 579374 364046 579430 364102
rect 579498 364046 579554 364102
rect 579622 364046 579678 364102
rect 579250 363922 579306 363978
rect 579374 363922 579430 363978
rect 579498 363922 579554 363978
rect 579622 363922 579678 363978
rect 579250 346294 579306 346350
rect 579374 346294 579430 346350
rect 579498 346294 579554 346350
rect 579622 346294 579678 346350
rect 579250 346170 579306 346226
rect 579374 346170 579430 346226
rect 579498 346170 579554 346226
rect 579622 346170 579678 346226
rect 579250 346046 579306 346102
rect 579374 346046 579430 346102
rect 579498 346046 579554 346102
rect 579622 346046 579678 346102
rect 579250 345922 579306 345978
rect 579374 345922 579430 345978
rect 579498 345922 579554 345978
rect 579622 345922 579678 345978
rect 579250 328294 579306 328350
rect 579374 328294 579430 328350
rect 579498 328294 579554 328350
rect 579622 328294 579678 328350
rect 579250 328170 579306 328226
rect 579374 328170 579430 328226
rect 579498 328170 579554 328226
rect 579622 328170 579678 328226
rect 579250 328046 579306 328102
rect 579374 328046 579430 328102
rect 579498 328046 579554 328102
rect 579622 328046 579678 328102
rect 579250 327922 579306 327978
rect 579374 327922 579430 327978
rect 579498 327922 579554 327978
rect 579622 327922 579678 327978
rect 402970 316294 403026 316350
rect 403094 316294 403150 316350
rect 403218 316294 403274 316350
rect 403342 316294 403398 316350
rect 402970 316170 403026 316226
rect 403094 316170 403150 316226
rect 403218 316170 403274 316226
rect 403342 316170 403398 316226
rect 402970 316046 403026 316102
rect 403094 316046 403150 316102
rect 403218 316046 403274 316102
rect 403342 316046 403398 316102
rect 402970 315922 403026 315978
rect 403094 315922 403150 315978
rect 403218 315922 403274 315978
rect 403342 315922 403398 315978
rect 402970 298294 403026 298350
rect 403094 298294 403150 298350
rect 403218 298294 403274 298350
rect 403342 298294 403398 298350
rect 420970 316294 421026 316350
rect 421094 316294 421150 316350
rect 421218 316294 421274 316350
rect 421342 316294 421398 316350
rect 420970 316170 421026 316226
rect 421094 316170 421150 316226
rect 421218 316170 421274 316226
rect 421342 316170 421398 316226
rect 420970 316046 421026 316102
rect 421094 316046 421150 316102
rect 421218 316046 421274 316102
rect 421342 316046 421398 316102
rect 420970 315922 421026 315978
rect 421094 315922 421150 315978
rect 421218 315922 421274 315978
rect 421342 315922 421398 315978
rect 420970 298366 421026 298422
rect 421094 298366 421150 298422
rect 421218 298366 421274 298422
rect 421342 298366 421398 298422
rect 438970 316294 439026 316350
rect 439094 316294 439150 316350
rect 439218 316294 439274 316350
rect 439342 316294 439398 316350
rect 438970 316170 439026 316226
rect 439094 316170 439150 316226
rect 439218 316170 439274 316226
rect 439342 316170 439398 316226
rect 438970 316046 439026 316102
rect 439094 316046 439150 316102
rect 439218 316046 439274 316102
rect 439342 316046 439398 316102
rect 438970 315922 439026 315978
rect 439094 315922 439150 315978
rect 439218 315922 439274 315978
rect 439342 315922 439398 315978
rect 438970 298366 439026 298422
rect 439094 298366 439150 298422
rect 439218 298366 439274 298422
rect 439342 298366 439398 298422
rect 456970 316294 457026 316350
rect 457094 316294 457150 316350
rect 457218 316294 457274 316350
rect 457342 316294 457398 316350
rect 456970 316170 457026 316226
rect 457094 316170 457150 316226
rect 457218 316170 457274 316226
rect 457342 316170 457398 316226
rect 456970 316046 457026 316102
rect 457094 316046 457150 316102
rect 457218 316046 457274 316102
rect 457342 316046 457398 316102
rect 456970 315922 457026 315978
rect 457094 315922 457150 315978
rect 457218 315922 457274 315978
rect 457342 315922 457398 315978
rect 456970 298366 457026 298422
rect 457094 298366 457150 298422
rect 457218 298366 457274 298422
rect 457342 298366 457398 298422
rect 474970 316294 475026 316350
rect 475094 316294 475150 316350
rect 475218 316294 475274 316350
rect 475342 316294 475398 316350
rect 474970 316170 475026 316226
rect 475094 316170 475150 316226
rect 475218 316170 475274 316226
rect 475342 316170 475398 316226
rect 474970 316046 475026 316102
rect 475094 316046 475150 316102
rect 475218 316046 475274 316102
rect 475342 316046 475398 316102
rect 474970 315922 475026 315978
rect 475094 315922 475150 315978
rect 475218 315922 475274 315978
rect 475342 315922 475398 315978
rect 474970 298366 475026 298422
rect 475094 298366 475150 298422
rect 475218 298366 475274 298422
rect 475342 298366 475398 298422
rect 492970 316294 493026 316350
rect 493094 316294 493150 316350
rect 493218 316294 493274 316350
rect 493342 316294 493398 316350
rect 492970 316170 493026 316226
rect 493094 316170 493150 316226
rect 493218 316170 493274 316226
rect 493342 316170 493398 316226
rect 492970 316046 493026 316102
rect 493094 316046 493150 316102
rect 493218 316046 493274 316102
rect 493342 316046 493398 316102
rect 492970 315922 493026 315978
rect 493094 315922 493150 315978
rect 493218 315922 493274 315978
rect 493342 315922 493398 315978
rect 492970 298366 493026 298422
rect 493094 298366 493150 298422
rect 493218 298366 493274 298422
rect 493342 298366 493398 298422
rect 510970 316294 511026 316350
rect 511094 316294 511150 316350
rect 511218 316294 511274 316350
rect 511342 316294 511398 316350
rect 510970 316170 511026 316226
rect 511094 316170 511150 316226
rect 511218 316170 511274 316226
rect 511342 316170 511398 316226
rect 510970 316046 511026 316102
rect 511094 316046 511150 316102
rect 511218 316046 511274 316102
rect 511342 316046 511398 316102
rect 510970 315922 511026 315978
rect 511094 315922 511150 315978
rect 511218 315922 511274 315978
rect 511342 315922 511398 315978
rect 510970 298366 511026 298422
rect 511094 298366 511150 298422
rect 511218 298366 511274 298422
rect 511342 298366 511398 298422
rect 528970 316294 529026 316350
rect 529094 316294 529150 316350
rect 529218 316294 529274 316350
rect 529342 316294 529398 316350
rect 528970 316170 529026 316226
rect 529094 316170 529150 316226
rect 529218 316170 529274 316226
rect 529342 316170 529398 316226
rect 528970 316046 529026 316102
rect 529094 316046 529150 316102
rect 529218 316046 529274 316102
rect 529342 316046 529398 316102
rect 528970 315922 529026 315978
rect 529094 315922 529150 315978
rect 529218 315922 529274 315978
rect 529342 315922 529398 315978
rect 528970 298366 529026 298422
rect 529094 298366 529150 298422
rect 529218 298366 529274 298422
rect 529342 298366 529398 298422
rect 546970 316294 547026 316350
rect 547094 316294 547150 316350
rect 547218 316294 547274 316350
rect 547342 316294 547398 316350
rect 546970 316170 547026 316226
rect 547094 316170 547150 316226
rect 547218 316170 547274 316226
rect 547342 316170 547398 316226
rect 546970 316046 547026 316102
rect 547094 316046 547150 316102
rect 547218 316046 547274 316102
rect 547342 316046 547398 316102
rect 546970 315922 547026 315978
rect 547094 315922 547150 315978
rect 547218 315922 547274 315978
rect 547342 315922 547398 315978
rect 546970 298366 547026 298422
rect 547094 298366 547150 298422
rect 547218 298366 547274 298422
rect 547342 298366 547398 298422
rect 564970 316294 565026 316350
rect 565094 316294 565150 316350
rect 565218 316294 565274 316350
rect 565342 316294 565398 316350
rect 564970 316170 565026 316226
rect 565094 316170 565150 316226
rect 565218 316170 565274 316226
rect 565342 316170 565398 316226
rect 564970 316046 565026 316102
rect 565094 316046 565150 316102
rect 565218 316046 565274 316102
rect 565342 316046 565398 316102
rect 564970 315922 565026 315978
rect 565094 315922 565150 315978
rect 565218 315922 565274 315978
rect 565342 315922 565398 315978
rect 564970 298366 565026 298422
rect 565094 298366 565150 298422
rect 565218 298366 565274 298422
rect 565342 298366 565398 298422
rect 579250 310294 579306 310350
rect 579374 310294 579430 310350
rect 579498 310294 579554 310350
rect 579622 310294 579678 310350
rect 579250 310170 579306 310226
rect 579374 310170 579430 310226
rect 579498 310170 579554 310226
rect 579622 310170 579678 310226
rect 579250 310046 579306 310102
rect 579374 310046 579430 310102
rect 579498 310046 579554 310102
rect 579622 310046 579678 310102
rect 579250 309922 579306 309978
rect 579374 309922 579430 309978
rect 579498 309922 579554 309978
rect 579622 309922 579678 309978
rect 402970 298170 403026 298226
rect 403094 298170 403150 298226
rect 403218 298170 403274 298226
rect 403342 298170 403398 298226
rect 402970 298046 403026 298102
rect 403094 298046 403150 298102
rect 403218 298046 403274 298102
rect 403342 298046 403398 298102
rect 402970 297922 403026 297978
rect 403094 297922 403150 297978
rect 403218 297922 403274 297978
rect 403342 297922 403398 297978
rect 402970 280294 403026 280350
rect 403094 280294 403150 280350
rect 403218 280294 403274 280350
rect 403342 280294 403398 280350
rect 402970 280170 403026 280226
rect 403094 280170 403150 280226
rect 403218 280170 403274 280226
rect 403342 280170 403398 280226
rect 402970 280046 403026 280102
rect 403094 280046 403150 280102
rect 403218 280046 403274 280102
rect 403342 280046 403398 280102
rect 402970 279922 403026 279978
rect 403094 279922 403150 279978
rect 403218 279922 403274 279978
rect 403342 279922 403398 279978
rect 402970 262294 403026 262350
rect 403094 262294 403150 262350
rect 403218 262294 403274 262350
rect 403342 262294 403398 262350
rect 402970 262170 403026 262226
rect 403094 262170 403150 262226
rect 403218 262170 403274 262226
rect 403342 262170 403398 262226
rect 402970 262046 403026 262102
rect 403094 262046 403150 262102
rect 403218 262046 403274 262102
rect 403342 262046 403398 262102
rect 402970 261922 403026 261978
rect 403094 261922 403150 261978
rect 403218 261922 403274 261978
rect 403342 261922 403398 261978
rect 402970 244294 403026 244350
rect 403094 244294 403150 244350
rect 403218 244294 403274 244350
rect 403342 244294 403398 244350
rect 402970 244170 403026 244226
rect 403094 244170 403150 244226
rect 403218 244170 403274 244226
rect 403342 244170 403398 244226
rect 402970 244046 403026 244102
rect 403094 244046 403150 244102
rect 403218 244046 403274 244102
rect 403342 244046 403398 244102
rect 402970 243922 403026 243978
rect 403094 243922 403150 243978
rect 403218 243922 403274 243978
rect 403342 243922 403398 243978
rect 402970 226294 403026 226350
rect 403094 226294 403150 226350
rect 403218 226294 403274 226350
rect 403342 226294 403398 226350
rect 402970 226170 403026 226226
rect 403094 226170 403150 226226
rect 403218 226170 403274 226226
rect 403342 226170 403398 226226
rect 402970 226046 403026 226102
rect 403094 226046 403150 226102
rect 403218 226046 403274 226102
rect 403342 226046 403398 226102
rect 402970 225922 403026 225978
rect 403094 225922 403150 225978
rect 403218 225922 403274 225978
rect 403342 225922 403398 225978
rect 402970 208294 403026 208350
rect 403094 208294 403150 208350
rect 403218 208294 403274 208350
rect 403342 208294 403398 208350
rect 402970 208170 403026 208226
rect 403094 208170 403150 208226
rect 403218 208170 403274 208226
rect 403342 208170 403398 208226
rect 402970 208046 403026 208102
rect 403094 208046 403150 208102
rect 403218 208046 403274 208102
rect 403342 208046 403398 208102
rect 402970 207922 403026 207978
rect 403094 207922 403150 207978
rect 403218 207922 403274 207978
rect 403342 207922 403398 207978
rect 402970 190294 403026 190350
rect 403094 190294 403150 190350
rect 403218 190294 403274 190350
rect 403342 190294 403398 190350
rect 402970 190170 403026 190226
rect 403094 190170 403150 190226
rect 403218 190170 403274 190226
rect 403342 190170 403398 190226
rect 402970 190046 403026 190102
rect 403094 190046 403150 190102
rect 403218 190046 403274 190102
rect 403342 190046 403398 190102
rect 402970 189922 403026 189978
rect 403094 189922 403150 189978
rect 403218 189922 403274 189978
rect 403342 189922 403398 189978
rect 402970 172294 403026 172350
rect 403094 172294 403150 172350
rect 403218 172294 403274 172350
rect 403342 172294 403398 172350
rect 402970 172170 403026 172226
rect 403094 172170 403150 172226
rect 403218 172170 403274 172226
rect 403342 172170 403398 172226
rect 402970 172046 403026 172102
rect 403094 172046 403150 172102
rect 403218 172046 403274 172102
rect 403342 172046 403398 172102
rect 402970 171922 403026 171978
rect 403094 171922 403150 171978
rect 403218 171922 403274 171978
rect 403342 171922 403398 171978
rect 579250 292294 579306 292350
rect 579374 292294 579430 292350
rect 579498 292294 579554 292350
rect 579622 292294 579678 292350
rect 579250 292170 579306 292226
rect 579374 292170 579430 292226
rect 579498 292170 579554 292226
rect 579622 292170 579678 292226
rect 579250 292046 579306 292102
rect 579374 292046 579430 292102
rect 579498 292046 579554 292102
rect 579622 292046 579678 292102
rect 579250 291922 579306 291978
rect 579374 291922 579430 291978
rect 579498 291922 579554 291978
rect 579622 291922 579678 291978
rect 579250 274294 579306 274350
rect 579374 274294 579430 274350
rect 579498 274294 579554 274350
rect 579622 274294 579678 274350
rect 579250 274170 579306 274226
rect 579374 274170 579430 274226
rect 579498 274170 579554 274226
rect 579622 274170 579678 274226
rect 579250 274046 579306 274102
rect 579374 274046 579430 274102
rect 579498 274046 579554 274102
rect 579622 274046 579678 274102
rect 579250 273922 579306 273978
rect 579374 273922 579430 273978
rect 579498 273922 579554 273978
rect 579622 273922 579678 273978
rect 579250 256294 579306 256350
rect 579374 256294 579430 256350
rect 579498 256294 579554 256350
rect 579622 256294 579678 256350
rect 579250 256170 579306 256226
rect 579374 256170 579430 256226
rect 579498 256170 579554 256226
rect 579622 256170 579678 256226
rect 579250 256046 579306 256102
rect 579374 256046 579430 256102
rect 579498 256046 579554 256102
rect 579622 256046 579678 256102
rect 579250 255922 579306 255978
rect 579374 255922 579430 255978
rect 579498 255922 579554 255978
rect 579622 255922 579678 255978
rect 579250 238294 579306 238350
rect 579374 238294 579430 238350
rect 579498 238294 579554 238350
rect 579622 238294 579678 238350
rect 579250 238170 579306 238226
rect 579374 238170 579430 238226
rect 579498 238170 579554 238226
rect 579622 238170 579678 238226
rect 579250 238046 579306 238102
rect 579374 238046 579430 238102
rect 579498 238046 579554 238102
rect 579622 238046 579678 238102
rect 579250 237922 579306 237978
rect 579374 237922 579430 237978
rect 579498 237922 579554 237978
rect 579622 237922 579678 237978
rect 579250 220294 579306 220350
rect 579374 220294 579430 220350
rect 579498 220294 579554 220350
rect 579622 220294 579678 220350
rect 579250 220170 579306 220226
rect 579374 220170 579430 220226
rect 579498 220170 579554 220226
rect 579622 220170 579678 220226
rect 579250 220046 579306 220102
rect 579374 220046 579430 220102
rect 579498 220046 579554 220102
rect 579622 220046 579678 220102
rect 579250 219922 579306 219978
rect 579374 219922 579430 219978
rect 579498 219922 579554 219978
rect 579622 219922 579678 219978
rect 579250 202294 579306 202350
rect 579374 202294 579430 202350
rect 579498 202294 579554 202350
rect 579622 202294 579678 202350
rect 579250 202170 579306 202226
rect 579374 202170 579430 202226
rect 579498 202170 579554 202226
rect 579622 202170 579678 202226
rect 579250 202046 579306 202102
rect 579374 202046 579430 202102
rect 579498 202046 579554 202102
rect 579622 202046 579678 202102
rect 579250 201922 579306 201978
rect 579374 201922 579430 201978
rect 579498 201922 579554 201978
rect 579622 201922 579678 201978
rect 579250 184294 579306 184350
rect 579374 184294 579430 184350
rect 579498 184294 579554 184350
rect 579622 184294 579678 184350
rect 579250 184170 579306 184226
rect 579374 184170 579430 184226
rect 579498 184170 579554 184226
rect 579622 184170 579678 184226
rect 579250 184046 579306 184102
rect 579374 184046 579430 184102
rect 579498 184046 579554 184102
rect 579622 184046 579678 184102
rect 579250 183922 579306 183978
rect 579374 183922 579430 183978
rect 579498 183922 579554 183978
rect 579622 183922 579678 183978
rect 579250 166294 579306 166350
rect 579374 166294 579430 166350
rect 579498 166294 579554 166350
rect 579622 166294 579678 166350
rect 579250 166170 579306 166226
rect 579374 166170 579430 166226
rect 579498 166170 579554 166226
rect 579622 166170 579678 166226
rect 579250 166046 579306 166102
rect 579374 166046 579430 166102
rect 579498 166046 579554 166102
rect 579622 166046 579678 166102
rect 579250 165922 579306 165978
rect 579374 165922 579430 165978
rect 579498 165922 579554 165978
rect 579622 165922 579678 165978
rect 402970 154294 403026 154350
rect 403094 154294 403150 154350
rect 403218 154294 403274 154350
rect 403342 154294 403398 154350
rect 402970 154170 403026 154226
rect 403094 154170 403150 154226
rect 403218 154170 403274 154226
rect 403342 154170 403398 154226
rect 402970 154046 403026 154102
rect 403094 154046 403150 154102
rect 403218 154046 403274 154102
rect 403342 154046 403398 154102
rect 402970 153922 403026 153978
rect 403094 153922 403150 153978
rect 403218 153922 403274 153978
rect 403342 153922 403398 153978
rect 402970 136294 403026 136350
rect 403094 136294 403150 136350
rect 403218 136294 403274 136350
rect 403342 136294 403398 136350
rect 402970 136170 403026 136226
rect 403094 136170 403150 136226
rect 403218 136170 403274 136226
rect 403342 136170 403398 136226
rect 402970 136046 403026 136102
rect 403094 136046 403150 136102
rect 403218 136046 403274 136102
rect 403342 136046 403398 136102
rect 402970 135922 403026 135978
rect 403094 135922 403150 135978
rect 403218 135922 403274 135978
rect 403342 135922 403398 135978
rect 402970 118294 403026 118350
rect 403094 118294 403150 118350
rect 403218 118294 403274 118350
rect 403342 118294 403398 118350
rect 402970 118170 403026 118226
rect 403094 118170 403150 118226
rect 403218 118170 403274 118226
rect 403342 118170 403398 118226
rect 402970 118046 403026 118102
rect 403094 118046 403150 118102
rect 403218 118046 403274 118102
rect 403342 118046 403398 118102
rect 402970 117922 403026 117978
rect 403094 117922 403150 117978
rect 403218 117922 403274 117978
rect 403342 117922 403398 117978
rect 402970 100294 403026 100350
rect 403094 100294 403150 100350
rect 403218 100294 403274 100350
rect 403342 100294 403398 100350
rect 402970 100170 403026 100226
rect 403094 100170 403150 100226
rect 403218 100170 403274 100226
rect 403342 100170 403398 100226
rect 402970 100046 403026 100102
rect 403094 100046 403150 100102
rect 403218 100046 403274 100102
rect 403342 100046 403398 100102
rect 402970 99922 403026 99978
rect 403094 99922 403150 99978
rect 403218 99922 403274 99978
rect 403342 99922 403398 99978
rect 402970 82294 403026 82350
rect 403094 82294 403150 82350
rect 403218 82294 403274 82350
rect 403342 82294 403398 82350
rect 402970 82170 403026 82226
rect 403094 82170 403150 82226
rect 403218 82170 403274 82226
rect 403342 82170 403398 82226
rect 402970 82046 403026 82102
rect 403094 82046 403150 82102
rect 403218 82046 403274 82102
rect 403342 82046 403398 82102
rect 402970 81922 403026 81978
rect 403094 81922 403150 81978
rect 403218 81922 403274 81978
rect 403342 81922 403398 81978
rect 402970 64294 403026 64350
rect 403094 64294 403150 64350
rect 403218 64294 403274 64350
rect 403342 64294 403398 64350
rect 402970 64170 403026 64226
rect 403094 64170 403150 64226
rect 403218 64170 403274 64226
rect 403342 64170 403398 64226
rect 402970 64046 403026 64102
rect 403094 64046 403150 64102
rect 403218 64046 403274 64102
rect 403342 64046 403398 64102
rect 402970 63922 403026 63978
rect 403094 63922 403150 63978
rect 403218 63922 403274 63978
rect 403342 63922 403398 63978
rect 402970 46294 403026 46350
rect 403094 46294 403150 46350
rect 403218 46294 403274 46350
rect 403342 46294 403398 46350
rect 402970 46170 403026 46226
rect 403094 46170 403150 46226
rect 403218 46170 403274 46226
rect 403342 46170 403398 46226
rect 402970 46046 403026 46102
rect 403094 46046 403150 46102
rect 403218 46046 403274 46102
rect 403342 46046 403398 46102
rect 402970 45922 403026 45978
rect 403094 45922 403150 45978
rect 403218 45922 403274 45978
rect 403342 45922 403398 45978
rect 402970 28294 403026 28350
rect 403094 28294 403150 28350
rect 403218 28294 403274 28350
rect 403342 28294 403398 28350
rect 402970 28170 403026 28226
rect 403094 28170 403150 28226
rect 403218 28170 403274 28226
rect 403342 28170 403398 28226
rect 402970 28046 403026 28102
rect 403094 28046 403150 28102
rect 403218 28046 403274 28102
rect 403342 28046 403398 28102
rect 402970 27922 403026 27978
rect 403094 27922 403150 27978
rect 403218 27922 403274 27978
rect 403342 27922 403398 27978
rect 402970 10294 403026 10350
rect 403094 10294 403150 10350
rect 403218 10294 403274 10350
rect 403342 10294 403398 10350
rect 402970 10170 403026 10226
rect 403094 10170 403150 10226
rect 403218 10170 403274 10226
rect 403342 10170 403398 10226
rect 402970 10046 403026 10102
rect 403094 10046 403150 10102
rect 403218 10046 403274 10102
rect 403342 10046 403398 10102
rect 402970 9922 403026 9978
rect 403094 9922 403150 9978
rect 403218 9922 403274 9978
rect 403342 9922 403398 9978
rect 402970 -1176 403026 -1120
rect 403094 -1176 403150 -1120
rect 403218 -1176 403274 -1120
rect 403342 -1176 403398 -1120
rect 402970 -1300 403026 -1244
rect 403094 -1300 403150 -1244
rect 403218 -1300 403274 -1244
rect 403342 -1300 403398 -1244
rect 402970 -1424 403026 -1368
rect 403094 -1424 403150 -1368
rect 403218 -1424 403274 -1368
rect 403342 -1424 403398 -1368
rect 402970 -1548 403026 -1492
rect 403094 -1548 403150 -1492
rect 403218 -1548 403274 -1492
rect 403342 -1548 403398 -1492
rect 417250 148294 417306 148350
rect 417374 148294 417430 148350
rect 417498 148294 417554 148350
rect 417622 148294 417678 148350
rect 417250 148170 417306 148226
rect 417374 148170 417430 148226
rect 417498 148170 417554 148226
rect 417622 148170 417678 148226
rect 417250 148046 417306 148102
rect 417374 148046 417430 148102
rect 417498 148046 417554 148102
rect 417622 148046 417678 148102
rect 417250 147922 417306 147978
rect 417374 147922 417430 147978
rect 417498 147922 417554 147978
rect 417622 147922 417678 147978
rect 417250 130294 417306 130350
rect 417374 130294 417430 130350
rect 417498 130294 417554 130350
rect 417622 130294 417678 130350
rect 417250 130170 417306 130226
rect 417374 130170 417430 130226
rect 417498 130170 417554 130226
rect 417622 130170 417678 130226
rect 417250 130046 417306 130102
rect 417374 130046 417430 130102
rect 417498 130046 417554 130102
rect 417622 130046 417678 130102
rect 417250 129922 417306 129978
rect 417374 129922 417430 129978
rect 417498 129922 417554 129978
rect 417622 129922 417678 129978
rect 417250 112294 417306 112350
rect 417374 112294 417430 112350
rect 417498 112294 417554 112350
rect 417622 112294 417678 112350
rect 417250 112170 417306 112226
rect 417374 112170 417430 112226
rect 417498 112170 417554 112226
rect 417622 112170 417678 112226
rect 417250 112046 417306 112102
rect 417374 112046 417430 112102
rect 417498 112046 417554 112102
rect 417622 112046 417678 112102
rect 417250 111922 417306 111978
rect 417374 111922 417430 111978
rect 417498 111922 417554 111978
rect 417622 111922 417678 111978
rect 417250 94294 417306 94350
rect 417374 94294 417430 94350
rect 417498 94294 417554 94350
rect 417622 94294 417678 94350
rect 417250 94170 417306 94226
rect 417374 94170 417430 94226
rect 417498 94170 417554 94226
rect 417622 94170 417678 94226
rect 417250 94046 417306 94102
rect 417374 94046 417430 94102
rect 417498 94046 417554 94102
rect 417622 94046 417678 94102
rect 417250 93922 417306 93978
rect 417374 93922 417430 93978
rect 417498 93922 417554 93978
rect 417622 93922 417678 93978
rect 417250 76294 417306 76350
rect 417374 76294 417430 76350
rect 417498 76294 417554 76350
rect 417622 76294 417678 76350
rect 417250 76170 417306 76226
rect 417374 76170 417430 76226
rect 417498 76170 417554 76226
rect 417622 76170 417678 76226
rect 417250 76046 417306 76102
rect 417374 76046 417430 76102
rect 417498 76046 417554 76102
rect 417622 76046 417678 76102
rect 417250 75922 417306 75978
rect 417374 75922 417430 75978
rect 417498 75922 417554 75978
rect 417622 75922 417678 75978
rect 417250 58294 417306 58350
rect 417374 58294 417430 58350
rect 417498 58294 417554 58350
rect 417622 58294 417678 58350
rect 417250 58170 417306 58226
rect 417374 58170 417430 58226
rect 417498 58170 417554 58226
rect 417622 58170 417678 58226
rect 417250 58046 417306 58102
rect 417374 58046 417430 58102
rect 417498 58046 417554 58102
rect 417622 58046 417678 58102
rect 417250 57922 417306 57978
rect 417374 57922 417430 57978
rect 417498 57922 417554 57978
rect 417622 57922 417678 57978
rect 417250 40294 417306 40350
rect 417374 40294 417430 40350
rect 417498 40294 417554 40350
rect 417622 40294 417678 40350
rect 417250 40170 417306 40226
rect 417374 40170 417430 40226
rect 417498 40170 417554 40226
rect 417622 40170 417678 40226
rect 417250 40046 417306 40102
rect 417374 40046 417430 40102
rect 417498 40046 417554 40102
rect 417622 40046 417678 40102
rect 417250 39922 417306 39978
rect 417374 39922 417430 39978
rect 417498 39922 417554 39978
rect 417622 39922 417678 39978
rect 417250 22294 417306 22350
rect 417374 22294 417430 22350
rect 417498 22294 417554 22350
rect 417622 22294 417678 22350
rect 417250 22170 417306 22226
rect 417374 22170 417430 22226
rect 417498 22170 417554 22226
rect 417622 22170 417678 22226
rect 417250 22046 417306 22102
rect 417374 22046 417430 22102
rect 417498 22046 417554 22102
rect 417622 22046 417678 22102
rect 417250 21922 417306 21978
rect 417374 21922 417430 21978
rect 417498 21922 417554 21978
rect 417622 21922 417678 21978
rect 417250 4294 417306 4350
rect 417374 4294 417430 4350
rect 417498 4294 417554 4350
rect 417622 4294 417678 4350
rect 417250 4170 417306 4226
rect 417374 4170 417430 4226
rect 417498 4170 417554 4226
rect 417622 4170 417678 4226
rect 417250 4046 417306 4102
rect 417374 4046 417430 4102
rect 417498 4046 417554 4102
rect 417622 4046 417678 4102
rect 417250 3922 417306 3978
rect 417374 3922 417430 3978
rect 417498 3922 417554 3978
rect 417622 3922 417678 3978
rect 417250 -216 417306 -160
rect 417374 -216 417430 -160
rect 417498 -216 417554 -160
rect 417622 -216 417678 -160
rect 417250 -340 417306 -284
rect 417374 -340 417430 -284
rect 417498 -340 417554 -284
rect 417622 -340 417678 -284
rect 417250 -464 417306 -408
rect 417374 -464 417430 -408
rect 417498 -464 417554 -408
rect 417622 -464 417678 -408
rect 417250 -588 417306 -532
rect 417374 -588 417430 -532
rect 417498 -588 417554 -532
rect 417622 -588 417678 -532
rect 420970 154294 421026 154350
rect 421094 154294 421150 154350
rect 421218 154294 421274 154350
rect 421342 154294 421398 154350
rect 420970 154170 421026 154226
rect 421094 154170 421150 154226
rect 421218 154170 421274 154226
rect 421342 154170 421398 154226
rect 420970 154046 421026 154102
rect 421094 154046 421150 154102
rect 421218 154046 421274 154102
rect 421342 154046 421398 154102
rect 420970 153922 421026 153978
rect 421094 153922 421150 153978
rect 421218 153922 421274 153978
rect 421342 153922 421398 153978
rect 420970 136294 421026 136350
rect 421094 136294 421150 136350
rect 421218 136294 421274 136350
rect 421342 136294 421398 136350
rect 420970 136170 421026 136226
rect 421094 136170 421150 136226
rect 421218 136170 421274 136226
rect 421342 136170 421398 136226
rect 420970 136046 421026 136102
rect 421094 136046 421150 136102
rect 421218 136046 421274 136102
rect 421342 136046 421398 136102
rect 420970 135922 421026 135978
rect 421094 135922 421150 135978
rect 421218 135922 421274 135978
rect 421342 135922 421398 135978
rect 420970 118294 421026 118350
rect 421094 118294 421150 118350
rect 421218 118294 421274 118350
rect 421342 118294 421398 118350
rect 420970 118170 421026 118226
rect 421094 118170 421150 118226
rect 421218 118170 421274 118226
rect 421342 118170 421398 118226
rect 420970 118046 421026 118102
rect 421094 118046 421150 118102
rect 421218 118046 421274 118102
rect 421342 118046 421398 118102
rect 420970 117922 421026 117978
rect 421094 117922 421150 117978
rect 421218 117922 421274 117978
rect 421342 117922 421398 117978
rect 420970 100294 421026 100350
rect 421094 100294 421150 100350
rect 421218 100294 421274 100350
rect 421342 100294 421398 100350
rect 420970 100170 421026 100226
rect 421094 100170 421150 100226
rect 421218 100170 421274 100226
rect 421342 100170 421398 100226
rect 420970 100046 421026 100102
rect 421094 100046 421150 100102
rect 421218 100046 421274 100102
rect 421342 100046 421398 100102
rect 420970 99922 421026 99978
rect 421094 99922 421150 99978
rect 421218 99922 421274 99978
rect 421342 99922 421398 99978
rect 420970 82294 421026 82350
rect 421094 82294 421150 82350
rect 421218 82294 421274 82350
rect 421342 82294 421398 82350
rect 420970 82170 421026 82226
rect 421094 82170 421150 82226
rect 421218 82170 421274 82226
rect 421342 82170 421398 82226
rect 420970 82046 421026 82102
rect 421094 82046 421150 82102
rect 421218 82046 421274 82102
rect 421342 82046 421398 82102
rect 420970 81922 421026 81978
rect 421094 81922 421150 81978
rect 421218 81922 421274 81978
rect 421342 81922 421398 81978
rect 420970 64294 421026 64350
rect 421094 64294 421150 64350
rect 421218 64294 421274 64350
rect 421342 64294 421398 64350
rect 420970 64170 421026 64226
rect 421094 64170 421150 64226
rect 421218 64170 421274 64226
rect 421342 64170 421398 64226
rect 420970 64046 421026 64102
rect 421094 64046 421150 64102
rect 421218 64046 421274 64102
rect 421342 64046 421398 64102
rect 420970 63922 421026 63978
rect 421094 63922 421150 63978
rect 421218 63922 421274 63978
rect 421342 63922 421398 63978
rect 420970 46294 421026 46350
rect 421094 46294 421150 46350
rect 421218 46294 421274 46350
rect 421342 46294 421398 46350
rect 420970 46170 421026 46226
rect 421094 46170 421150 46226
rect 421218 46170 421274 46226
rect 421342 46170 421398 46226
rect 420970 46046 421026 46102
rect 421094 46046 421150 46102
rect 421218 46046 421274 46102
rect 421342 46046 421398 46102
rect 420970 45922 421026 45978
rect 421094 45922 421150 45978
rect 421218 45922 421274 45978
rect 421342 45922 421398 45978
rect 420970 28294 421026 28350
rect 421094 28294 421150 28350
rect 421218 28294 421274 28350
rect 421342 28294 421398 28350
rect 420970 28170 421026 28226
rect 421094 28170 421150 28226
rect 421218 28170 421274 28226
rect 421342 28170 421398 28226
rect 420970 28046 421026 28102
rect 421094 28046 421150 28102
rect 421218 28046 421274 28102
rect 421342 28046 421398 28102
rect 420970 27922 421026 27978
rect 421094 27922 421150 27978
rect 421218 27922 421274 27978
rect 421342 27922 421398 27978
rect 420970 10294 421026 10350
rect 421094 10294 421150 10350
rect 421218 10294 421274 10350
rect 421342 10294 421398 10350
rect 420970 10170 421026 10226
rect 421094 10170 421150 10226
rect 421218 10170 421274 10226
rect 421342 10170 421398 10226
rect 420970 10046 421026 10102
rect 421094 10046 421150 10102
rect 421218 10046 421274 10102
rect 421342 10046 421398 10102
rect 420970 9922 421026 9978
rect 421094 9922 421150 9978
rect 421218 9922 421274 9978
rect 421342 9922 421398 9978
rect 420970 -1176 421026 -1120
rect 421094 -1176 421150 -1120
rect 421218 -1176 421274 -1120
rect 421342 -1176 421398 -1120
rect 420970 -1300 421026 -1244
rect 421094 -1300 421150 -1244
rect 421218 -1300 421274 -1244
rect 421342 -1300 421398 -1244
rect 420970 -1424 421026 -1368
rect 421094 -1424 421150 -1368
rect 421218 -1424 421274 -1368
rect 421342 -1424 421398 -1368
rect 420970 -1548 421026 -1492
rect 421094 -1548 421150 -1492
rect 421218 -1548 421274 -1492
rect 421342 -1548 421398 -1492
rect 435250 148294 435306 148350
rect 435374 148294 435430 148350
rect 435498 148294 435554 148350
rect 435622 148294 435678 148350
rect 435250 148170 435306 148226
rect 435374 148170 435430 148226
rect 435498 148170 435554 148226
rect 435622 148170 435678 148226
rect 435250 148046 435306 148102
rect 435374 148046 435430 148102
rect 435498 148046 435554 148102
rect 435622 148046 435678 148102
rect 435250 147922 435306 147978
rect 435374 147922 435430 147978
rect 435498 147922 435554 147978
rect 435622 147922 435678 147978
rect 435250 130294 435306 130350
rect 435374 130294 435430 130350
rect 435498 130294 435554 130350
rect 435622 130294 435678 130350
rect 435250 130170 435306 130226
rect 435374 130170 435430 130226
rect 435498 130170 435554 130226
rect 435622 130170 435678 130226
rect 435250 130046 435306 130102
rect 435374 130046 435430 130102
rect 435498 130046 435554 130102
rect 435622 130046 435678 130102
rect 435250 129922 435306 129978
rect 435374 129922 435430 129978
rect 435498 129922 435554 129978
rect 435622 129922 435678 129978
rect 435250 112294 435306 112350
rect 435374 112294 435430 112350
rect 435498 112294 435554 112350
rect 435622 112294 435678 112350
rect 435250 112170 435306 112226
rect 435374 112170 435430 112226
rect 435498 112170 435554 112226
rect 435622 112170 435678 112226
rect 435250 112046 435306 112102
rect 435374 112046 435430 112102
rect 435498 112046 435554 112102
rect 435622 112046 435678 112102
rect 435250 111922 435306 111978
rect 435374 111922 435430 111978
rect 435498 111922 435554 111978
rect 435622 111922 435678 111978
rect 435250 94294 435306 94350
rect 435374 94294 435430 94350
rect 435498 94294 435554 94350
rect 435622 94294 435678 94350
rect 435250 94170 435306 94226
rect 435374 94170 435430 94226
rect 435498 94170 435554 94226
rect 435622 94170 435678 94226
rect 435250 94046 435306 94102
rect 435374 94046 435430 94102
rect 435498 94046 435554 94102
rect 435622 94046 435678 94102
rect 435250 93922 435306 93978
rect 435374 93922 435430 93978
rect 435498 93922 435554 93978
rect 435622 93922 435678 93978
rect 435250 76294 435306 76350
rect 435374 76294 435430 76350
rect 435498 76294 435554 76350
rect 435622 76294 435678 76350
rect 435250 76170 435306 76226
rect 435374 76170 435430 76226
rect 435498 76170 435554 76226
rect 435622 76170 435678 76226
rect 435250 76046 435306 76102
rect 435374 76046 435430 76102
rect 435498 76046 435554 76102
rect 435622 76046 435678 76102
rect 435250 75922 435306 75978
rect 435374 75922 435430 75978
rect 435498 75922 435554 75978
rect 435622 75922 435678 75978
rect 435250 58294 435306 58350
rect 435374 58294 435430 58350
rect 435498 58294 435554 58350
rect 435622 58294 435678 58350
rect 435250 58170 435306 58226
rect 435374 58170 435430 58226
rect 435498 58170 435554 58226
rect 435622 58170 435678 58226
rect 435250 58046 435306 58102
rect 435374 58046 435430 58102
rect 435498 58046 435554 58102
rect 435622 58046 435678 58102
rect 435250 57922 435306 57978
rect 435374 57922 435430 57978
rect 435498 57922 435554 57978
rect 435622 57922 435678 57978
rect 435250 40294 435306 40350
rect 435374 40294 435430 40350
rect 435498 40294 435554 40350
rect 435622 40294 435678 40350
rect 435250 40170 435306 40226
rect 435374 40170 435430 40226
rect 435498 40170 435554 40226
rect 435622 40170 435678 40226
rect 435250 40046 435306 40102
rect 435374 40046 435430 40102
rect 435498 40046 435554 40102
rect 435622 40046 435678 40102
rect 435250 39922 435306 39978
rect 435374 39922 435430 39978
rect 435498 39922 435554 39978
rect 435622 39922 435678 39978
rect 435250 22294 435306 22350
rect 435374 22294 435430 22350
rect 435498 22294 435554 22350
rect 435622 22294 435678 22350
rect 435250 22170 435306 22226
rect 435374 22170 435430 22226
rect 435498 22170 435554 22226
rect 435622 22170 435678 22226
rect 435250 22046 435306 22102
rect 435374 22046 435430 22102
rect 435498 22046 435554 22102
rect 435622 22046 435678 22102
rect 435250 21922 435306 21978
rect 435374 21922 435430 21978
rect 435498 21922 435554 21978
rect 435622 21922 435678 21978
rect 435250 4294 435306 4350
rect 435374 4294 435430 4350
rect 435498 4294 435554 4350
rect 435622 4294 435678 4350
rect 435250 4170 435306 4226
rect 435374 4170 435430 4226
rect 435498 4170 435554 4226
rect 435622 4170 435678 4226
rect 435250 4046 435306 4102
rect 435374 4046 435430 4102
rect 435498 4046 435554 4102
rect 435622 4046 435678 4102
rect 435250 3922 435306 3978
rect 435374 3922 435430 3978
rect 435498 3922 435554 3978
rect 435622 3922 435678 3978
rect 435250 -216 435306 -160
rect 435374 -216 435430 -160
rect 435498 -216 435554 -160
rect 435622 -216 435678 -160
rect 435250 -340 435306 -284
rect 435374 -340 435430 -284
rect 435498 -340 435554 -284
rect 435622 -340 435678 -284
rect 435250 -464 435306 -408
rect 435374 -464 435430 -408
rect 435498 -464 435554 -408
rect 435622 -464 435678 -408
rect 435250 -588 435306 -532
rect 435374 -588 435430 -532
rect 435498 -588 435554 -532
rect 435622 -588 435678 -532
rect 438970 154294 439026 154350
rect 439094 154294 439150 154350
rect 439218 154294 439274 154350
rect 439342 154294 439398 154350
rect 438970 154170 439026 154226
rect 439094 154170 439150 154226
rect 439218 154170 439274 154226
rect 439342 154170 439398 154226
rect 438970 154046 439026 154102
rect 439094 154046 439150 154102
rect 439218 154046 439274 154102
rect 439342 154046 439398 154102
rect 438970 153922 439026 153978
rect 439094 153922 439150 153978
rect 439218 153922 439274 153978
rect 439342 153922 439398 153978
rect 438970 136294 439026 136350
rect 439094 136294 439150 136350
rect 439218 136294 439274 136350
rect 439342 136294 439398 136350
rect 438970 136170 439026 136226
rect 439094 136170 439150 136226
rect 439218 136170 439274 136226
rect 439342 136170 439398 136226
rect 438970 136046 439026 136102
rect 439094 136046 439150 136102
rect 439218 136046 439274 136102
rect 439342 136046 439398 136102
rect 438970 135922 439026 135978
rect 439094 135922 439150 135978
rect 439218 135922 439274 135978
rect 439342 135922 439398 135978
rect 438970 118294 439026 118350
rect 439094 118294 439150 118350
rect 439218 118294 439274 118350
rect 439342 118294 439398 118350
rect 438970 118170 439026 118226
rect 439094 118170 439150 118226
rect 439218 118170 439274 118226
rect 439342 118170 439398 118226
rect 438970 118046 439026 118102
rect 439094 118046 439150 118102
rect 439218 118046 439274 118102
rect 439342 118046 439398 118102
rect 438970 117922 439026 117978
rect 439094 117922 439150 117978
rect 439218 117922 439274 117978
rect 439342 117922 439398 117978
rect 438970 100294 439026 100350
rect 439094 100294 439150 100350
rect 439218 100294 439274 100350
rect 439342 100294 439398 100350
rect 438970 100170 439026 100226
rect 439094 100170 439150 100226
rect 439218 100170 439274 100226
rect 439342 100170 439398 100226
rect 438970 100046 439026 100102
rect 439094 100046 439150 100102
rect 439218 100046 439274 100102
rect 439342 100046 439398 100102
rect 438970 99922 439026 99978
rect 439094 99922 439150 99978
rect 439218 99922 439274 99978
rect 439342 99922 439398 99978
rect 438970 82294 439026 82350
rect 439094 82294 439150 82350
rect 439218 82294 439274 82350
rect 439342 82294 439398 82350
rect 438970 82170 439026 82226
rect 439094 82170 439150 82226
rect 439218 82170 439274 82226
rect 439342 82170 439398 82226
rect 438970 82046 439026 82102
rect 439094 82046 439150 82102
rect 439218 82046 439274 82102
rect 439342 82046 439398 82102
rect 438970 81922 439026 81978
rect 439094 81922 439150 81978
rect 439218 81922 439274 81978
rect 439342 81922 439398 81978
rect 438970 64294 439026 64350
rect 439094 64294 439150 64350
rect 439218 64294 439274 64350
rect 439342 64294 439398 64350
rect 438970 64170 439026 64226
rect 439094 64170 439150 64226
rect 439218 64170 439274 64226
rect 439342 64170 439398 64226
rect 438970 64046 439026 64102
rect 439094 64046 439150 64102
rect 439218 64046 439274 64102
rect 439342 64046 439398 64102
rect 438970 63922 439026 63978
rect 439094 63922 439150 63978
rect 439218 63922 439274 63978
rect 439342 63922 439398 63978
rect 438970 46294 439026 46350
rect 439094 46294 439150 46350
rect 439218 46294 439274 46350
rect 439342 46294 439398 46350
rect 438970 46170 439026 46226
rect 439094 46170 439150 46226
rect 439218 46170 439274 46226
rect 439342 46170 439398 46226
rect 438970 46046 439026 46102
rect 439094 46046 439150 46102
rect 439218 46046 439274 46102
rect 439342 46046 439398 46102
rect 438970 45922 439026 45978
rect 439094 45922 439150 45978
rect 439218 45922 439274 45978
rect 439342 45922 439398 45978
rect 438970 28294 439026 28350
rect 439094 28294 439150 28350
rect 439218 28294 439274 28350
rect 439342 28294 439398 28350
rect 438970 28170 439026 28226
rect 439094 28170 439150 28226
rect 439218 28170 439274 28226
rect 439342 28170 439398 28226
rect 438970 28046 439026 28102
rect 439094 28046 439150 28102
rect 439218 28046 439274 28102
rect 439342 28046 439398 28102
rect 438970 27922 439026 27978
rect 439094 27922 439150 27978
rect 439218 27922 439274 27978
rect 439342 27922 439398 27978
rect 438970 10294 439026 10350
rect 439094 10294 439150 10350
rect 439218 10294 439274 10350
rect 439342 10294 439398 10350
rect 438970 10170 439026 10226
rect 439094 10170 439150 10226
rect 439218 10170 439274 10226
rect 439342 10170 439398 10226
rect 438970 10046 439026 10102
rect 439094 10046 439150 10102
rect 439218 10046 439274 10102
rect 439342 10046 439398 10102
rect 438970 9922 439026 9978
rect 439094 9922 439150 9978
rect 439218 9922 439274 9978
rect 439342 9922 439398 9978
rect 438970 -1176 439026 -1120
rect 439094 -1176 439150 -1120
rect 439218 -1176 439274 -1120
rect 439342 -1176 439398 -1120
rect 438970 -1300 439026 -1244
rect 439094 -1300 439150 -1244
rect 439218 -1300 439274 -1244
rect 439342 -1300 439398 -1244
rect 438970 -1424 439026 -1368
rect 439094 -1424 439150 -1368
rect 439218 -1424 439274 -1368
rect 439342 -1424 439398 -1368
rect 438970 -1548 439026 -1492
rect 439094 -1548 439150 -1492
rect 439218 -1548 439274 -1492
rect 439342 -1548 439398 -1492
rect 453250 148294 453306 148350
rect 453374 148294 453430 148350
rect 453498 148294 453554 148350
rect 453622 148294 453678 148350
rect 453250 148170 453306 148226
rect 453374 148170 453430 148226
rect 453498 148170 453554 148226
rect 453622 148170 453678 148226
rect 453250 148046 453306 148102
rect 453374 148046 453430 148102
rect 453498 148046 453554 148102
rect 453622 148046 453678 148102
rect 453250 147922 453306 147978
rect 453374 147922 453430 147978
rect 453498 147922 453554 147978
rect 453622 147922 453678 147978
rect 453250 130294 453306 130350
rect 453374 130294 453430 130350
rect 453498 130294 453554 130350
rect 453622 130294 453678 130350
rect 453250 130170 453306 130226
rect 453374 130170 453430 130226
rect 453498 130170 453554 130226
rect 453622 130170 453678 130226
rect 453250 130046 453306 130102
rect 453374 130046 453430 130102
rect 453498 130046 453554 130102
rect 453622 130046 453678 130102
rect 453250 129922 453306 129978
rect 453374 129922 453430 129978
rect 453498 129922 453554 129978
rect 453622 129922 453678 129978
rect 453250 112294 453306 112350
rect 453374 112294 453430 112350
rect 453498 112294 453554 112350
rect 453622 112294 453678 112350
rect 453250 112170 453306 112226
rect 453374 112170 453430 112226
rect 453498 112170 453554 112226
rect 453622 112170 453678 112226
rect 453250 112046 453306 112102
rect 453374 112046 453430 112102
rect 453498 112046 453554 112102
rect 453622 112046 453678 112102
rect 453250 111922 453306 111978
rect 453374 111922 453430 111978
rect 453498 111922 453554 111978
rect 453622 111922 453678 111978
rect 453250 94294 453306 94350
rect 453374 94294 453430 94350
rect 453498 94294 453554 94350
rect 453622 94294 453678 94350
rect 453250 94170 453306 94226
rect 453374 94170 453430 94226
rect 453498 94170 453554 94226
rect 453622 94170 453678 94226
rect 453250 94046 453306 94102
rect 453374 94046 453430 94102
rect 453498 94046 453554 94102
rect 453622 94046 453678 94102
rect 453250 93922 453306 93978
rect 453374 93922 453430 93978
rect 453498 93922 453554 93978
rect 453622 93922 453678 93978
rect 453250 76294 453306 76350
rect 453374 76294 453430 76350
rect 453498 76294 453554 76350
rect 453622 76294 453678 76350
rect 453250 76170 453306 76226
rect 453374 76170 453430 76226
rect 453498 76170 453554 76226
rect 453622 76170 453678 76226
rect 453250 76046 453306 76102
rect 453374 76046 453430 76102
rect 453498 76046 453554 76102
rect 453622 76046 453678 76102
rect 453250 75922 453306 75978
rect 453374 75922 453430 75978
rect 453498 75922 453554 75978
rect 453622 75922 453678 75978
rect 453250 58294 453306 58350
rect 453374 58294 453430 58350
rect 453498 58294 453554 58350
rect 453622 58294 453678 58350
rect 453250 58170 453306 58226
rect 453374 58170 453430 58226
rect 453498 58170 453554 58226
rect 453622 58170 453678 58226
rect 453250 58046 453306 58102
rect 453374 58046 453430 58102
rect 453498 58046 453554 58102
rect 453622 58046 453678 58102
rect 453250 57922 453306 57978
rect 453374 57922 453430 57978
rect 453498 57922 453554 57978
rect 453622 57922 453678 57978
rect 453250 40294 453306 40350
rect 453374 40294 453430 40350
rect 453498 40294 453554 40350
rect 453622 40294 453678 40350
rect 453250 40170 453306 40226
rect 453374 40170 453430 40226
rect 453498 40170 453554 40226
rect 453622 40170 453678 40226
rect 453250 40046 453306 40102
rect 453374 40046 453430 40102
rect 453498 40046 453554 40102
rect 453622 40046 453678 40102
rect 453250 39922 453306 39978
rect 453374 39922 453430 39978
rect 453498 39922 453554 39978
rect 453622 39922 453678 39978
rect 453250 22294 453306 22350
rect 453374 22294 453430 22350
rect 453498 22294 453554 22350
rect 453622 22294 453678 22350
rect 453250 22170 453306 22226
rect 453374 22170 453430 22226
rect 453498 22170 453554 22226
rect 453622 22170 453678 22226
rect 453250 22046 453306 22102
rect 453374 22046 453430 22102
rect 453498 22046 453554 22102
rect 453622 22046 453678 22102
rect 453250 21922 453306 21978
rect 453374 21922 453430 21978
rect 453498 21922 453554 21978
rect 453622 21922 453678 21978
rect 453250 4294 453306 4350
rect 453374 4294 453430 4350
rect 453498 4294 453554 4350
rect 453622 4294 453678 4350
rect 453250 4170 453306 4226
rect 453374 4170 453430 4226
rect 453498 4170 453554 4226
rect 453622 4170 453678 4226
rect 453250 4046 453306 4102
rect 453374 4046 453430 4102
rect 453498 4046 453554 4102
rect 453622 4046 453678 4102
rect 453250 3922 453306 3978
rect 453374 3922 453430 3978
rect 453498 3922 453554 3978
rect 453622 3922 453678 3978
rect 453250 -216 453306 -160
rect 453374 -216 453430 -160
rect 453498 -216 453554 -160
rect 453622 -216 453678 -160
rect 453250 -340 453306 -284
rect 453374 -340 453430 -284
rect 453498 -340 453554 -284
rect 453622 -340 453678 -284
rect 453250 -464 453306 -408
rect 453374 -464 453430 -408
rect 453498 -464 453554 -408
rect 453622 -464 453678 -408
rect 453250 -588 453306 -532
rect 453374 -588 453430 -532
rect 453498 -588 453554 -532
rect 453622 -588 453678 -532
rect 456970 154294 457026 154350
rect 457094 154294 457150 154350
rect 457218 154294 457274 154350
rect 457342 154294 457398 154350
rect 456970 154170 457026 154226
rect 457094 154170 457150 154226
rect 457218 154170 457274 154226
rect 457342 154170 457398 154226
rect 456970 154046 457026 154102
rect 457094 154046 457150 154102
rect 457218 154046 457274 154102
rect 457342 154046 457398 154102
rect 456970 153922 457026 153978
rect 457094 153922 457150 153978
rect 457218 153922 457274 153978
rect 457342 153922 457398 153978
rect 456970 136294 457026 136350
rect 457094 136294 457150 136350
rect 457218 136294 457274 136350
rect 457342 136294 457398 136350
rect 456970 136170 457026 136226
rect 457094 136170 457150 136226
rect 457218 136170 457274 136226
rect 457342 136170 457398 136226
rect 456970 136046 457026 136102
rect 457094 136046 457150 136102
rect 457218 136046 457274 136102
rect 457342 136046 457398 136102
rect 456970 135922 457026 135978
rect 457094 135922 457150 135978
rect 457218 135922 457274 135978
rect 457342 135922 457398 135978
rect 456970 118294 457026 118350
rect 457094 118294 457150 118350
rect 457218 118294 457274 118350
rect 457342 118294 457398 118350
rect 456970 118170 457026 118226
rect 457094 118170 457150 118226
rect 457218 118170 457274 118226
rect 457342 118170 457398 118226
rect 456970 118046 457026 118102
rect 457094 118046 457150 118102
rect 457218 118046 457274 118102
rect 457342 118046 457398 118102
rect 456970 117922 457026 117978
rect 457094 117922 457150 117978
rect 457218 117922 457274 117978
rect 457342 117922 457398 117978
rect 456970 100294 457026 100350
rect 457094 100294 457150 100350
rect 457218 100294 457274 100350
rect 457342 100294 457398 100350
rect 456970 100170 457026 100226
rect 457094 100170 457150 100226
rect 457218 100170 457274 100226
rect 457342 100170 457398 100226
rect 456970 100046 457026 100102
rect 457094 100046 457150 100102
rect 457218 100046 457274 100102
rect 457342 100046 457398 100102
rect 456970 99922 457026 99978
rect 457094 99922 457150 99978
rect 457218 99922 457274 99978
rect 457342 99922 457398 99978
rect 456970 82294 457026 82350
rect 457094 82294 457150 82350
rect 457218 82294 457274 82350
rect 457342 82294 457398 82350
rect 456970 82170 457026 82226
rect 457094 82170 457150 82226
rect 457218 82170 457274 82226
rect 457342 82170 457398 82226
rect 456970 82046 457026 82102
rect 457094 82046 457150 82102
rect 457218 82046 457274 82102
rect 457342 82046 457398 82102
rect 456970 81922 457026 81978
rect 457094 81922 457150 81978
rect 457218 81922 457274 81978
rect 457342 81922 457398 81978
rect 456970 64294 457026 64350
rect 457094 64294 457150 64350
rect 457218 64294 457274 64350
rect 457342 64294 457398 64350
rect 456970 64170 457026 64226
rect 457094 64170 457150 64226
rect 457218 64170 457274 64226
rect 457342 64170 457398 64226
rect 456970 64046 457026 64102
rect 457094 64046 457150 64102
rect 457218 64046 457274 64102
rect 457342 64046 457398 64102
rect 456970 63922 457026 63978
rect 457094 63922 457150 63978
rect 457218 63922 457274 63978
rect 457342 63922 457398 63978
rect 456970 46294 457026 46350
rect 457094 46294 457150 46350
rect 457218 46294 457274 46350
rect 457342 46294 457398 46350
rect 456970 46170 457026 46226
rect 457094 46170 457150 46226
rect 457218 46170 457274 46226
rect 457342 46170 457398 46226
rect 456970 46046 457026 46102
rect 457094 46046 457150 46102
rect 457218 46046 457274 46102
rect 457342 46046 457398 46102
rect 456970 45922 457026 45978
rect 457094 45922 457150 45978
rect 457218 45922 457274 45978
rect 457342 45922 457398 45978
rect 456970 28294 457026 28350
rect 457094 28294 457150 28350
rect 457218 28294 457274 28350
rect 457342 28294 457398 28350
rect 456970 28170 457026 28226
rect 457094 28170 457150 28226
rect 457218 28170 457274 28226
rect 457342 28170 457398 28226
rect 456970 28046 457026 28102
rect 457094 28046 457150 28102
rect 457218 28046 457274 28102
rect 457342 28046 457398 28102
rect 456970 27922 457026 27978
rect 457094 27922 457150 27978
rect 457218 27922 457274 27978
rect 457342 27922 457398 27978
rect 456970 10294 457026 10350
rect 457094 10294 457150 10350
rect 457218 10294 457274 10350
rect 457342 10294 457398 10350
rect 456970 10170 457026 10226
rect 457094 10170 457150 10226
rect 457218 10170 457274 10226
rect 457342 10170 457398 10226
rect 456970 10046 457026 10102
rect 457094 10046 457150 10102
rect 457218 10046 457274 10102
rect 457342 10046 457398 10102
rect 456970 9922 457026 9978
rect 457094 9922 457150 9978
rect 457218 9922 457274 9978
rect 457342 9922 457398 9978
rect 456970 -1176 457026 -1120
rect 457094 -1176 457150 -1120
rect 457218 -1176 457274 -1120
rect 457342 -1176 457398 -1120
rect 456970 -1300 457026 -1244
rect 457094 -1300 457150 -1244
rect 457218 -1300 457274 -1244
rect 457342 -1300 457398 -1244
rect 456970 -1424 457026 -1368
rect 457094 -1424 457150 -1368
rect 457218 -1424 457274 -1368
rect 457342 -1424 457398 -1368
rect 456970 -1548 457026 -1492
rect 457094 -1548 457150 -1492
rect 457218 -1548 457274 -1492
rect 457342 -1548 457398 -1492
rect 471250 148294 471306 148350
rect 471374 148294 471430 148350
rect 471498 148294 471554 148350
rect 471622 148294 471678 148350
rect 471250 148170 471306 148226
rect 471374 148170 471430 148226
rect 471498 148170 471554 148226
rect 471622 148170 471678 148226
rect 471250 148046 471306 148102
rect 471374 148046 471430 148102
rect 471498 148046 471554 148102
rect 471622 148046 471678 148102
rect 471250 147922 471306 147978
rect 471374 147922 471430 147978
rect 471498 147922 471554 147978
rect 471622 147922 471678 147978
rect 471250 130294 471306 130350
rect 471374 130294 471430 130350
rect 471498 130294 471554 130350
rect 471622 130294 471678 130350
rect 471250 130170 471306 130226
rect 471374 130170 471430 130226
rect 471498 130170 471554 130226
rect 471622 130170 471678 130226
rect 471250 130046 471306 130102
rect 471374 130046 471430 130102
rect 471498 130046 471554 130102
rect 471622 130046 471678 130102
rect 471250 129922 471306 129978
rect 471374 129922 471430 129978
rect 471498 129922 471554 129978
rect 471622 129922 471678 129978
rect 471250 112294 471306 112350
rect 471374 112294 471430 112350
rect 471498 112294 471554 112350
rect 471622 112294 471678 112350
rect 471250 112170 471306 112226
rect 471374 112170 471430 112226
rect 471498 112170 471554 112226
rect 471622 112170 471678 112226
rect 471250 112046 471306 112102
rect 471374 112046 471430 112102
rect 471498 112046 471554 112102
rect 471622 112046 471678 112102
rect 471250 111922 471306 111978
rect 471374 111922 471430 111978
rect 471498 111922 471554 111978
rect 471622 111922 471678 111978
rect 471250 94294 471306 94350
rect 471374 94294 471430 94350
rect 471498 94294 471554 94350
rect 471622 94294 471678 94350
rect 471250 94170 471306 94226
rect 471374 94170 471430 94226
rect 471498 94170 471554 94226
rect 471622 94170 471678 94226
rect 471250 94046 471306 94102
rect 471374 94046 471430 94102
rect 471498 94046 471554 94102
rect 471622 94046 471678 94102
rect 471250 93922 471306 93978
rect 471374 93922 471430 93978
rect 471498 93922 471554 93978
rect 471622 93922 471678 93978
rect 471250 76294 471306 76350
rect 471374 76294 471430 76350
rect 471498 76294 471554 76350
rect 471622 76294 471678 76350
rect 471250 76170 471306 76226
rect 471374 76170 471430 76226
rect 471498 76170 471554 76226
rect 471622 76170 471678 76226
rect 471250 76046 471306 76102
rect 471374 76046 471430 76102
rect 471498 76046 471554 76102
rect 471622 76046 471678 76102
rect 471250 75922 471306 75978
rect 471374 75922 471430 75978
rect 471498 75922 471554 75978
rect 471622 75922 471678 75978
rect 471250 58294 471306 58350
rect 471374 58294 471430 58350
rect 471498 58294 471554 58350
rect 471622 58294 471678 58350
rect 471250 58170 471306 58226
rect 471374 58170 471430 58226
rect 471498 58170 471554 58226
rect 471622 58170 471678 58226
rect 471250 58046 471306 58102
rect 471374 58046 471430 58102
rect 471498 58046 471554 58102
rect 471622 58046 471678 58102
rect 471250 57922 471306 57978
rect 471374 57922 471430 57978
rect 471498 57922 471554 57978
rect 471622 57922 471678 57978
rect 471250 40294 471306 40350
rect 471374 40294 471430 40350
rect 471498 40294 471554 40350
rect 471622 40294 471678 40350
rect 471250 40170 471306 40226
rect 471374 40170 471430 40226
rect 471498 40170 471554 40226
rect 471622 40170 471678 40226
rect 471250 40046 471306 40102
rect 471374 40046 471430 40102
rect 471498 40046 471554 40102
rect 471622 40046 471678 40102
rect 471250 39922 471306 39978
rect 471374 39922 471430 39978
rect 471498 39922 471554 39978
rect 471622 39922 471678 39978
rect 471250 22294 471306 22350
rect 471374 22294 471430 22350
rect 471498 22294 471554 22350
rect 471622 22294 471678 22350
rect 471250 22170 471306 22226
rect 471374 22170 471430 22226
rect 471498 22170 471554 22226
rect 471622 22170 471678 22226
rect 471250 22046 471306 22102
rect 471374 22046 471430 22102
rect 471498 22046 471554 22102
rect 471622 22046 471678 22102
rect 471250 21922 471306 21978
rect 471374 21922 471430 21978
rect 471498 21922 471554 21978
rect 471622 21922 471678 21978
rect 471250 4294 471306 4350
rect 471374 4294 471430 4350
rect 471498 4294 471554 4350
rect 471622 4294 471678 4350
rect 471250 4170 471306 4226
rect 471374 4170 471430 4226
rect 471498 4170 471554 4226
rect 471622 4170 471678 4226
rect 471250 4046 471306 4102
rect 471374 4046 471430 4102
rect 471498 4046 471554 4102
rect 471622 4046 471678 4102
rect 471250 3922 471306 3978
rect 471374 3922 471430 3978
rect 471498 3922 471554 3978
rect 471622 3922 471678 3978
rect 471250 -216 471306 -160
rect 471374 -216 471430 -160
rect 471498 -216 471554 -160
rect 471622 -216 471678 -160
rect 471250 -340 471306 -284
rect 471374 -340 471430 -284
rect 471498 -340 471554 -284
rect 471622 -340 471678 -284
rect 471250 -464 471306 -408
rect 471374 -464 471430 -408
rect 471498 -464 471554 -408
rect 471622 -464 471678 -408
rect 471250 -588 471306 -532
rect 471374 -588 471430 -532
rect 471498 -588 471554 -532
rect 471622 -588 471678 -532
rect 474970 154294 475026 154350
rect 475094 154294 475150 154350
rect 475218 154294 475274 154350
rect 475342 154294 475398 154350
rect 474970 154170 475026 154226
rect 475094 154170 475150 154226
rect 475218 154170 475274 154226
rect 475342 154170 475398 154226
rect 474970 154046 475026 154102
rect 475094 154046 475150 154102
rect 475218 154046 475274 154102
rect 475342 154046 475398 154102
rect 474970 153922 475026 153978
rect 475094 153922 475150 153978
rect 475218 153922 475274 153978
rect 475342 153922 475398 153978
rect 474970 136294 475026 136350
rect 475094 136294 475150 136350
rect 475218 136294 475274 136350
rect 475342 136294 475398 136350
rect 474970 136170 475026 136226
rect 475094 136170 475150 136226
rect 475218 136170 475274 136226
rect 475342 136170 475398 136226
rect 474970 136046 475026 136102
rect 475094 136046 475150 136102
rect 475218 136046 475274 136102
rect 475342 136046 475398 136102
rect 474970 135922 475026 135978
rect 475094 135922 475150 135978
rect 475218 135922 475274 135978
rect 475342 135922 475398 135978
rect 474970 118294 475026 118350
rect 475094 118294 475150 118350
rect 475218 118294 475274 118350
rect 475342 118294 475398 118350
rect 474970 118170 475026 118226
rect 475094 118170 475150 118226
rect 475218 118170 475274 118226
rect 475342 118170 475398 118226
rect 474970 118046 475026 118102
rect 475094 118046 475150 118102
rect 475218 118046 475274 118102
rect 475342 118046 475398 118102
rect 474970 117922 475026 117978
rect 475094 117922 475150 117978
rect 475218 117922 475274 117978
rect 475342 117922 475398 117978
rect 474970 100294 475026 100350
rect 475094 100294 475150 100350
rect 475218 100294 475274 100350
rect 475342 100294 475398 100350
rect 474970 100170 475026 100226
rect 475094 100170 475150 100226
rect 475218 100170 475274 100226
rect 475342 100170 475398 100226
rect 474970 100046 475026 100102
rect 475094 100046 475150 100102
rect 475218 100046 475274 100102
rect 475342 100046 475398 100102
rect 474970 99922 475026 99978
rect 475094 99922 475150 99978
rect 475218 99922 475274 99978
rect 475342 99922 475398 99978
rect 474970 82294 475026 82350
rect 475094 82294 475150 82350
rect 475218 82294 475274 82350
rect 475342 82294 475398 82350
rect 474970 82170 475026 82226
rect 475094 82170 475150 82226
rect 475218 82170 475274 82226
rect 475342 82170 475398 82226
rect 474970 82046 475026 82102
rect 475094 82046 475150 82102
rect 475218 82046 475274 82102
rect 475342 82046 475398 82102
rect 474970 81922 475026 81978
rect 475094 81922 475150 81978
rect 475218 81922 475274 81978
rect 475342 81922 475398 81978
rect 474970 64294 475026 64350
rect 475094 64294 475150 64350
rect 475218 64294 475274 64350
rect 475342 64294 475398 64350
rect 474970 64170 475026 64226
rect 475094 64170 475150 64226
rect 475218 64170 475274 64226
rect 475342 64170 475398 64226
rect 474970 64046 475026 64102
rect 475094 64046 475150 64102
rect 475218 64046 475274 64102
rect 475342 64046 475398 64102
rect 474970 63922 475026 63978
rect 475094 63922 475150 63978
rect 475218 63922 475274 63978
rect 475342 63922 475398 63978
rect 474970 46294 475026 46350
rect 475094 46294 475150 46350
rect 475218 46294 475274 46350
rect 475342 46294 475398 46350
rect 474970 46170 475026 46226
rect 475094 46170 475150 46226
rect 475218 46170 475274 46226
rect 475342 46170 475398 46226
rect 474970 46046 475026 46102
rect 475094 46046 475150 46102
rect 475218 46046 475274 46102
rect 475342 46046 475398 46102
rect 474970 45922 475026 45978
rect 475094 45922 475150 45978
rect 475218 45922 475274 45978
rect 475342 45922 475398 45978
rect 474970 28294 475026 28350
rect 475094 28294 475150 28350
rect 475218 28294 475274 28350
rect 475342 28294 475398 28350
rect 474970 28170 475026 28226
rect 475094 28170 475150 28226
rect 475218 28170 475274 28226
rect 475342 28170 475398 28226
rect 474970 28046 475026 28102
rect 475094 28046 475150 28102
rect 475218 28046 475274 28102
rect 475342 28046 475398 28102
rect 474970 27922 475026 27978
rect 475094 27922 475150 27978
rect 475218 27922 475274 27978
rect 475342 27922 475398 27978
rect 474970 10294 475026 10350
rect 475094 10294 475150 10350
rect 475218 10294 475274 10350
rect 475342 10294 475398 10350
rect 474970 10170 475026 10226
rect 475094 10170 475150 10226
rect 475218 10170 475274 10226
rect 475342 10170 475398 10226
rect 474970 10046 475026 10102
rect 475094 10046 475150 10102
rect 475218 10046 475274 10102
rect 475342 10046 475398 10102
rect 474970 9922 475026 9978
rect 475094 9922 475150 9978
rect 475218 9922 475274 9978
rect 475342 9922 475398 9978
rect 474970 -1176 475026 -1120
rect 475094 -1176 475150 -1120
rect 475218 -1176 475274 -1120
rect 475342 -1176 475398 -1120
rect 474970 -1300 475026 -1244
rect 475094 -1300 475150 -1244
rect 475218 -1300 475274 -1244
rect 475342 -1300 475398 -1244
rect 474970 -1424 475026 -1368
rect 475094 -1424 475150 -1368
rect 475218 -1424 475274 -1368
rect 475342 -1424 475398 -1368
rect 474970 -1548 475026 -1492
rect 475094 -1548 475150 -1492
rect 475218 -1548 475274 -1492
rect 475342 -1548 475398 -1492
rect 489250 148294 489306 148350
rect 489374 148294 489430 148350
rect 489498 148294 489554 148350
rect 489622 148294 489678 148350
rect 489250 148170 489306 148226
rect 489374 148170 489430 148226
rect 489498 148170 489554 148226
rect 489622 148170 489678 148226
rect 489250 148046 489306 148102
rect 489374 148046 489430 148102
rect 489498 148046 489554 148102
rect 489622 148046 489678 148102
rect 489250 147922 489306 147978
rect 489374 147922 489430 147978
rect 489498 147922 489554 147978
rect 489622 147922 489678 147978
rect 489250 130294 489306 130350
rect 489374 130294 489430 130350
rect 489498 130294 489554 130350
rect 489622 130294 489678 130350
rect 489250 130170 489306 130226
rect 489374 130170 489430 130226
rect 489498 130170 489554 130226
rect 489622 130170 489678 130226
rect 489250 130046 489306 130102
rect 489374 130046 489430 130102
rect 489498 130046 489554 130102
rect 489622 130046 489678 130102
rect 489250 129922 489306 129978
rect 489374 129922 489430 129978
rect 489498 129922 489554 129978
rect 489622 129922 489678 129978
rect 489250 112294 489306 112350
rect 489374 112294 489430 112350
rect 489498 112294 489554 112350
rect 489622 112294 489678 112350
rect 489250 112170 489306 112226
rect 489374 112170 489430 112226
rect 489498 112170 489554 112226
rect 489622 112170 489678 112226
rect 489250 112046 489306 112102
rect 489374 112046 489430 112102
rect 489498 112046 489554 112102
rect 489622 112046 489678 112102
rect 489250 111922 489306 111978
rect 489374 111922 489430 111978
rect 489498 111922 489554 111978
rect 489622 111922 489678 111978
rect 489250 94294 489306 94350
rect 489374 94294 489430 94350
rect 489498 94294 489554 94350
rect 489622 94294 489678 94350
rect 489250 94170 489306 94226
rect 489374 94170 489430 94226
rect 489498 94170 489554 94226
rect 489622 94170 489678 94226
rect 489250 94046 489306 94102
rect 489374 94046 489430 94102
rect 489498 94046 489554 94102
rect 489622 94046 489678 94102
rect 489250 93922 489306 93978
rect 489374 93922 489430 93978
rect 489498 93922 489554 93978
rect 489622 93922 489678 93978
rect 489250 76294 489306 76350
rect 489374 76294 489430 76350
rect 489498 76294 489554 76350
rect 489622 76294 489678 76350
rect 489250 76170 489306 76226
rect 489374 76170 489430 76226
rect 489498 76170 489554 76226
rect 489622 76170 489678 76226
rect 489250 76046 489306 76102
rect 489374 76046 489430 76102
rect 489498 76046 489554 76102
rect 489622 76046 489678 76102
rect 489250 75922 489306 75978
rect 489374 75922 489430 75978
rect 489498 75922 489554 75978
rect 489622 75922 489678 75978
rect 489250 58294 489306 58350
rect 489374 58294 489430 58350
rect 489498 58294 489554 58350
rect 489622 58294 489678 58350
rect 489250 58170 489306 58226
rect 489374 58170 489430 58226
rect 489498 58170 489554 58226
rect 489622 58170 489678 58226
rect 489250 58046 489306 58102
rect 489374 58046 489430 58102
rect 489498 58046 489554 58102
rect 489622 58046 489678 58102
rect 489250 57922 489306 57978
rect 489374 57922 489430 57978
rect 489498 57922 489554 57978
rect 489622 57922 489678 57978
rect 489250 40294 489306 40350
rect 489374 40294 489430 40350
rect 489498 40294 489554 40350
rect 489622 40294 489678 40350
rect 489250 40170 489306 40226
rect 489374 40170 489430 40226
rect 489498 40170 489554 40226
rect 489622 40170 489678 40226
rect 489250 40046 489306 40102
rect 489374 40046 489430 40102
rect 489498 40046 489554 40102
rect 489622 40046 489678 40102
rect 489250 39922 489306 39978
rect 489374 39922 489430 39978
rect 489498 39922 489554 39978
rect 489622 39922 489678 39978
rect 489250 22294 489306 22350
rect 489374 22294 489430 22350
rect 489498 22294 489554 22350
rect 489622 22294 489678 22350
rect 489250 22170 489306 22226
rect 489374 22170 489430 22226
rect 489498 22170 489554 22226
rect 489622 22170 489678 22226
rect 489250 22046 489306 22102
rect 489374 22046 489430 22102
rect 489498 22046 489554 22102
rect 489622 22046 489678 22102
rect 489250 21922 489306 21978
rect 489374 21922 489430 21978
rect 489498 21922 489554 21978
rect 489622 21922 489678 21978
rect 489250 4294 489306 4350
rect 489374 4294 489430 4350
rect 489498 4294 489554 4350
rect 489622 4294 489678 4350
rect 489250 4170 489306 4226
rect 489374 4170 489430 4226
rect 489498 4170 489554 4226
rect 489622 4170 489678 4226
rect 489250 4046 489306 4102
rect 489374 4046 489430 4102
rect 489498 4046 489554 4102
rect 489622 4046 489678 4102
rect 489250 3922 489306 3978
rect 489374 3922 489430 3978
rect 489498 3922 489554 3978
rect 489622 3922 489678 3978
rect 489250 -216 489306 -160
rect 489374 -216 489430 -160
rect 489498 -216 489554 -160
rect 489622 -216 489678 -160
rect 489250 -340 489306 -284
rect 489374 -340 489430 -284
rect 489498 -340 489554 -284
rect 489622 -340 489678 -284
rect 489250 -464 489306 -408
rect 489374 -464 489430 -408
rect 489498 -464 489554 -408
rect 489622 -464 489678 -408
rect 489250 -588 489306 -532
rect 489374 -588 489430 -532
rect 489498 -588 489554 -532
rect 489622 -588 489678 -532
rect 492970 154294 493026 154350
rect 493094 154294 493150 154350
rect 493218 154294 493274 154350
rect 493342 154294 493398 154350
rect 492970 154170 493026 154226
rect 493094 154170 493150 154226
rect 493218 154170 493274 154226
rect 493342 154170 493398 154226
rect 492970 154046 493026 154102
rect 493094 154046 493150 154102
rect 493218 154046 493274 154102
rect 493342 154046 493398 154102
rect 492970 153922 493026 153978
rect 493094 153922 493150 153978
rect 493218 153922 493274 153978
rect 493342 153922 493398 153978
rect 492970 136294 493026 136350
rect 493094 136294 493150 136350
rect 493218 136294 493274 136350
rect 493342 136294 493398 136350
rect 492970 136170 493026 136226
rect 493094 136170 493150 136226
rect 493218 136170 493274 136226
rect 493342 136170 493398 136226
rect 492970 136046 493026 136102
rect 493094 136046 493150 136102
rect 493218 136046 493274 136102
rect 493342 136046 493398 136102
rect 492970 135922 493026 135978
rect 493094 135922 493150 135978
rect 493218 135922 493274 135978
rect 493342 135922 493398 135978
rect 492970 118294 493026 118350
rect 493094 118294 493150 118350
rect 493218 118294 493274 118350
rect 493342 118294 493398 118350
rect 492970 118170 493026 118226
rect 493094 118170 493150 118226
rect 493218 118170 493274 118226
rect 493342 118170 493398 118226
rect 492970 118046 493026 118102
rect 493094 118046 493150 118102
rect 493218 118046 493274 118102
rect 493342 118046 493398 118102
rect 492970 117922 493026 117978
rect 493094 117922 493150 117978
rect 493218 117922 493274 117978
rect 493342 117922 493398 117978
rect 492970 100294 493026 100350
rect 493094 100294 493150 100350
rect 493218 100294 493274 100350
rect 493342 100294 493398 100350
rect 492970 100170 493026 100226
rect 493094 100170 493150 100226
rect 493218 100170 493274 100226
rect 493342 100170 493398 100226
rect 492970 100046 493026 100102
rect 493094 100046 493150 100102
rect 493218 100046 493274 100102
rect 493342 100046 493398 100102
rect 492970 99922 493026 99978
rect 493094 99922 493150 99978
rect 493218 99922 493274 99978
rect 493342 99922 493398 99978
rect 492970 82294 493026 82350
rect 493094 82294 493150 82350
rect 493218 82294 493274 82350
rect 493342 82294 493398 82350
rect 492970 82170 493026 82226
rect 493094 82170 493150 82226
rect 493218 82170 493274 82226
rect 493342 82170 493398 82226
rect 492970 82046 493026 82102
rect 493094 82046 493150 82102
rect 493218 82046 493274 82102
rect 493342 82046 493398 82102
rect 492970 81922 493026 81978
rect 493094 81922 493150 81978
rect 493218 81922 493274 81978
rect 493342 81922 493398 81978
rect 492970 64294 493026 64350
rect 493094 64294 493150 64350
rect 493218 64294 493274 64350
rect 493342 64294 493398 64350
rect 492970 64170 493026 64226
rect 493094 64170 493150 64226
rect 493218 64170 493274 64226
rect 493342 64170 493398 64226
rect 492970 64046 493026 64102
rect 493094 64046 493150 64102
rect 493218 64046 493274 64102
rect 493342 64046 493398 64102
rect 492970 63922 493026 63978
rect 493094 63922 493150 63978
rect 493218 63922 493274 63978
rect 493342 63922 493398 63978
rect 492970 46294 493026 46350
rect 493094 46294 493150 46350
rect 493218 46294 493274 46350
rect 493342 46294 493398 46350
rect 492970 46170 493026 46226
rect 493094 46170 493150 46226
rect 493218 46170 493274 46226
rect 493342 46170 493398 46226
rect 492970 46046 493026 46102
rect 493094 46046 493150 46102
rect 493218 46046 493274 46102
rect 493342 46046 493398 46102
rect 492970 45922 493026 45978
rect 493094 45922 493150 45978
rect 493218 45922 493274 45978
rect 493342 45922 493398 45978
rect 492970 28294 493026 28350
rect 493094 28294 493150 28350
rect 493218 28294 493274 28350
rect 493342 28294 493398 28350
rect 492970 28170 493026 28226
rect 493094 28170 493150 28226
rect 493218 28170 493274 28226
rect 493342 28170 493398 28226
rect 492970 28046 493026 28102
rect 493094 28046 493150 28102
rect 493218 28046 493274 28102
rect 493342 28046 493398 28102
rect 492970 27922 493026 27978
rect 493094 27922 493150 27978
rect 493218 27922 493274 27978
rect 493342 27922 493398 27978
rect 492970 10294 493026 10350
rect 493094 10294 493150 10350
rect 493218 10294 493274 10350
rect 493342 10294 493398 10350
rect 492970 10170 493026 10226
rect 493094 10170 493150 10226
rect 493218 10170 493274 10226
rect 493342 10170 493398 10226
rect 492970 10046 493026 10102
rect 493094 10046 493150 10102
rect 493218 10046 493274 10102
rect 493342 10046 493398 10102
rect 492970 9922 493026 9978
rect 493094 9922 493150 9978
rect 493218 9922 493274 9978
rect 493342 9922 493398 9978
rect 492970 -1176 493026 -1120
rect 493094 -1176 493150 -1120
rect 493218 -1176 493274 -1120
rect 493342 -1176 493398 -1120
rect 492970 -1300 493026 -1244
rect 493094 -1300 493150 -1244
rect 493218 -1300 493274 -1244
rect 493342 -1300 493398 -1244
rect 492970 -1424 493026 -1368
rect 493094 -1424 493150 -1368
rect 493218 -1424 493274 -1368
rect 493342 -1424 493398 -1368
rect 492970 -1548 493026 -1492
rect 493094 -1548 493150 -1492
rect 493218 -1548 493274 -1492
rect 493342 -1548 493398 -1492
rect 507250 148294 507306 148350
rect 507374 148294 507430 148350
rect 507498 148294 507554 148350
rect 507622 148294 507678 148350
rect 507250 148170 507306 148226
rect 507374 148170 507430 148226
rect 507498 148170 507554 148226
rect 507622 148170 507678 148226
rect 507250 148046 507306 148102
rect 507374 148046 507430 148102
rect 507498 148046 507554 148102
rect 507622 148046 507678 148102
rect 507250 147922 507306 147978
rect 507374 147922 507430 147978
rect 507498 147922 507554 147978
rect 507622 147922 507678 147978
rect 507250 130294 507306 130350
rect 507374 130294 507430 130350
rect 507498 130294 507554 130350
rect 507622 130294 507678 130350
rect 507250 130170 507306 130226
rect 507374 130170 507430 130226
rect 507498 130170 507554 130226
rect 507622 130170 507678 130226
rect 507250 130046 507306 130102
rect 507374 130046 507430 130102
rect 507498 130046 507554 130102
rect 507622 130046 507678 130102
rect 507250 129922 507306 129978
rect 507374 129922 507430 129978
rect 507498 129922 507554 129978
rect 507622 129922 507678 129978
rect 507250 112294 507306 112350
rect 507374 112294 507430 112350
rect 507498 112294 507554 112350
rect 507622 112294 507678 112350
rect 507250 112170 507306 112226
rect 507374 112170 507430 112226
rect 507498 112170 507554 112226
rect 507622 112170 507678 112226
rect 507250 112046 507306 112102
rect 507374 112046 507430 112102
rect 507498 112046 507554 112102
rect 507622 112046 507678 112102
rect 507250 111922 507306 111978
rect 507374 111922 507430 111978
rect 507498 111922 507554 111978
rect 507622 111922 507678 111978
rect 507250 94294 507306 94350
rect 507374 94294 507430 94350
rect 507498 94294 507554 94350
rect 507622 94294 507678 94350
rect 507250 94170 507306 94226
rect 507374 94170 507430 94226
rect 507498 94170 507554 94226
rect 507622 94170 507678 94226
rect 507250 94046 507306 94102
rect 507374 94046 507430 94102
rect 507498 94046 507554 94102
rect 507622 94046 507678 94102
rect 507250 93922 507306 93978
rect 507374 93922 507430 93978
rect 507498 93922 507554 93978
rect 507622 93922 507678 93978
rect 507250 76294 507306 76350
rect 507374 76294 507430 76350
rect 507498 76294 507554 76350
rect 507622 76294 507678 76350
rect 507250 76170 507306 76226
rect 507374 76170 507430 76226
rect 507498 76170 507554 76226
rect 507622 76170 507678 76226
rect 507250 76046 507306 76102
rect 507374 76046 507430 76102
rect 507498 76046 507554 76102
rect 507622 76046 507678 76102
rect 507250 75922 507306 75978
rect 507374 75922 507430 75978
rect 507498 75922 507554 75978
rect 507622 75922 507678 75978
rect 507250 58294 507306 58350
rect 507374 58294 507430 58350
rect 507498 58294 507554 58350
rect 507622 58294 507678 58350
rect 507250 58170 507306 58226
rect 507374 58170 507430 58226
rect 507498 58170 507554 58226
rect 507622 58170 507678 58226
rect 507250 58046 507306 58102
rect 507374 58046 507430 58102
rect 507498 58046 507554 58102
rect 507622 58046 507678 58102
rect 507250 57922 507306 57978
rect 507374 57922 507430 57978
rect 507498 57922 507554 57978
rect 507622 57922 507678 57978
rect 507250 40294 507306 40350
rect 507374 40294 507430 40350
rect 507498 40294 507554 40350
rect 507622 40294 507678 40350
rect 507250 40170 507306 40226
rect 507374 40170 507430 40226
rect 507498 40170 507554 40226
rect 507622 40170 507678 40226
rect 507250 40046 507306 40102
rect 507374 40046 507430 40102
rect 507498 40046 507554 40102
rect 507622 40046 507678 40102
rect 507250 39922 507306 39978
rect 507374 39922 507430 39978
rect 507498 39922 507554 39978
rect 507622 39922 507678 39978
rect 507250 22294 507306 22350
rect 507374 22294 507430 22350
rect 507498 22294 507554 22350
rect 507622 22294 507678 22350
rect 507250 22170 507306 22226
rect 507374 22170 507430 22226
rect 507498 22170 507554 22226
rect 507622 22170 507678 22226
rect 507250 22046 507306 22102
rect 507374 22046 507430 22102
rect 507498 22046 507554 22102
rect 507622 22046 507678 22102
rect 507250 21922 507306 21978
rect 507374 21922 507430 21978
rect 507498 21922 507554 21978
rect 507622 21922 507678 21978
rect 507250 4294 507306 4350
rect 507374 4294 507430 4350
rect 507498 4294 507554 4350
rect 507622 4294 507678 4350
rect 507250 4170 507306 4226
rect 507374 4170 507430 4226
rect 507498 4170 507554 4226
rect 507622 4170 507678 4226
rect 507250 4046 507306 4102
rect 507374 4046 507430 4102
rect 507498 4046 507554 4102
rect 507622 4046 507678 4102
rect 507250 3922 507306 3978
rect 507374 3922 507430 3978
rect 507498 3922 507554 3978
rect 507622 3922 507678 3978
rect 507250 -216 507306 -160
rect 507374 -216 507430 -160
rect 507498 -216 507554 -160
rect 507622 -216 507678 -160
rect 507250 -340 507306 -284
rect 507374 -340 507430 -284
rect 507498 -340 507554 -284
rect 507622 -340 507678 -284
rect 507250 -464 507306 -408
rect 507374 -464 507430 -408
rect 507498 -464 507554 -408
rect 507622 -464 507678 -408
rect 507250 -588 507306 -532
rect 507374 -588 507430 -532
rect 507498 -588 507554 -532
rect 507622 -588 507678 -532
rect 510970 154294 511026 154350
rect 511094 154294 511150 154350
rect 511218 154294 511274 154350
rect 511342 154294 511398 154350
rect 510970 154170 511026 154226
rect 511094 154170 511150 154226
rect 511218 154170 511274 154226
rect 511342 154170 511398 154226
rect 510970 154046 511026 154102
rect 511094 154046 511150 154102
rect 511218 154046 511274 154102
rect 511342 154046 511398 154102
rect 510970 153922 511026 153978
rect 511094 153922 511150 153978
rect 511218 153922 511274 153978
rect 511342 153922 511398 153978
rect 510970 136294 511026 136350
rect 511094 136294 511150 136350
rect 511218 136294 511274 136350
rect 511342 136294 511398 136350
rect 510970 136170 511026 136226
rect 511094 136170 511150 136226
rect 511218 136170 511274 136226
rect 511342 136170 511398 136226
rect 510970 136046 511026 136102
rect 511094 136046 511150 136102
rect 511218 136046 511274 136102
rect 511342 136046 511398 136102
rect 510970 135922 511026 135978
rect 511094 135922 511150 135978
rect 511218 135922 511274 135978
rect 511342 135922 511398 135978
rect 510970 118294 511026 118350
rect 511094 118294 511150 118350
rect 511218 118294 511274 118350
rect 511342 118294 511398 118350
rect 510970 118170 511026 118226
rect 511094 118170 511150 118226
rect 511218 118170 511274 118226
rect 511342 118170 511398 118226
rect 510970 118046 511026 118102
rect 511094 118046 511150 118102
rect 511218 118046 511274 118102
rect 511342 118046 511398 118102
rect 510970 117922 511026 117978
rect 511094 117922 511150 117978
rect 511218 117922 511274 117978
rect 511342 117922 511398 117978
rect 510970 100294 511026 100350
rect 511094 100294 511150 100350
rect 511218 100294 511274 100350
rect 511342 100294 511398 100350
rect 510970 100170 511026 100226
rect 511094 100170 511150 100226
rect 511218 100170 511274 100226
rect 511342 100170 511398 100226
rect 510970 100046 511026 100102
rect 511094 100046 511150 100102
rect 511218 100046 511274 100102
rect 511342 100046 511398 100102
rect 510970 99922 511026 99978
rect 511094 99922 511150 99978
rect 511218 99922 511274 99978
rect 511342 99922 511398 99978
rect 525250 148294 525306 148350
rect 525374 148294 525430 148350
rect 525498 148294 525554 148350
rect 525622 148294 525678 148350
rect 525250 148170 525306 148226
rect 525374 148170 525430 148226
rect 525498 148170 525554 148226
rect 525622 148170 525678 148226
rect 525250 148046 525306 148102
rect 525374 148046 525430 148102
rect 525498 148046 525554 148102
rect 525622 148046 525678 148102
rect 525250 147922 525306 147978
rect 525374 147922 525430 147978
rect 525498 147922 525554 147978
rect 525622 147922 525678 147978
rect 525250 130294 525306 130350
rect 525374 130294 525430 130350
rect 525498 130294 525554 130350
rect 525622 130294 525678 130350
rect 525250 130170 525306 130226
rect 525374 130170 525430 130226
rect 525498 130170 525554 130226
rect 525622 130170 525678 130226
rect 525250 130046 525306 130102
rect 525374 130046 525430 130102
rect 525498 130046 525554 130102
rect 525622 130046 525678 130102
rect 525250 129922 525306 129978
rect 525374 129922 525430 129978
rect 525498 129922 525554 129978
rect 525622 129922 525678 129978
rect 525250 112294 525306 112350
rect 525374 112294 525430 112350
rect 525498 112294 525554 112350
rect 525622 112294 525678 112350
rect 525250 112170 525306 112226
rect 525374 112170 525430 112226
rect 525498 112170 525554 112226
rect 525622 112170 525678 112226
rect 525250 112046 525306 112102
rect 525374 112046 525430 112102
rect 525498 112046 525554 112102
rect 525622 112046 525678 112102
rect 525250 111922 525306 111978
rect 525374 111922 525430 111978
rect 525498 111922 525554 111978
rect 525622 111922 525678 111978
rect 524518 94294 524574 94350
rect 524642 94294 524698 94350
rect 524518 94170 524574 94226
rect 524642 94170 524698 94226
rect 524518 94046 524574 94102
rect 524642 94046 524698 94102
rect 524518 93922 524574 93978
rect 524642 93922 524698 93978
rect 525250 94294 525306 94350
rect 525374 94294 525430 94350
rect 525498 94294 525554 94350
rect 525622 94294 525678 94350
rect 525250 94170 525306 94226
rect 525374 94170 525430 94226
rect 525498 94170 525554 94226
rect 525622 94170 525678 94226
rect 525250 94046 525306 94102
rect 525374 94046 525430 94102
rect 525498 94046 525554 94102
rect 525622 94046 525678 94102
rect 525250 93922 525306 93978
rect 525374 93922 525430 93978
rect 525498 93922 525554 93978
rect 525622 93922 525678 93978
rect 510970 82294 511026 82350
rect 511094 82294 511150 82350
rect 511218 82294 511274 82350
rect 511342 82294 511398 82350
rect 510970 82170 511026 82226
rect 511094 82170 511150 82226
rect 511218 82170 511274 82226
rect 511342 82170 511398 82226
rect 510970 82046 511026 82102
rect 511094 82046 511150 82102
rect 511218 82046 511274 82102
rect 511342 82046 511398 82102
rect 510970 81922 511026 81978
rect 511094 81922 511150 81978
rect 511218 81922 511274 81978
rect 511342 81922 511398 81978
rect 524518 76294 524574 76350
rect 524642 76294 524698 76350
rect 524518 76170 524574 76226
rect 524642 76170 524698 76226
rect 524518 76046 524574 76102
rect 524642 76046 524698 76102
rect 524518 75922 524574 75978
rect 524642 75922 524698 75978
rect 525250 76294 525306 76350
rect 525374 76294 525430 76350
rect 525498 76294 525554 76350
rect 525622 76294 525678 76350
rect 525250 76170 525306 76226
rect 525374 76170 525430 76226
rect 525498 76170 525554 76226
rect 525622 76170 525678 76226
rect 525250 76046 525306 76102
rect 525374 76046 525430 76102
rect 525498 76046 525554 76102
rect 525622 76046 525678 76102
rect 525250 75922 525306 75978
rect 525374 75922 525430 75978
rect 525498 75922 525554 75978
rect 525622 75922 525678 75978
rect 510970 64294 511026 64350
rect 511094 64294 511150 64350
rect 511218 64294 511274 64350
rect 511342 64294 511398 64350
rect 510970 64170 511026 64226
rect 511094 64170 511150 64226
rect 511218 64170 511274 64226
rect 511342 64170 511398 64226
rect 510970 64046 511026 64102
rect 511094 64046 511150 64102
rect 511218 64046 511274 64102
rect 511342 64046 511398 64102
rect 510970 63922 511026 63978
rect 511094 63922 511150 63978
rect 511218 63922 511274 63978
rect 511342 63922 511398 63978
rect 510970 46294 511026 46350
rect 511094 46294 511150 46350
rect 511218 46294 511274 46350
rect 511342 46294 511398 46350
rect 510970 46170 511026 46226
rect 511094 46170 511150 46226
rect 511218 46170 511274 46226
rect 511342 46170 511398 46226
rect 510970 46046 511026 46102
rect 511094 46046 511150 46102
rect 511218 46046 511274 46102
rect 511342 46046 511398 46102
rect 510970 45922 511026 45978
rect 511094 45922 511150 45978
rect 511218 45922 511274 45978
rect 511342 45922 511398 45978
rect 510970 28294 511026 28350
rect 511094 28294 511150 28350
rect 511218 28294 511274 28350
rect 511342 28294 511398 28350
rect 510970 28170 511026 28226
rect 511094 28170 511150 28226
rect 511218 28170 511274 28226
rect 511342 28170 511398 28226
rect 510970 28046 511026 28102
rect 511094 28046 511150 28102
rect 511218 28046 511274 28102
rect 511342 28046 511398 28102
rect 510970 27922 511026 27978
rect 511094 27922 511150 27978
rect 511218 27922 511274 27978
rect 511342 27922 511398 27978
rect 510970 10294 511026 10350
rect 511094 10294 511150 10350
rect 511218 10294 511274 10350
rect 511342 10294 511398 10350
rect 510970 10170 511026 10226
rect 511094 10170 511150 10226
rect 511218 10170 511274 10226
rect 511342 10170 511398 10226
rect 510970 10046 511026 10102
rect 511094 10046 511150 10102
rect 511218 10046 511274 10102
rect 511342 10046 511398 10102
rect 510970 9922 511026 9978
rect 511094 9922 511150 9978
rect 511218 9922 511274 9978
rect 511342 9922 511398 9978
rect 510970 -1176 511026 -1120
rect 511094 -1176 511150 -1120
rect 511218 -1176 511274 -1120
rect 511342 -1176 511398 -1120
rect 510970 -1300 511026 -1244
rect 511094 -1300 511150 -1244
rect 511218 -1300 511274 -1244
rect 511342 -1300 511398 -1244
rect 510970 -1424 511026 -1368
rect 511094 -1424 511150 -1368
rect 511218 -1424 511274 -1368
rect 511342 -1424 511398 -1368
rect 510970 -1548 511026 -1492
rect 511094 -1548 511150 -1492
rect 511218 -1548 511274 -1492
rect 511342 -1548 511398 -1492
rect 525250 58294 525306 58350
rect 525374 58294 525430 58350
rect 525498 58294 525554 58350
rect 525622 58294 525678 58350
rect 525250 58170 525306 58226
rect 525374 58170 525430 58226
rect 525498 58170 525554 58226
rect 525622 58170 525678 58226
rect 525250 58046 525306 58102
rect 525374 58046 525430 58102
rect 525498 58046 525554 58102
rect 525622 58046 525678 58102
rect 525250 57922 525306 57978
rect 525374 57922 525430 57978
rect 525498 57922 525554 57978
rect 525622 57922 525678 57978
rect 525250 40294 525306 40350
rect 525374 40294 525430 40350
rect 525498 40294 525554 40350
rect 525622 40294 525678 40350
rect 525250 40170 525306 40226
rect 525374 40170 525430 40226
rect 525498 40170 525554 40226
rect 525622 40170 525678 40226
rect 525250 40046 525306 40102
rect 525374 40046 525430 40102
rect 525498 40046 525554 40102
rect 525622 40046 525678 40102
rect 525250 39922 525306 39978
rect 525374 39922 525430 39978
rect 525498 39922 525554 39978
rect 525622 39922 525678 39978
rect 525250 22294 525306 22350
rect 525374 22294 525430 22350
rect 525498 22294 525554 22350
rect 525622 22294 525678 22350
rect 525250 22170 525306 22226
rect 525374 22170 525430 22226
rect 525498 22170 525554 22226
rect 525622 22170 525678 22226
rect 525250 22046 525306 22102
rect 525374 22046 525430 22102
rect 525498 22046 525554 22102
rect 525622 22046 525678 22102
rect 525250 21922 525306 21978
rect 525374 21922 525430 21978
rect 525498 21922 525554 21978
rect 525622 21922 525678 21978
rect 525250 4294 525306 4350
rect 525374 4294 525430 4350
rect 525498 4294 525554 4350
rect 525622 4294 525678 4350
rect 525250 4170 525306 4226
rect 525374 4170 525430 4226
rect 525498 4170 525554 4226
rect 525622 4170 525678 4226
rect 528970 154294 529026 154350
rect 529094 154294 529150 154350
rect 529218 154294 529274 154350
rect 529342 154294 529398 154350
rect 528970 154170 529026 154226
rect 529094 154170 529150 154226
rect 529218 154170 529274 154226
rect 529342 154170 529398 154226
rect 528970 154046 529026 154102
rect 529094 154046 529150 154102
rect 529218 154046 529274 154102
rect 529342 154046 529398 154102
rect 528970 153922 529026 153978
rect 529094 153922 529150 153978
rect 529218 153922 529274 153978
rect 529342 153922 529398 153978
rect 528970 136294 529026 136350
rect 529094 136294 529150 136350
rect 529218 136294 529274 136350
rect 529342 136294 529398 136350
rect 528970 136170 529026 136226
rect 529094 136170 529150 136226
rect 529218 136170 529274 136226
rect 529342 136170 529398 136226
rect 528970 136046 529026 136102
rect 529094 136046 529150 136102
rect 529218 136046 529274 136102
rect 529342 136046 529398 136102
rect 528970 135922 529026 135978
rect 529094 135922 529150 135978
rect 529218 135922 529274 135978
rect 529342 135922 529398 135978
rect 528970 118294 529026 118350
rect 529094 118294 529150 118350
rect 529218 118294 529274 118350
rect 529342 118294 529398 118350
rect 528970 118170 529026 118226
rect 529094 118170 529150 118226
rect 529218 118170 529274 118226
rect 529342 118170 529398 118226
rect 528970 118046 529026 118102
rect 529094 118046 529150 118102
rect 529218 118046 529274 118102
rect 529342 118046 529398 118102
rect 528970 117922 529026 117978
rect 529094 117922 529150 117978
rect 529218 117922 529274 117978
rect 529342 117922 529398 117978
rect 543250 148294 543306 148350
rect 543374 148294 543430 148350
rect 543498 148294 543554 148350
rect 543622 148294 543678 148350
rect 543250 148170 543306 148226
rect 543374 148170 543430 148226
rect 543498 148170 543554 148226
rect 543622 148170 543678 148226
rect 543250 148046 543306 148102
rect 543374 148046 543430 148102
rect 543498 148046 543554 148102
rect 543622 148046 543678 148102
rect 543250 147922 543306 147978
rect 543374 147922 543430 147978
rect 543498 147922 543554 147978
rect 543622 147922 543678 147978
rect 543250 130294 543306 130350
rect 543374 130294 543430 130350
rect 543498 130294 543554 130350
rect 543622 130294 543678 130350
rect 543250 130170 543306 130226
rect 543374 130170 543430 130226
rect 543498 130170 543554 130226
rect 543622 130170 543678 130226
rect 543250 130046 543306 130102
rect 543374 130046 543430 130102
rect 543498 130046 543554 130102
rect 543622 130046 543678 130102
rect 543250 129922 543306 129978
rect 543374 129922 543430 129978
rect 543498 129922 543554 129978
rect 543622 129922 543678 129978
rect 543250 112294 543306 112350
rect 543374 112294 543430 112350
rect 543498 112294 543554 112350
rect 543622 112294 543678 112350
rect 543250 112170 543306 112226
rect 543374 112170 543430 112226
rect 543498 112170 543554 112226
rect 543622 112170 543678 112226
rect 543250 112046 543306 112102
rect 543374 112046 543430 112102
rect 543498 112046 543554 112102
rect 543622 112046 543678 112102
rect 543250 111922 543306 111978
rect 543374 111922 543430 111978
rect 543498 111922 543554 111978
rect 543622 111922 543678 111978
rect 528970 100294 529026 100350
rect 529094 100294 529150 100350
rect 529218 100294 529274 100350
rect 529342 100294 529398 100350
rect 528970 100170 529026 100226
rect 529094 100170 529150 100226
rect 529218 100170 529274 100226
rect 529342 100170 529398 100226
rect 528970 100046 529026 100102
rect 529094 100046 529150 100102
rect 529218 100046 529274 100102
rect 529342 100046 529398 100102
rect 528970 99922 529026 99978
rect 529094 99922 529150 99978
rect 529218 99922 529274 99978
rect 529342 99922 529398 99978
rect 539878 100294 539934 100350
rect 540002 100294 540058 100350
rect 539878 100170 539934 100226
rect 540002 100170 540058 100226
rect 539878 100046 539934 100102
rect 540002 100046 540058 100102
rect 539878 99922 539934 99978
rect 540002 99922 540058 99978
rect 543250 94294 543306 94350
rect 543374 94294 543430 94350
rect 543498 94294 543554 94350
rect 543622 94294 543678 94350
rect 543250 94170 543306 94226
rect 543374 94170 543430 94226
rect 543498 94170 543554 94226
rect 543622 94170 543678 94226
rect 543250 94046 543306 94102
rect 543374 94046 543430 94102
rect 543498 94046 543554 94102
rect 543622 94046 543678 94102
rect 543250 93922 543306 93978
rect 543374 93922 543430 93978
rect 543498 93922 543554 93978
rect 543622 93922 543678 93978
rect 528970 82294 529026 82350
rect 529094 82294 529150 82350
rect 529218 82294 529274 82350
rect 529342 82294 529398 82350
rect 528970 82170 529026 82226
rect 529094 82170 529150 82226
rect 529218 82170 529274 82226
rect 529342 82170 529398 82226
rect 528970 82046 529026 82102
rect 529094 82046 529150 82102
rect 529218 82046 529274 82102
rect 529342 82046 529398 82102
rect 528970 81922 529026 81978
rect 529094 81922 529150 81978
rect 529218 81922 529274 81978
rect 529342 81922 529398 81978
rect 539878 82294 539934 82350
rect 540002 82294 540058 82350
rect 539878 82170 539934 82226
rect 540002 82170 540058 82226
rect 539878 82046 539934 82102
rect 540002 82046 540058 82102
rect 539878 81922 539934 81978
rect 540002 81922 540058 81978
rect 543250 76294 543306 76350
rect 543374 76294 543430 76350
rect 543498 76294 543554 76350
rect 543622 76294 543678 76350
rect 543250 76170 543306 76226
rect 543374 76170 543430 76226
rect 543498 76170 543554 76226
rect 543622 76170 543678 76226
rect 543250 76046 543306 76102
rect 543374 76046 543430 76102
rect 543498 76046 543554 76102
rect 543622 76046 543678 76102
rect 543250 75922 543306 75978
rect 543374 75922 543430 75978
rect 543498 75922 543554 75978
rect 543622 75922 543678 75978
rect 528970 64294 529026 64350
rect 529094 64294 529150 64350
rect 529218 64294 529274 64350
rect 529342 64294 529398 64350
rect 528970 64170 529026 64226
rect 529094 64170 529150 64226
rect 529218 64170 529274 64226
rect 529342 64170 529398 64226
rect 528970 64046 529026 64102
rect 529094 64046 529150 64102
rect 529218 64046 529274 64102
rect 529342 64046 529398 64102
rect 528970 63922 529026 63978
rect 529094 63922 529150 63978
rect 529218 63922 529274 63978
rect 529342 63922 529398 63978
rect 539878 64294 539934 64350
rect 540002 64294 540058 64350
rect 539878 64170 539934 64226
rect 540002 64170 540058 64226
rect 539878 64046 539934 64102
rect 540002 64046 540058 64102
rect 539878 63922 539934 63978
rect 540002 63922 540058 63978
rect 528970 46294 529026 46350
rect 529094 46294 529150 46350
rect 529218 46294 529274 46350
rect 529342 46294 529398 46350
rect 528970 46170 529026 46226
rect 529094 46170 529150 46226
rect 529218 46170 529274 46226
rect 529342 46170 529398 46226
rect 528970 46046 529026 46102
rect 529094 46046 529150 46102
rect 529218 46046 529274 46102
rect 529342 46046 529398 46102
rect 528970 45922 529026 45978
rect 529094 45922 529150 45978
rect 529218 45922 529274 45978
rect 529342 45922 529398 45978
rect 528970 28294 529026 28350
rect 529094 28294 529150 28350
rect 529218 28294 529274 28350
rect 529342 28294 529398 28350
rect 528970 28170 529026 28226
rect 529094 28170 529150 28226
rect 529218 28170 529274 28226
rect 529342 28170 529398 28226
rect 528970 28046 529026 28102
rect 529094 28046 529150 28102
rect 529218 28046 529274 28102
rect 529342 28046 529398 28102
rect 528970 27922 529026 27978
rect 529094 27922 529150 27978
rect 529218 27922 529274 27978
rect 529342 27922 529398 27978
rect 528970 10294 529026 10350
rect 529094 10294 529150 10350
rect 529218 10294 529274 10350
rect 529342 10294 529398 10350
rect 528970 10170 529026 10226
rect 529094 10170 529150 10226
rect 529218 10170 529274 10226
rect 529342 10170 529398 10226
rect 528970 10046 529026 10102
rect 529094 10046 529150 10102
rect 529218 10046 529274 10102
rect 529342 10046 529398 10102
rect 528970 9922 529026 9978
rect 529094 9922 529150 9978
rect 529218 9922 529274 9978
rect 529342 9922 529398 9978
rect 525250 4046 525306 4102
rect 525374 4046 525430 4102
rect 525498 4046 525554 4102
rect 525622 4046 525678 4102
rect 525250 3922 525306 3978
rect 525374 3922 525430 3978
rect 525498 3922 525554 3978
rect 525622 3922 525678 3978
rect 525250 -216 525306 -160
rect 525374 -216 525430 -160
rect 525498 -216 525554 -160
rect 525622 -216 525678 -160
rect 525250 -340 525306 -284
rect 525374 -340 525430 -284
rect 525498 -340 525554 -284
rect 525622 -340 525678 -284
rect 525250 -464 525306 -408
rect 525374 -464 525430 -408
rect 525498 -464 525554 -408
rect 525622 -464 525678 -408
rect 525250 -588 525306 -532
rect 525374 -588 525430 -532
rect 525498 -588 525554 -532
rect 525622 -588 525678 -532
rect 528970 -1176 529026 -1120
rect 529094 -1176 529150 -1120
rect 529218 -1176 529274 -1120
rect 529342 -1176 529398 -1120
rect 528970 -1300 529026 -1244
rect 529094 -1300 529150 -1244
rect 529218 -1300 529274 -1244
rect 529342 -1300 529398 -1244
rect 528970 -1424 529026 -1368
rect 529094 -1424 529150 -1368
rect 529218 -1424 529274 -1368
rect 529342 -1424 529398 -1368
rect 528970 -1548 529026 -1492
rect 529094 -1548 529150 -1492
rect 529218 -1548 529274 -1492
rect 529342 -1548 529398 -1492
rect 543250 58294 543306 58350
rect 543374 58294 543430 58350
rect 543498 58294 543554 58350
rect 543622 58294 543678 58350
rect 543250 58170 543306 58226
rect 543374 58170 543430 58226
rect 543498 58170 543554 58226
rect 543622 58170 543678 58226
rect 543250 58046 543306 58102
rect 543374 58046 543430 58102
rect 543498 58046 543554 58102
rect 543622 58046 543678 58102
rect 543250 57922 543306 57978
rect 543374 57922 543430 57978
rect 543498 57922 543554 57978
rect 543622 57922 543678 57978
rect 543250 40294 543306 40350
rect 543374 40294 543430 40350
rect 543498 40294 543554 40350
rect 543622 40294 543678 40350
rect 543250 40170 543306 40226
rect 543374 40170 543430 40226
rect 543498 40170 543554 40226
rect 543622 40170 543678 40226
rect 543250 40046 543306 40102
rect 543374 40046 543430 40102
rect 543498 40046 543554 40102
rect 543622 40046 543678 40102
rect 543250 39922 543306 39978
rect 543374 39922 543430 39978
rect 543498 39922 543554 39978
rect 543622 39922 543678 39978
rect 543250 22294 543306 22350
rect 543374 22294 543430 22350
rect 543498 22294 543554 22350
rect 543622 22294 543678 22350
rect 543250 22170 543306 22226
rect 543374 22170 543430 22226
rect 543498 22170 543554 22226
rect 543622 22170 543678 22226
rect 543250 22046 543306 22102
rect 543374 22046 543430 22102
rect 543498 22046 543554 22102
rect 543622 22046 543678 22102
rect 543250 21922 543306 21978
rect 543374 21922 543430 21978
rect 543498 21922 543554 21978
rect 543622 21922 543678 21978
rect 543250 4294 543306 4350
rect 543374 4294 543430 4350
rect 543498 4294 543554 4350
rect 543622 4294 543678 4350
rect 543250 4170 543306 4226
rect 543374 4170 543430 4226
rect 543498 4170 543554 4226
rect 543622 4170 543678 4226
rect 543250 4046 543306 4102
rect 543374 4046 543430 4102
rect 543498 4046 543554 4102
rect 543622 4046 543678 4102
rect 543250 3922 543306 3978
rect 543374 3922 543430 3978
rect 543498 3922 543554 3978
rect 543622 3922 543678 3978
rect 543250 -216 543306 -160
rect 543374 -216 543430 -160
rect 543498 -216 543554 -160
rect 543622 -216 543678 -160
rect 543250 -340 543306 -284
rect 543374 -340 543430 -284
rect 543498 -340 543554 -284
rect 543622 -340 543678 -284
rect 543250 -464 543306 -408
rect 543374 -464 543430 -408
rect 543498 -464 543554 -408
rect 543622 -464 543678 -408
rect 543250 -588 543306 -532
rect 543374 -588 543430 -532
rect 543498 -588 543554 -532
rect 543622 -588 543678 -532
rect 546970 154294 547026 154350
rect 547094 154294 547150 154350
rect 547218 154294 547274 154350
rect 547342 154294 547398 154350
rect 546970 154170 547026 154226
rect 547094 154170 547150 154226
rect 547218 154170 547274 154226
rect 547342 154170 547398 154226
rect 546970 154046 547026 154102
rect 547094 154046 547150 154102
rect 547218 154046 547274 154102
rect 547342 154046 547398 154102
rect 546970 153922 547026 153978
rect 547094 153922 547150 153978
rect 547218 153922 547274 153978
rect 547342 153922 547398 153978
rect 546970 136294 547026 136350
rect 547094 136294 547150 136350
rect 547218 136294 547274 136350
rect 547342 136294 547398 136350
rect 546970 136170 547026 136226
rect 547094 136170 547150 136226
rect 547218 136170 547274 136226
rect 547342 136170 547398 136226
rect 546970 136046 547026 136102
rect 547094 136046 547150 136102
rect 547218 136046 547274 136102
rect 547342 136046 547398 136102
rect 546970 135922 547026 135978
rect 547094 135922 547150 135978
rect 547218 135922 547274 135978
rect 547342 135922 547398 135978
rect 546970 118294 547026 118350
rect 547094 118294 547150 118350
rect 547218 118294 547274 118350
rect 547342 118294 547398 118350
rect 546970 118170 547026 118226
rect 547094 118170 547150 118226
rect 547218 118170 547274 118226
rect 547342 118170 547398 118226
rect 546970 118046 547026 118102
rect 547094 118046 547150 118102
rect 547218 118046 547274 118102
rect 547342 118046 547398 118102
rect 546970 117922 547026 117978
rect 547094 117922 547150 117978
rect 547218 117922 547274 117978
rect 547342 117922 547398 117978
rect 546970 100294 547026 100350
rect 547094 100294 547150 100350
rect 547218 100294 547274 100350
rect 547342 100294 547398 100350
rect 546970 100170 547026 100226
rect 547094 100170 547150 100226
rect 547218 100170 547274 100226
rect 547342 100170 547398 100226
rect 546970 100046 547026 100102
rect 547094 100046 547150 100102
rect 547218 100046 547274 100102
rect 547342 100046 547398 100102
rect 546970 99922 547026 99978
rect 547094 99922 547150 99978
rect 547218 99922 547274 99978
rect 547342 99922 547398 99978
rect 546970 82294 547026 82350
rect 547094 82294 547150 82350
rect 547218 82294 547274 82350
rect 547342 82294 547398 82350
rect 546970 82170 547026 82226
rect 547094 82170 547150 82226
rect 547218 82170 547274 82226
rect 547342 82170 547398 82226
rect 546970 82046 547026 82102
rect 547094 82046 547150 82102
rect 547218 82046 547274 82102
rect 547342 82046 547398 82102
rect 546970 81922 547026 81978
rect 547094 81922 547150 81978
rect 547218 81922 547274 81978
rect 547342 81922 547398 81978
rect 546970 64294 547026 64350
rect 547094 64294 547150 64350
rect 547218 64294 547274 64350
rect 547342 64294 547398 64350
rect 546970 64170 547026 64226
rect 547094 64170 547150 64226
rect 547218 64170 547274 64226
rect 547342 64170 547398 64226
rect 546970 64046 547026 64102
rect 547094 64046 547150 64102
rect 547218 64046 547274 64102
rect 547342 64046 547398 64102
rect 546970 63922 547026 63978
rect 547094 63922 547150 63978
rect 547218 63922 547274 63978
rect 547342 63922 547398 63978
rect 546970 46294 547026 46350
rect 547094 46294 547150 46350
rect 547218 46294 547274 46350
rect 547342 46294 547398 46350
rect 546970 46170 547026 46226
rect 547094 46170 547150 46226
rect 547218 46170 547274 46226
rect 547342 46170 547398 46226
rect 546970 46046 547026 46102
rect 547094 46046 547150 46102
rect 547218 46046 547274 46102
rect 547342 46046 547398 46102
rect 546970 45922 547026 45978
rect 547094 45922 547150 45978
rect 547218 45922 547274 45978
rect 547342 45922 547398 45978
rect 546970 28294 547026 28350
rect 547094 28294 547150 28350
rect 547218 28294 547274 28350
rect 547342 28294 547398 28350
rect 546970 28170 547026 28226
rect 547094 28170 547150 28226
rect 547218 28170 547274 28226
rect 547342 28170 547398 28226
rect 546970 28046 547026 28102
rect 547094 28046 547150 28102
rect 547218 28046 547274 28102
rect 547342 28046 547398 28102
rect 546970 27922 547026 27978
rect 547094 27922 547150 27978
rect 547218 27922 547274 27978
rect 547342 27922 547398 27978
rect 546970 10294 547026 10350
rect 547094 10294 547150 10350
rect 547218 10294 547274 10350
rect 547342 10294 547398 10350
rect 546970 10170 547026 10226
rect 547094 10170 547150 10226
rect 547218 10170 547274 10226
rect 547342 10170 547398 10226
rect 546970 10046 547026 10102
rect 547094 10046 547150 10102
rect 547218 10046 547274 10102
rect 547342 10046 547398 10102
rect 546970 9922 547026 9978
rect 547094 9922 547150 9978
rect 547218 9922 547274 9978
rect 547342 9922 547398 9978
rect 561250 148294 561306 148350
rect 561374 148294 561430 148350
rect 561498 148294 561554 148350
rect 561622 148294 561678 148350
rect 561250 148170 561306 148226
rect 561374 148170 561430 148226
rect 561498 148170 561554 148226
rect 561622 148170 561678 148226
rect 561250 148046 561306 148102
rect 561374 148046 561430 148102
rect 561498 148046 561554 148102
rect 561622 148046 561678 148102
rect 561250 147922 561306 147978
rect 561374 147922 561430 147978
rect 561498 147922 561554 147978
rect 561622 147922 561678 147978
rect 561250 130294 561306 130350
rect 561374 130294 561430 130350
rect 561498 130294 561554 130350
rect 561622 130294 561678 130350
rect 561250 130170 561306 130226
rect 561374 130170 561430 130226
rect 561498 130170 561554 130226
rect 561622 130170 561678 130226
rect 561250 130046 561306 130102
rect 561374 130046 561430 130102
rect 561498 130046 561554 130102
rect 561622 130046 561678 130102
rect 561250 129922 561306 129978
rect 561374 129922 561430 129978
rect 561498 129922 561554 129978
rect 561622 129922 561678 129978
rect 561250 112294 561306 112350
rect 561374 112294 561430 112350
rect 561498 112294 561554 112350
rect 561622 112294 561678 112350
rect 561250 112170 561306 112226
rect 561374 112170 561430 112226
rect 561498 112170 561554 112226
rect 561622 112170 561678 112226
rect 561250 112046 561306 112102
rect 561374 112046 561430 112102
rect 561498 112046 561554 112102
rect 561622 112046 561678 112102
rect 561250 111922 561306 111978
rect 561374 111922 561430 111978
rect 561498 111922 561554 111978
rect 561622 111922 561678 111978
rect 555238 94294 555294 94350
rect 555362 94294 555418 94350
rect 555238 94170 555294 94226
rect 555362 94170 555418 94226
rect 555238 94046 555294 94102
rect 555362 94046 555418 94102
rect 555238 93922 555294 93978
rect 555362 93922 555418 93978
rect 561250 94294 561306 94350
rect 561374 94294 561430 94350
rect 561498 94294 561554 94350
rect 561622 94294 561678 94350
rect 561250 94170 561306 94226
rect 561374 94170 561430 94226
rect 561498 94170 561554 94226
rect 561622 94170 561678 94226
rect 561250 94046 561306 94102
rect 561374 94046 561430 94102
rect 561498 94046 561554 94102
rect 561622 94046 561678 94102
rect 561250 93922 561306 93978
rect 561374 93922 561430 93978
rect 561498 93922 561554 93978
rect 561622 93922 561678 93978
rect 555238 76294 555294 76350
rect 555362 76294 555418 76350
rect 555238 76170 555294 76226
rect 555362 76170 555418 76226
rect 555238 76046 555294 76102
rect 555362 76046 555418 76102
rect 555238 75922 555294 75978
rect 555362 75922 555418 75978
rect 561250 76294 561306 76350
rect 561374 76294 561430 76350
rect 561498 76294 561554 76350
rect 561622 76294 561678 76350
rect 561250 76170 561306 76226
rect 561374 76170 561430 76226
rect 561498 76170 561554 76226
rect 561622 76170 561678 76226
rect 561250 76046 561306 76102
rect 561374 76046 561430 76102
rect 561498 76046 561554 76102
rect 561622 76046 561678 76102
rect 561250 75922 561306 75978
rect 561374 75922 561430 75978
rect 561498 75922 561554 75978
rect 561622 75922 561678 75978
rect 561250 58294 561306 58350
rect 561374 58294 561430 58350
rect 561498 58294 561554 58350
rect 561622 58294 561678 58350
rect 561250 58170 561306 58226
rect 561374 58170 561430 58226
rect 561498 58170 561554 58226
rect 561622 58170 561678 58226
rect 561250 58046 561306 58102
rect 561374 58046 561430 58102
rect 561498 58046 561554 58102
rect 561622 58046 561678 58102
rect 561250 57922 561306 57978
rect 561374 57922 561430 57978
rect 561498 57922 561554 57978
rect 561622 57922 561678 57978
rect 561250 40294 561306 40350
rect 561374 40294 561430 40350
rect 561498 40294 561554 40350
rect 561622 40294 561678 40350
rect 561250 40170 561306 40226
rect 561374 40170 561430 40226
rect 561498 40170 561554 40226
rect 561622 40170 561678 40226
rect 561250 40046 561306 40102
rect 561374 40046 561430 40102
rect 561498 40046 561554 40102
rect 561622 40046 561678 40102
rect 561250 39922 561306 39978
rect 561374 39922 561430 39978
rect 561498 39922 561554 39978
rect 561622 39922 561678 39978
rect 561250 22294 561306 22350
rect 561374 22294 561430 22350
rect 561498 22294 561554 22350
rect 561622 22294 561678 22350
rect 561250 22170 561306 22226
rect 561374 22170 561430 22226
rect 561498 22170 561554 22226
rect 561622 22170 561678 22226
rect 561250 22046 561306 22102
rect 561374 22046 561430 22102
rect 561498 22046 561554 22102
rect 561622 22046 561678 22102
rect 561250 21922 561306 21978
rect 561374 21922 561430 21978
rect 561498 21922 561554 21978
rect 561622 21922 561678 21978
rect 561250 4294 561306 4350
rect 561374 4294 561430 4350
rect 561498 4294 561554 4350
rect 561622 4294 561678 4350
rect 561250 4170 561306 4226
rect 561374 4170 561430 4226
rect 561498 4170 561554 4226
rect 561622 4170 561678 4226
rect 561250 4046 561306 4102
rect 561374 4046 561430 4102
rect 561498 4046 561554 4102
rect 561622 4046 561678 4102
rect 561250 3922 561306 3978
rect 561374 3922 561430 3978
rect 561498 3922 561554 3978
rect 561622 3922 561678 3978
rect 546970 -1176 547026 -1120
rect 547094 -1176 547150 -1120
rect 547218 -1176 547274 -1120
rect 547342 -1176 547398 -1120
rect 546970 -1300 547026 -1244
rect 547094 -1300 547150 -1244
rect 547218 -1300 547274 -1244
rect 547342 -1300 547398 -1244
rect 546970 -1424 547026 -1368
rect 547094 -1424 547150 -1368
rect 547218 -1424 547274 -1368
rect 547342 -1424 547398 -1368
rect 546970 -1548 547026 -1492
rect 547094 -1548 547150 -1492
rect 547218 -1548 547274 -1492
rect 547342 -1548 547398 -1492
rect 564970 154294 565026 154350
rect 565094 154294 565150 154350
rect 565218 154294 565274 154350
rect 565342 154294 565398 154350
rect 564970 154170 565026 154226
rect 565094 154170 565150 154226
rect 565218 154170 565274 154226
rect 565342 154170 565398 154226
rect 564970 154046 565026 154102
rect 565094 154046 565150 154102
rect 565218 154046 565274 154102
rect 565342 154046 565398 154102
rect 564970 153922 565026 153978
rect 565094 153922 565150 153978
rect 565218 153922 565274 153978
rect 565342 153922 565398 153978
rect 564970 136294 565026 136350
rect 565094 136294 565150 136350
rect 565218 136294 565274 136350
rect 565342 136294 565398 136350
rect 564970 136170 565026 136226
rect 565094 136170 565150 136226
rect 565218 136170 565274 136226
rect 565342 136170 565398 136226
rect 564970 136046 565026 136102
rect 565094 136046 565150 136102
rect 565218 136046 565274 136102
rect 565342 136046 565398 136102
rect 564970 135922 565026 135978
rect 565094 135922 565150 135978
rect 565218 135922 565274 135978
rect 565342 135922 565398 135978
rect 564970 118294 565026 118350
rect 565094 118294 565150 118350
rect 565218 118294 565274 118350
rect 565342 118294 565398 118350
rect 564970 118170 565026 118226
rect 565094 118170 565150 118226
rect 565218 118170 565274 118226
rect 565342 118170 565398 118226
rect 564970 118046 565026 118102
rect 565094 118046 565150 118102
rect 565218 118046 565274 118102
rect 565342 118046 565398 118102
rect 564970 117922 565026 117978
rect 565094 117922 565150 117978
rect 565218 117922 565274 117978
rect 565342 117922 565398 117978
rect 564970 100294 565026 100350
rect 565094 100294 565150 100350
rect 565218 100294 565274 100350
rect 565342 100294 565398 100350
rect 564970 100170 565026 100226
rect 565094 100170 565150 100226
rect 565218 100170 565274 100226
rect 565342 100170 565398 100226
rect 564970 100046 565026 100102
rect 565094 100046 565150 100102
rect 565218 100046 565274 100102
rect 565342 100046 565398 100102
rect 564970 99922 565026 99978
rect 565094 99922 565150 99978
rect 565218 99922 565274 99978
rect 565342 99922 565398 99978
rect 564970 82294 565026 82350
rect 565094 82294 565150 82350
rect 565218 82294 565274 82350
rect 565342 82294 565398 82350
rect 564970 82170 565026 82226
rect 565094 82170 565150 82226
rect 565218 82170 565274 82226
rect 565342 82170 565398 82226
rect 564970 82046 565026 82102
rect 565094 82046 565150 82102
rect 565218 82046 565274 82102
rect 565342 82046 565398 82102
rect 564970 81922 565026 81978
rect 565094 81922 565150 81978
rect 565218 81922 565274 81978
rect 565342 81922 565398 81978
rect 564970 64294 565026 64350
rect 565094 64294 565150 64350
rect 565218 64294 565274 64350
rect 565342 64294 565398 64350
rect 564970 64170 565026 64226
rect 565094 64170 565150 64226
rect 565218 64170 565274 64226
rect 565342 64170 565398 64226
rect 564970 64046 565026 64102
rect 565094 64046 565150 64102
rect 565218 64046 565274 64102
rect 565342 64046 565398 64102
rect 564970 63922 565026 63978
rect 565094 63922 565150 63978
rect 565218 63922 565274 63978
rect 565342 63922 565398 63978
rect 564970 46294 565026 46350
rect 565094 46294 565150 46350
rect 565218 46294 565274 46350
rect 565342 46294 565398 46350
rect 564970 46170 565026 46226
rect 565094 46170 565150 46226
rect 565218 46170 565274 46226
rect 565342 46170 565398 46226
rect 564970 46046 565026 46102
rect 565094 46046 565150 46102
rect 565218 46046 565274 46102
rect 565342 46046 565398 46102
rect 564970 45922 565026 45978
rect 565094 45922 565150 45978
rect 565218 45922 565274 45978
rect 565342 45922 565398 45978
rect 564970 28294 565026 28350
rect 565094 28294 565150 28350
rect 565218 28294 565274 28350
rect 565342 28294 565398 28350
rect 564970 28170 565026 28226
rect 565094 28170 565150 28226
rect 565218 28170 565274 28226
rect 565342 28170 565398 28226
rect 564970 28046 565026 28102
rect 565094 28046 565150 28102
rect 565218 28046 565274 28102
rect 565342 28046 565398 28102
rect 564970 27922 565026 27978
rect 565094 27922 565150 27978
rect 565218 27922 565274 27978
rect 565342 27922 565398 27978
rect 564970 10294 565026 10350
rect 565094 10294 565150 10350
rect 565218 10294 565274 10350
rect 565342 10294 565398 10350
rect 564970 10170 565026 10226
rect 565094 10170 565150 10226
rect 565218 10170 565274 10226
rect 565342 10170 565398 10226
rect 564970 10046 565026 10102
rect 565094 10046 565150 10102
rect 565218 10046 565274 10102
rect 565342 10046 565398 10102
rect 564970 9922 565026 9978
rect 565094 9922 565150 9978
rect 565218 9922 565274 9978
rect 565342 9922 565398 9978
rect 561250 -216 561306 -160
rect 561374 -216 561430 -160
rect 561498 -216 561554 -160
rect 561622 -216 561678 -160
rect 561250 -340 561306 -284
rect 561374 -340 561430 -284
rect 561498 -340 561554 -284
rect 561622 -340 561678 -284
rect 561250 -464 561306 -408
rect 561374 -464 561430 -408
rect 561498 -464 561554 -408
rect 561622 -464 561678 -408
rect 561250 -588 561306 -532
rect 561374 -588 561430 -532
rect 561498 -588 561554 -532
rect 561622 -588 561678 -532
rect 564970 -1176 565026 -1120
rect 565094 -1176 565150 -1120
rect 565218 -1176 565274 -1120
rect 565342 -1176 565398 -1120
rect 564970 -1300 565026 -1244
rect 565094 -1300 565150 -1244
rect 565218 -1300 565274 -1244
rect 565342 -1300 565398 -1244
rect 564970 -1424 565026 -1368
rect 565094 -1424 565150 -1368
rect 565218 -1424 565274 -1368
rect 565342 -1424 565398 -1368
rect 564970 -1548 565026 -1492
rect 565094 -1548 565150 -1492
rect 565218 -1548 565274 -1492
rect 565342 -1548 565398 -1492
rect 579250 148294 579306 148350
rect 579374 148294 579430 148350
rect 579498 148294 579554 148350
rect 579622 148294 579678 148350
rect 579250 148170 579306 148226
rect 579374 148170 579430 148226
rect 579498 148170 579554 148226
rect 579622 148170 579678 148226
rect 579250 148046 579306 148102
rect 579374 148046 579430 148102
rect 579498 148046 579554 148102
rect 579622 148046 579678 148102
rect 579250 147922 579306 147978
rect 579374 147922 579430 147978
rect 579498 147922 579554 147978
rect 579622 147922 579678 147978
rect 579250 130294 579306 130350
rect 579374 130294 579430 130350
rect 579498 130294 579554 130350
rect 579622 130294 579678 130350
rect 579250 130170 579306 130226
rect 579374 130170 579430 130226
rect 579498 130170 579554 130226
rect 579622 130170 579678 130226
rect 579250 130046 579306 130102
rect 579374 130046 579430 130102
rect 579498 130046 579554 130102
rect 579622 130046 579678 130102
rect 579250 129922 579306 129978
rect 579374 129922 579430 129978
rect 579498 129922 579554 129978
rect 579622 129922 579678 129978
rect 579250 112294 579306 112350
rect 579374 112294 579430 112350
rect 579498 112294 579554 112350
rect 579622 112294 579678 112350
rect 579250 112170 579306 112226
rect 579374 112170 579430 112226
rect 579498 112170 579554 112226
rect 579622 112170 579678 112226
rect 579250 112046 579306 112102
rect 579374 112046 579430 112102
rect 579498 112046 579554 112102
rect 579622 112046 579678 112102
rect 579250 111922 579306 111978
rect 579374 111922 579430 111978
rect 579498 111922 579554 111978
rect 579622 111922 579678 111978
rect 579250 94294 579306 94350
rect 579374 94294 579430 94350
rect 579498 94294 579554 94350
rect 579622 94294 579678 94350
rect 579250 94170 579306 94226
rect 579374 94170 579430 94226
rect 579498 94170 579554 94226
rect 579622 94170 579678 94226
rect 579250 94046 579306 94102
rect 579374 94046 579430 94102
rect 579498 94046 579554 94102
rect 579622 94046 579678 94102
rect 579250 93922 579306 93978
rect 579374 93922 579430 93978
rect 579498 93922 579554 93978
rect 579622 93922 579678 93978
rect 579250 76294 579306 76350
rect 579374 76294 579430 76350
rect 579498 76294 579554 76350
rect 579622 76294 579678 76350
rect 579250 76170 579306 76226
rect 579374 76170 579430 76226
rect 579498 76170 579554 76226
rect 579622 76170 579678 76226
rect 579250 76046 579306 76102
rect 579374 76046 579430 76102
rect 579498 76046 579554 76102
rect 579622 76046 579678 76102
rect 579250 75922 579306 75978
rect 579374 75922 579430 75978
rect 579498 75922 579554 75978
rect 579622 75922 579678 75978
rect 579250 58294 579306 58350
rect 579374 58294 579430 58350
rect 579498 58294 579554 58350
rect 579622 58294 579678 58350
rect 579250 58170 579306 58226
rect 579374 58170 579430 58226
rect 579498 58170 579554 58226
rect 579622 58170 579678 58226
rect 579250 58046 579306 58102
rect 579374 58046 579430 58102
rect 579498 58046 579554 58102
rect 579622 58046 579678 58102
rect 579250 57922 579306 57978
rect 579374 57922 579430 57978
rect 579498 57922 579554 57978
rect 579622 57922 579678 57978
rect 579250 40294 579306 40350
rect 579374 40294 579430 40350
rect 579498 40294 579554 40350
rect 579622 40294 579678 40350
rect 579250 40170 579306 40226
rect 579374 40170 579430 40226
rect 579498 40170 579554 40226
rect 579622 40170 579678 40226
rect 579250 40046 579306 40102
rect 579374 40046 579430 40102
rect 579498 40046 579554 40102
rect 579622 40046 579678 40102
rect 579250 39922 579306 39978
rect 579374 39922 579430 39978
rect 579498 39922 579554 39978
rect 579622 39922 579678 39978
rect 579250 22294 579306 22350
rect 579374 22294 579430 22350
rect 579498 22294 579554 22350
rect 579622 22294 579678 22350
rect 579250 22170 579306 22226
rect 579374 22170 579430 22226
rect 579498 22170 579554 22226
rect 579622 22170 579678 22226
rect 579250 22046 579306 22102
rect 579374 22046 579430 22102
rect 579498 22046 579554 22102
rect 579622 22046 579678 22102
rect 579250 21922 579306 21978
rect 579374 21922 579430 21978
rect 579498 21922 579554 21978
rect 579622 21922 579678 21978
rect 579250 4294 579306 4350
rect 579374 4294 579430 4350
rect 579498 4294 579554 4350
rect 579622 4294 579678 4350
rect 579250 4170 579306 4226
rect 579374 4170 579430 4226
rect 579498 4170 579554 4226
rect 579622 4170 579678 4226
rect 579250 4046 579306 4102
rect 579374 4046 579430 4102
rect 579498 4046 579554 4102
rect 579622 4046 579678 4102
rect 579250 3922 579306 3978
rect 579374 3922 579430 3978
rect 579498 3922 579554 3978
rect 579622 3922 579678 3978
rect 579250 -216 579306 -160
rect 579374 -216 579430 -160
rect 579498 -216 579554 -160
rect 579622 -216 579678 -160
rect 579250 -340 579306 -284
rect 579374 -340 579430 -284
rect 579498 -340 579554 -284
rect 579622 -340 579678 -284
rect 579250 -464 579306 -408
rect 579374 -464 579430 -408
rect 579498 -464 579554 -408
rect 579622 -464 579678 -408
rect 579250 -588 579306 -532
rect 579374 -588 579430 -532
rect 579498 -588 579554 -532
rect 579622 -588 579678 -532
rect 582970 598116 583026 598172
rect 583094 598116 583150 598172
rect 583218 598116 583274 598172
rect 583342 598116 583398 598172
rect 582970 597992 583026 598048
rect 583094 597992 583150 598048
rect 583218 597992 583274 598048
rect 583342 597992 583398 598048
rect 582970 597868 583026 597924
rect 583094 597868 583150 597924
rect 583218 597868 583274 597924
rect 583342 597868 583398 597924
rect 582970 597744 583026 597800
rect 583094 597744 583150 597800
rect 583218 597744 583274 597800
rect 583342 597744 583398 597800
rect 597456 598116 597512 598172
rect 597580 598116 597636 598172
rect 597704 598116 597760 598172
rect 597828 598116 597884 598172
rect 597456 597992 597512 598048
rect 597580 597992 597636 598048
rect 597704 597992 597760 598048
rect 597828 597992 597884 598048
rect 597456 597868 597512 597924
rect 597580 597868 597636 597924
rect 597704 597868 597760 597924
rect 597828 597868 597884 597924
rect 597456 597744 597512 597800
rect 597580 597744 597636 597800
rect 597704 597744 597760 597800
rect 597828 597744 597884 597800
rect 582970 586294 583026 586350
rect 583094 586294 583150 586350
rect 583218 586294 583274 586350
rect 583342 586294 583398 586350
rect 582970 586170 583026 586226
rect 583094 586170 583150 586226
rect 583218 586170 583274 586226
rect 583342 586170 583398 586226
rect 582970 586046 583026 586102
rect 583094 586046 583150 586102
rect 583218 586046 583274 586102
rect 583342 586046 583398 586102
rect 582970 585922 583026 585978
rect 583094 585922 583150 585978
rect 583218 585922 583274 585978
rect 583342 585922 583398 585978
rect 582970 568294 583026 568350
rect 583094 568294 583150 568350
rect 583218 568294 583274 568350
rect 583342 568294 583398 568350
rect 582970 568170 583026 568226
rect 583094 568170 583150 568226
rect 583218 568170 583274 568226
rect 583342 568170 583398 568226
rect 582970 568046 583026 568102
rect 583094 568046 583150 568102
rect 583218 568046 583274 568102
rect 583342 568046 583398 568102
rect 582970 567922 583026 567978
rect 583094 567922 583150 567978
rect 583218 567922 583274 567978
rect 583342 567922 583398 567978
rect 582970 550294 583026 550350
rect 583094 550294 583150 550350
rect 583218 550294 583274 550350
rect 583342 550294 583398 550350
rect 582970 550170 583026 550226
rect 583094 550170 583150 550226
rect 583218 550170 583274 550226
rect 583342 550170 583398 550226
rect 582970 550046 583026 550102
rect 583094 550046 583150 550102
rect 583218 550046 583274 550102
rect 583342 550046 583398 550102
rect 582970 549922 583026 549978
rect 583094 549922 583150 549978
rect 583218 549922 583274 549978
rect 583342 549922 583398 549978
rect 582970 532294 583026 532350
rect 583094 532294 583150 532350
rect 583218 532294 583274 532350
rect 583342 532294 583398 532350
rect 582970 532170 583026 532226
rect 583094 532170 583150 532226
rect 583218 532170 583274 532226
rect 583342 532170 583398 532226
rect 582970 532046 583026 532102
rect 583094 532046 583150 532102
rect 583218 532046 583274 532102
rect 583342 532046 583398 532102
rect 582970 531922 583026 531978
rect 583094 531922 583150 531978
rect 583218 531922 583274 531978
rect 583342 531922 583398 531978
rect 582970 514294 583026 514350
rect 583094 514294 583150 514350
rect 583218 514294 583274 514350
rect 583342 514294 583398 514350
rect 582970 514170 583026 514226
rect 583094 514170 583150 514226
rect 583218 514170 583274 514226
rect 583342 514170 583398 514226
rect 582970 514046 583026 514102
rect 583094 514046 583150 514102
rect 583218 514046 583274 514102
rect 583342 514046 583398 514102
rect 582970 513922 583026 513978
rect 583094 513922 583150 513978
rect 583218 513922 583274 513978
rect 583342 513922 583398 513978
rect 582970 496294 583026 496350
rect 583094 496294 583150 496350
rect 583218 496294 583274 496350
rect 583342 496294 583398 496350
rect 582970 496170 583026 496226
rect 583094 496170 583150 496226
rect 583218 496170 583274 496226
rect 583342 496170 583398 496226
rect 582970 496046 583026 496102
rect 583094 496046 583150 496102
rect 583218 496046 583274 496102
rect 583342 496046 583398 496102
rect 582970 495922 583026 495978
rect 583094 495922 583150 495978
rect 583218 495922 583274 495978
rect 583342 495922 583398 495978
rect 582970 478294 583026 478350
rect 583094 478294 583150 478350
rect 583218 478294 583274 478350
rect 583342 478294 583398 478350
rect 582970 478170 583026 478226
rect 583094 478170 583150 478226
rect 583218 478170 583274 478226
rect 583342 478170 583398 478226
rect 582970 478046 583026 478102
rect 583094 478046 583150 478102
rect 583218 478046 583274 478102
rect 583342 478046 583398 478102
rect 582970 477922 583026 477978
rect 583094 477922 583150 477978
rect 583218 477922 583274 477978
rect 583342 477922 583398 477978
rect 582970 460294 583026 460350
rect 583094 460294 583150 460350
rect 583218 460294 583274 460350
rect 583342 460294 583398 460350
rect 582970 460170 583026 460226
rect 583094 460170 583150 460226
rect 583218 460170 583274 460226
rect 583342 460170 583398 460226
rect 582970 460046 583026 460102
rect 583094 460046 583150 460102
rect 583218 460046 583274 460102
rect 583342 460046 583398 460102
rect 582970 459922 583026 459978
rect 583094 459922 583150 459978
rect 583218 459922 583274 459978
rect 583342 459922 583398 459978
rect 582970 442294 583026 442350
rect 583094 442294 583150 442350
rect 583218 442294 583274 442350
rect 583342 442294 583398 442350
rect 582970 442170 583026 442226
rect 583094 442170 583150 442226
rect 583218 442170 583274 442226
rect 583342 442170 583398 442226
rect 582970 442046 583026 442102
rect 583094 442046 583150 442102
rect 583218 442046 583274 442102
rect 583342 442046 583398 442102
rect 582970 441922 583026 441978
rect 583094 441922 583150 441978
rect 583218 441922 583274 441978
rect 583342 441922 583398 441978
rect 582970 424294 583026 424350
rect 583094 424294 583150 424350
rect 583218 424294 583274 424350
rect 583342 424294 583398 424350
rect 582970 424170 583026 424226
rect 583094 424170 583150 424226
rect 583218 424170 583274 424226
rect 583342 424170 583398 424226
rect 582970 424046 583026 424102
rect 583094 424046 583150 424102
rect 583218 424046 583274 424102
rect 583342 424046 583398 424102
rect 582970 423922 583026 423978
rect 583094 423922 583150 423978
rect 583218 423922 583274 423978
rect 583342 423922 583398 423978
rect 582970 406294 583026 406350
rect 583094 406294 583150 406350
rect 583218 406294 583274 406350
rect 583342 406294 583398 406350
rect 582970 406170 583026 406226
rect 583094 406170 583150 406226
rect 583218 406170 583274 406226
rect 583342 406170 583398 406226
rect 582970 406046 583026 406102
rect 583094 406046 583150 406102
rect 583218 406046 583274 406102
rect 583342 406046 583398 406102
rect 582970 405922 583026 405978
rect 583094 405922 583150 405978
rect 583218 405922 583274 405978
rect 583342 405922 583398 405978
rect 582970 388294 583026 388350
rect 583094 388294 583150 388350
rect 583218 388294 583274 388350
rect 583342 388294 583398 388350
rect 582970 388170 583026 388226
rect 583094 388170 583150 388226
rect 583218 388170 583274 388226
rect 583342 388170 583398 388226
rect 582970 388046 583026 388102
rect 583094 388046 583150 388102
rect 583218 388046 583274 388102
rect 583342 388046 583398 388102
rect 582970 387922 583026 387978
rect 583094 387922 583150 387978
rect 583218 387922 583274 387978
rect 583342 387922 583398 387978
rect 582970 370294 583026 370350
rect 583094 370294 583150 370350
rect 583218 370294 583274 370350
rect 583342 370294 583398 370350
rect 582970 370170 583026 370226
rect 583094 370170 583150 370226
rect 583218 370170 583274 370226
rect 583342 370170 583398 370226
rect 582970 370046 583026 370102
rect 583094 370046 583150 370102
rect 583218 370046 583274 370102
rect 583342 370046 583398 370102
rect 582970 369922 583026 369978
rect 583094 369922 583150 369978
rect 583218 369922 583274 369978
rect 583342 369922 583398 369978
rect 582970 352294 583026 352350
rect 583094 352294 583150 352350
rect 583218 352294 583274 352350
rect 583342 352294 583398 352350
rect 582970 352170 583026 352226
rect 583094 352170 583150 352226
rect 583218 352170 583274 352226
rect 583342 352170 583398 352226
rect 582970 352046 583026 352102
rect 583094 352046 583150 352102
rect 583218 352046 583274 352102
rect 583342 352046 583398 352102
rect 582970 351922 583026 351978
rect 583094 351922 583150 351978
rect 583218 351922 583274 351978
rect 583342 351922 583398 351978
rect 582970 334294 583026 334350
rect 583094 334294 583150 334350
rect 583218 334294 583274 334350
rect 583342 334294 583398 334350
rect 582970 334170 583026 334226
rect 583094 334170 583150 334226
rect 583218 334170 583274 334226
rect 583342 334170 583398 334226
rect 582970 334046 583026 334102
rect 583094 334046 583150 334102
rect 583218 334046 583274 334102
rect 583342 334046 583398 334102
rect 582970 333922 583026 333978
rect 583094 333922 583150 333978
rect 583218 333922 583274 333978
rect 583342 333922 583398 333978
rect 582970 316294 583026 316350
rect 583094 316294 583150 316350
rect 583218 316294 583274 316350
rect 583342 316294 583398 316350
rect 582970 316170 583026 316226
rect 583094 316170 583150 316226
rect 583218 316170 583274 316226
rect 583342 316170 583398 316226
rect 582970 316046 583026 316102
rect 583094 316046 583150 316102
rect 583218 316046 583274 316102
rect 583342 316046 583398 316102
rect 582970 315922 583026 315978
rect 583094 315922 583150 315978
rect 583218 315922 583274 315978
rect 583342 315922 583398 315978
rect 582970 298294 583026 298350
rect 583094 298294 583150 298350
rect 583218 298294 583274 298350
rect 583342 298294 583398 298350
rect 582970 298170 583026 298226
rect 583094 298170 583150 298226
rect 583218 298170 583274 298226
rect 583342 298170 583398 298226
rect 582970 298046 583026 298102
rect 583094 298046 583150 298102
rect 583218 298046 583274 298102
rect 583342 298046 583398 298102
rect 582970 297922 583026 297978
rect 583094 297922 583150 297978
rect 583218 297922 583274 297978
rect 583342 297922 583398 297978
rect 582970 280294 583026 280350
rect 583094 280294 583150 280350
rect 583218 280294 583274 280350
rect 583342 280294 583398 280350
rect 582970 280170 583026 280226
rect 583094 280170 583150 280226
rect 583218 280170 583274 280226
rect 583342 280170 583398 280226
rect 582970 280046 583026 280102
rect 583094 280046 583150 280102
rect 583218 280046 583274 280102
rect 583342 280046 583398 280102
rect 582970 279922 583026 279978
rect 583094 279922 583150 279978
rect 583218 279922 583274 279978
rect 583342 279922 583398 279978
rect 582970 262294 583026 262350
rect 583094 262294 583150 262350
rect 583218 262294 583274 262350
rect 583342 262294 583398 262350
rect 582970 262170 583026 262226
rect 583094 262170 583150 262226
rect 583218 262170 583274 262226
rect 583342 262170 583398 262226
rect 582970 262046 583026 262102
rect 583094 262046 583150 262102
rect 583218 262046 583274 262102
rect 583342 262046 583398 262102
rect 582970 261922 583026 261978
rect 583094 261922 583150 261978
rect 583218 261922 583274 261978
rect 583342 261922 583398 261978
rect 582970 244294 583026 244350
rect 583094 244294 583150 244350
rect 583218 244294 583274 244350
rect 583342 244294 583398 244350
rect 582970 244170 583026 244226
rect 583094 244170 583150 244226
rect 583218 244170 583274 244226
rect 583342 244170 583398 244226
rect 582970 244046 583026 244102
rect 583094 244046 583150 244102
rect 583218 244046 583274 244102
rect 583342 244046 583398 244102
rect 582970 243922 583026 243978
rect 583094 243922 583150 243978
rect 583218 243922 583274 243978
rect 583342 243922 583398 243978
rect 582970 226294 583026 226350
rect 583094 226294 583150 226350
rect 583218 226294 583274 226350
rect 583342 226294 583398 226350
rect 582970 226170 583026 226226
rect 583094 226170 583150 226226
rect 583218 226170 583274 226226
rect 583342 226170 583398 226226
rect 582970 226046 583026 226102
rect 583094 226046 583150 226102
rect 583218 226046 583274 226102
rect 583342 226046 583398 226102
rect 582970 225922 583026 225978
rect 583094 225922 583150 225978
rect 583218 225922 583274 225978
rect 583342 225922 583398 225978
rect 582970 208294 583026 208350
rect 583094 208294 583150 208350
rect 583218 208294 583274 208350
rect 583342 208294 583398 208350
rect 582970 208170 583026 208226
rect 583094 208170 583150 208226
rect 583218 208170 583274 208226
rect 583342 208170 583398 208226
rect 582970 208046 583026 208102
rect 583094 208046 583150 208102
rect 583218 208046 583274 208102
rect 583342 208046 583398 208102
rect 582970 207922 583026 207978
rect 583094 207922 583150 207978
rect 583218 207922 583274 207978
rect 583342 207922 583398 207978
rect 582970 190294 583026 190350
rect 583094 190294 583150 190350
rect 583218 190294 583274 190350
rect 583342 190294 583398 190350
rect 582970 190170 583026 190226
rect 583094 190170 583150 190226
rect 583218 190170 583274 190226
rect 583342 190170 583398 190226
rect 582970 190046 583026 190102
rect 583094 190046 583150 190102
rect 583218 190046 583274 190102
rect 583342 190046 583398 190102
rect 582970 189922 583026 189978
rect 583094 189922 583150 189978
rect 583218 189922 583274 189978
rect 583342 189922 583398 189978
rect 582970 172294 583026 172350
rect 583094 172294 583150 172350
rect 583218 172294 583274 172350
rect 583342 172294 583398 172350
rect 582970 172170 583026 172226
rect 583094 172170 583150 172226
rect 583218 172170 583274 172226
rect 583342 172170 583398 172226
rect 582970 172046 583026 172102
rect 583094 172046 583150 172102
rect 583218 172046 583274 172102
rect 583342 172046 583398 172102
rect 582970 171922 583026 171978
rect 583094 171922 583150 171978
rect 583218 171922 583274 171978
rect 583342 171922 583398 171978
rect 582970 154294 583026 154350
rect 583094 154294 583150 154350
rect 583218 154294 583274 154350
rect 583342 154294 583398 154350
rect 582970 154170 583026 154226
rect 583094 154170 583150 154226
rect 583218 154170 583274 154226
rect 583342 154170 583398 154226
rect 582970 154046 583026 154102
rect 583094 154046 583150 154102
rect 583218 154046 583274 154102
rect 583342 154046 583398 154102
rect 582970 153922 583026 153978
rect 583094 153922 583150 153978
rect 583218 153922 583274 153978
rect 583342 153922 583398 153978
rect 582970 136294 583026 136350
rect 583094 136294 583150 136350
rect 583218 136294 583274 136350
rect 583342 136294 583398 136350
rect 582970 136170 583026 136226
rect 583094 136170 583150 136226
rect 583218 136170 583274 136226
rect 583342 136170 583398 136226
rect 582970 136046 583026 136102
rect 583094 136046 583150 136102
rect 583218 136046 583274 136102
rect 583342 136046 583398 136102
rect 582970 135922 583026 135978
rect 583094 135922 583150 135978
rect 583218 135922 583274 135978
rect 583342 135922 583398 135978
rect 582970 118294 583026 118350
rect 583094 118294 583150 118350
rect 583218 118294 583274 118350
rect 583342 118294 583398 118350
rect 582970 118170 583026 118226
rect 583094 118170 583150 118226
rect 583218 118170 583274 118226
rect 583342 118170 583398 118226
rect 582970 118046 583026 118102
rect 583094 118046 583150 118102
rect 583218 118046 583274 118102
rect 583342 118046 583398 118102
rect 582970 117922 583026 117978
rect 583094 117922 583150 117978
rect 583218 117922 583274 117978
rect 583342 117922 583398 117978
rect 582970 100294 583026 100350
rect 583094 100294 583150 100350
rect 583218 100294 583274 100350
rect 583342 100294 583398 100350
rect 582970 100170 583026 100226
rect 583094 100170 583150 100226
rect 583218 100170 583274 100226
rect 583342 100170 583398 100226
rect 582970 100046 583026 100102
rect 583094 100046 583150 100102
rect 583218 100046 583274 100102
rect 583342 100046 583398 100102
rect 582970 99922 583026 99978
rect 583094 99922 583150 99978
rect 583218 99922 583274 99978
rect 583342 99922 583398 99978
rect 582970 82294 583026 82350
rect 583094 82294 583150 82350
rect 583218 82294 583274 82350
rect 583342 82294 583398 82350
rect 582970 82170 583026 82226
rect 583094 82170 583150 82226
rect 583218 82170 583274 82226
rect 583342 82170 583398 82226
rect 582970 82046 583026 82102
rect 583094 82046 583150 82102
rect 583218 82046 583274 82102
rect 583342 82046 583398 82102
rect 582970 81922 583026 81978
rect 583094 81922 583150 81978
rect 583218 81922 583274 81978
rect 583342 81922 583398 81978
rect 582970 64294 583026 64350
rect 583094 64294 583150 64350
rect 583218 64294 583274 64350
rect 583342 64294 583398 64350
rect 582970 64170 583026 64226
rect 583094 64170 583150 64226
rect 583218 64170 583274 64226
rect 583342 64170 583398 64226
rect 582970 64046 583026 64102
rect 583094 64046 583150 64102
rect 583218 64046 583274 64102
rect 583342 64046 583398 64102
rect 582970 63922 583026 63978
rect 583094 63922 583150 63978
rect 583218 63922 583274 63978
rect 583342 63922 583398 63978
rect 582970 46294 583026 46350
rect 583094 46294 583150 46350
rect 583218 46294 583274 46350
rect 583342 46294 583398 46350
rect 582970 46170 583026 46226
rect 583094 46170 583150 46226
rect 583218 46170 583274 46226
rect 583342 46170 583398 46226
rect 582970 46046 583026 46102
rect 583094 46046 583150 46102
rect 583218 46046 583274 46102
rect 583342 46046 583398 46102
rect 582970 45922 583026 45978
rect 583094 45922 583150 45978
rect 583218 45922 583274 45978
rect 583342 45922 583398 45978
rect 582970 28294 583026 28350
rect 583094 28294 583150 28350
rect 583218 28294 583274 28350
rect 583342 28294 583398 28350
rect 582970 28170 583026 28226
rect 583094 28170 583150 28226
rect 583218 28170 583274 28226
rect 583342 28170 583398 28226
rect 582970 28046 583026 28102
rect 583094 28046 583150 28102
rect 583218 28046 583274 28102
rect 583342 28046 583398 28102
rect 582970 27922 583026 27978
rect 583094 27922 583150 27978
rect 583218 27922 583274 27978
rect 583342 27922 583398 27978
rect 582970 10294 583026 10350
rect 583094 10294 583150 10350
rect 583218 10294 583274 10350
rect 583342 10294 583398 10350
rect 582970 10170 583026 10226
rect 583094 10170 583150 10226
rect 583218 10170 583274 10226
rect 583342 10170 583398 10226
rect 582970 10046 583026 10102
rect 583094 10046 583150 10102
rect 583218 10046 583274 10102
rect 583342 10046 583398 10102
rect 582970 9922 583026 9978
rect 583094 9922 583150 9978
rect 583218 9922 583274 9978
rect 583342 9922 583398 9978
rect 596496 597156 596552 597212
rect 596620 597156 596676 597212
rect 596744 597156 596800 597212
rect 596868 597156 596924 597212
rect 596496 597032 596552 597088
rect 596620 597032 596676 597088
rect 596744 597032 596800 597088
rect 596868 597032 596924 597088
rect 596496 596908 596552 596964
rect 596620 596908 596676 596964
rect 596744 596908 596800 596964
rect 596868 596908 596924 596964
rect 596496 596784 596552 596840
rect 596620 596784 596676 596840
rect 596744 596784 596800 596840
rect 596868 596784 596924 596840
rect 596496 580294 596552 580350
rect 596620 580294 596676 580350
rect 596744 580294 596800 580350
rect 596868 580294 596924 580350
rect 596496 580170 596552 580226
rect 596620 580170 596676 580226
rect 596744 580170 596800 580226
rect 596868 580170 596924 580226
rect 596496 580046 596552 580102
rect 596620 580046 596676 580102
rect 596744 580046 596800 580102
rect 596868 580046 596924 580102
rect 596496 579922 596552 579978
rect 596620 579922 596676 579978
rect 596744 579922 596800 579978
rect 596868 579922 596924 579978
rect 596496 562294 596552 562350
rect 596620 562294 596676 562350
rect 596744 562294 596800 562350
rect 596868 562294 596924 562350
rect 596496 562170 596552 562226
rect 596620 562170 596676 562226
rect 596744 562170 596800 562226
rect 596868 562170 596924 562226
rect 596496 562046 596552 562102
rect 596620 562046 596676 562102
rect 596744 562046 596800 562102
rect 596868 562046 596924 562102
rect 596496 561922 596552 561978
rect 596620 561922 596676 561978
rect 596744 561922 596800 561978
rect 596868 561922 596924 561978
rect 596496 544294 596552 544350
rect 596620 544294 596676 544350
rect 596744 544294 596800 544350
rect 596868 544294 596924 544350
rect 596496 544170 596552 544226
rect 596620 544170 596676 544226
rect 596744 544170 596800 544226
rect 596868 544170 596924 544226
rect 596496 544046 596552 544102
rect 596620 544046 596676 544102
rect 596744 544046 596800 544102
rect 596868 544046 596924 544102
rect 596496 543922 596552 543978
rect 596620 543922 596676 543978
rect 596744 543922 596800 543978
rect 596868 543922 596924 543978
rect 596496 526294 596552 526350
rect 596620 526294 596676 526350
rect 596744 526294 596800 526350
rect 596868 526294 596924 526350
rect 596496 526170 596552 526226
rect 596620 526170 596676 526226
rect 596744 526170 596800 526226
rect 596868 526170 596924 526226
rect 596496 526046 596552 526102
rect 596620 526046 596676 526102
rect 596744 526046 596800 526102
rect 596868 526046 596924 526102
rect 596496 525922 596552 525978
rect 596620 525922 596676 525978
rect 596744 525922 596800 525978
rect 596868 525922 596924 525978
rect 596496 508294 596552 508350
rect 596620 508294 596676 508350
rect 596744 508294 596800 508350
rect 596868 508294 596924 508350
rect 596496 508170 596552 508226
rect 596620 508170 596676 508226
rect 596744 508170 596800 508226
rect 596868 508170 596924 508226
rect 596496 508046 596552 508102
rect 596620 508046 596676 508102
rect 596744 508046 596800 508102
rect 596868 508046 596924 508102
rect 596496 507922 596552 507978
rect 596620 507922 596676 507978
rect 596744 507922 596800 507978
rect 596868 507922 596924 507978
rect 596496 490294 596552 490350
rect 596620 490294 596676 490350
rect 596744 490294 596800 490350
rect 596868 490294 596924 490350
rect 596496 490170 596552 490226
rect 596620 490170 596676 490226
rect 596744 490170 596800 490226
rect 596868 490170 596924 490226
rect 596496 490046 596552 490102
rect 596620 490046 596676 490102
rect 596744 490046 596800 490102
rect 596868 490046 596924 490102
rect 596496 489922 596552 489978
rect 596620 489922 596676 489978
rect 596744 489922 596800 489978
rect 596868 489922 596924 489978
rect 596496 472294 596552 472350
rect 596620 472294 596676 472350
rect 596744 472294 596800 472350
rect 596868 472294 596924 472350
rect 596496 472170 596552 472226
rect 596620 472170 596676 472226
rect 596744 472170 596800 472226
rect 596868 472170 596924 472226
rect 596496 472046 596552 472102
rect 596620 472046 596676 472102
rect 596744 472046 596800 472102
rect 596868 472046 596924 472102
rect 596496 471922 596552 471978
rect 596620 471922 596676 471978
rect 596744 471922 596800 471978
rect 596868 471922 596924 471978
rect 596496 454294 596552 454350
rect 596620 454294 596676 454350
rect 596744 454294 596800 454350
rect 596868 454294 596924 454350
rect 596496 454170 596552 454226
rect 596620 454170 596676 454226
rect 596744 454170 596800 454226
rect 596868 454170 596924 454226
rect 596496 454046 596552 454102
rect 596620 454046 596676 454102
rect 596744 454046 596800 454102
rect 596868 454046 596924 454102
rect 596496 453922 596552 453978
rect 596620 453922 596676 453978
rect 596744 453922 596800 453978
rect 596868 453922 596924 453978
rect 596496 436294 596552 436350
rect 596620 436294 596676 436350
rect 596744 436294 596800 436350
rect 596868 436294 596924 436350
rect 596496 436170 596552 436226
rect 596620 436170 596676 436226
rect 596744 436170 596800 436226
rect 596868 436170 596924 436226
rect 596496 436046 596552 436102
rect 596620 436046 596676 436102
rect 596744 436046 596800 436102
rect 596868 436046 596924 436102
rect 596496 435922 596552 435978
rect 596620 435922 596676 435978
rect 596744 435922 596800 435978
rect 596868 435922 596924 435978
rect 596496 418294 596552 418350
rect 596620 418294 596676 418350
rect 596744 418294 596800 418350
rect 596868 418294 596924 418350
rect 596496 418170 596552 418226
rect 596620 418170 596676 418226
rect 596744 418170 596800 418226
rect 596868 418170 596924 418226
rect 596496 418046 596552 418102
rect 596620 418046 596676 418102
rect 596744 418046 596800 418102
rect 596868 418046 596924 418102
rect 596496 417922 596552 417978
rect 596620 417922 596676 417978
rect 596744 417922 596800 417978
rect 596868 417922 596924 417978
rect 596496 400294 596552 400350
rect 596620 400294 596676 400350
rect 596744 400294 596800 400350
rect 596868 400294 596924 400350
rect 596496 400170 596552 400226
rect 596620 400170 596676 400226
rect 596744 400170 596800 400226
rect 596868 400170 596924 400226
rect 596496 400046 596552 400102
rect 596620 400046 596676 400102
rect 596744 400046 596800 400102
rect 596868 400046 596924 400102
rect 596496 399922 596552 399978
rect 596620 399922 596676 399978
rect 596744 399922 596800 399978
rect 596868 399922 596924 399978
rect 596496 382294 596552 382350
rect 596620 382294 596676 382350
rect 596744 382294 596800 382350
rect 596868 382294 596924 382350
rect 596496 382170 596552 382226
rect 596620 382170 596676 382226
rect 596744 382170 596800 382226
rect 596868 382170 596924 382226
rect 596496 382046 596552 382102
rect 596620 382046 596676 382102
rect 596744 382046 596800 382102
rect 596868 382046 596924 382102
rect 596496 381922 596552 381978
rect 596620 381922 596676 381978
rect 596744 381922 596800 381978
rect 596868 381922 596924 381978
rect 596496 364294 596552 364350
rect 596620 364294 596676 364350
rect 596744 364294 596800 364350
rect 596868 364294 596924 364350
rect 596496 364170 596552 364226
rect 596620 364170 596676 364226
rect 596744 364170 596800 364226
rect 596868 364170 596924 364226
rect 596496 364046 596552 364102
rect 596620 364046 596676 364102
rect 596744 364046 596800 364102
rect 596868 364046 596924 364102
rect 596496 363922 596552 363978
rect 596620 363922 596676 363978
rect 596744 363922 596800 363978
rect 596868 363922 596924 363978
rect 596496 346294 596552 346350
rect 596620 346294 596676 346350
rect 596744 346294 596800 346350
rect 596868 346294 596924 346350
rect 596496 346170 596552 346226
rect 596620 346170 596676 346226
rect 596744 346170 596800 346226
rect 596868 346170 596924 346226
rect 596496 346046 596552 346102
rect 596620 346046 596676 346102
rect 596744 346046 596800 346102
rect 596868 346046 596924 346102
rect 596496 345922 596552 345978
rect 596620 345922 596676 345978
rect 596744 345922 596800 345978
rect 596868 345922 596924 345978
rect 596496 328294 596552 328350
rect 596620 328294 596676 328350
rect 596744 328294 596800 328350
rect 596868 328294 596924 328350
rect 596496 328170 596552 328226
rect 596620 328170 596676 328226
rect 596744 328170 596800 328226
rect 596868 328170 596924 328226
rect 596496 328046 596552 328102
rect 596620 328046 596676 328102
rect 596744 328046 596800 328102
rect 596868 328046 596924 328102
rect 596496 327922 596552 327978
rect 596620 327922 596676 327978
rect 596744 327922 596800 327978
rect 596868 327922 596924 327978
rect 596496 310294 596552 310350
rect 596620 310294 596676 310350
rect 596744 310294 596800 310350
rect 596868 310294 596924 310350
rect 596496 310170 596552 310226
rect 596620 310170 596676 310226
rect 596744 310170 596800 310226
rect 596868 310170 596924 310226
rect 596496 310046 596552 310102
rect 596620 310046 596676 310102
rect 596744 310046 596800 310102
rect 596868 310046 596924 310102
rect 596496 309922 596552 309978
rect 596620 309922 596676 309978
rect 596744 309922 596800 309978
rect 596868 309922 596924 309978
rect 596496 292294 596552 292350
rect 596620 292294 596676 292350
rect 596744 292294 596800 292350
rect 596868 292294 596924 292350
rect 596496 292170 596552 292226
rect 596620 292170 596676 292226
rect 596744 292170 596800 292226
rect 596868 292170 596924 292226
rect 596496 292046 596552 292102
rect 596620 292046 596676 292102
rect 596744 292046 596800 292102
rect 596868 292046 596924 292102
rect 596496 291922 596552 291978
rect 596620 291922 596676 291978
rect 596744 291922 596800 291978
rect 596868 291922 596924 291978
rect 596496 274294 596552 274350
rect 596620 274294 596676 274350
rect 596744 274294 596800 274350
rect 596868 274294 596924 274350
rect 596496 274170 596552 274226
rect 596620 274170 596676 274226
rect 596744 274170 596800 274226
rect 596868 274170 596924 274226
rect 596496 274046 596552 274102
rect 596620 274046 596676 274102
rect 596744 274046 596800 274102
rect 596868 274046 596924 274102
rect 596496 273922 596552 273978
rect 596620 273922 596676 273978
rect 596744 273922 596800 273978
rect 596868 273922 596924 273978
rect 596496 256294 596552 256350
rect 596620 256294 596676 256350
rect 596744 256294 596800 256350
rect 596868 256294 596924 256350
rect 596496 256170 596552 256226
rect 596620 256170 596676 256226
rect 596744 256170 596800 256226
rect 596868 256170 596924 256226
rect 596496 256046 596552 256102
rect 596620 256046 596676 256102
rect 596744 256046 596800 256102
rect 596868 256046 596924 256102
rect 596496 255922 596552 255978
rect 596620 255922 596676 255978
rect 596744 255922 596800 255978
rect 596868 255922 596924 255978
rect 596496 238294 596552 238350
rect 596620 238294 596676 238350
rect 596744 238294 596800 238350
rect 596868 238294 596924 238350
rect 596496 238170 596552 238226
rect 596620 238170 596676 238226
rect 596744 238170 596800 238226
rect 596868 238170 596924 238226
rect 596496 238046 596552 238102
rect 596620 238046 596676 238102
rect 596744 238046 596800 238102
rect 596868 238046 596924 238102
rect 596496 237922 596552 237978
rect 596620 237922 596676 237978
rect 596744 237922 596800 237978
rect 596868 237922 596924 237978
rect 596496 220294 596552 220350
rect 596620 220294 596676 220350
rect 596744 220294 596800 220350
rect 596868 220294 596924 220350
rect 596496 220170 596552 220226
rect 596620 220170 596676 220226
rect 596744 220170 596800 220226
rect 596868 220170 596924 220226
rect 596496 220046 596552 220102
rect 596620 220046 596676 220102
rect 596744 220046 596800 220102
rect 596868 220046 596924 220102
rect 596496 219922 596552 219978
rect 596620 219922 596676 219978
rect 596744 219922 596800 219978
rect 596868 219922 596924 219978
rect 596496 202294 596552 202350
rect 596620 202294 596676 202350
rect 596744 202294 596800 202350
rect 596868 202294 596924 202350
rect 596496 202170 596552 202226
rect 596620 202170 596676 202226
rect 596744 202170 596800 202226
rect 596868 202170 596924 202226
rect 596496 202046 596552 202102
rect 596620 202046 596676 202102
rect 596744 202046 596800 202102
rect 596868 202046 596924 202102
rect 596496 201922 596552 201978
rect 596620 201922 596676 201978
rect 596744 201922 596800 201978
rect 596868 201922 596924 201978
rect 596496 184294 596552 184350
rect 596620 184294 596676 184350
rect 596744 184294 596800 184350
rect 596868 184294 596924 184350
rect 596496 184170 596552 184226
rect 596620 184170 596676 184226
rect 596744 184170 596800 184226
rect 596868 184170 596924 184226
rect 596496 184046 596552 184102
rect 596620 184046 596676 184102
rect 596744 184046 596800 184102
rect 596868 184046 596924 184102
rect 596496 183922 596552 183978
rect 596620 183922 596676 183978
rect 596744 183922 596800 183978
rect 596868 183922 596924 183978
rect 596496 166294 596552 166350
rect 596620 166294 596676 166350
rect 596744 166294 596800 166350
rect 596868 166294 596924 166350
rect 596496 166170 596552 166226
rect 596620 166170 596676 166226
rect 596744 166170 596800 166226
rect 596868 166170 596924 166226
rect 596496 166046 596552 166102
rect 596620 166046 596676 166102
rect 596744 166046 596800 166102
rect 596868 166046 596924 166102
rect 596496 165922 596552 165978
rect 596620 165922 596676 165978
rect 596744 165922 596800 165978
rect 596868 165922 596924 165978
rect 596496 148294 596552 148350
rect 596620 148294 596676 148350
rect 596744 148294 596800 148350
rect 596868 148294 596924 148350
rect 596496 148170 596552 148226
rect 596620 148170 596676 148226
rect 596744 148170 596800 148226
rect 596868 148170 596924 148226
rect 596496 148046 596552 148102
rect 596620 148046 596676 148102
rect 596744 148046 596800 148102
rect 596868 148046 596924 148102
rect 596496 147922 596552 147978
rect 596620 147922 596676 147978
rect 596744 147922 596800 147978
rect 596868 147922 596924 147978
rect 596496 130294 596552 130350
rect 596620 130294 596676 130350
rect 596744 130294 596800 130350
rect 596868 130294 596924 130350
rect 596496 130170 596552 130226
rect 596620 130170 596676 130226
rect 596744 130170 596800 130226
rect 596868 130170 596924 130226
rect 596496 130046 596552 130102
rect 596620 130046 596676 130102
rect 596744 130046 596800 130102
rect 596868 130046 596924 130102
rect 596496 129922 596552 129978
rect 596620 129922 596676 129978
rect 596744 129922 596800 129978
rect 596868 129922 596924 129978
rect 596496 112294 596552 112350
rect 596620 112294 596676 112350
rect 596744 112294 596800 112350
rect 596868 112294 596924 112350
rect 596496 112170 596552 112226
rect 596620 112170 596676 112226
rect 596744 112170 596800 112226
rect 596868 112170 596924 112226
rect 596496 112046 596552 112102
rect 596620 112046 596676 112102
rect 596744 112046 596800 112102
rect 596868 112046 596924 112102
rect 596496 111922 596552 111978
rect 596620 111922 596676 111978
rect 596744 111922 596800 111978
rect 596868 111922 596924 111978
rect 596496 94294 596552 94350
rect 596620 94294 596676 94350
rect 596744 94294 596800 94350
rect 596868 94294 596924 94350
rect 596496 94170 596552 94226
rect 596620 94170 596676 94226
rect 596744 94170 596800 94226
rect 596868 94170 596924 94226
rect 596496 94046 596552 94102
rect 596620 94046 596676 94102
rect 596744 94046 596800 94102
rect 596868 94046 596924 94102
rect 596496 93922 596552 93978
rect 596620 93922 596676 93978
rect 596744 93922 596800 93978
rect 596868 93922 596924 93978
rect 596496 76294 596552 76350
rect 596620 76294 596676 76350
rect 596744 76294 596800 76350
rect 596868 76294 596924 76350
rect 596496 76170 596552 76226
rect 596620 76170 596676 76226
rect 596744 76170 596800 76226
rect 596868 76170 596924 76226
rect 596496 76046 596552 76102
rect 596620 76046 596676 76102
rect 596744 76046 596800 76102
rect 596868 76046 596924 76102
rect 596496 75922 596552 75978
rect 596620 75922 596676 75978
rect 596744 75922 596800 75978
rect 596868 75922 596924 75978
rect 596496 58294 596552 58350
rect 596620 58294 596676 58350
rect 596744 58294 596800 58350
rect 596868 58294 596924 58350
rect 596496 58170 596552 58226
rect 596620 58170 596676 58226
rect 596744 58170 596800 58226
rect 596868 58170 596924 58226
rect 596496 58046 596552 58102
rect 596620 58046 596676 58102
rect 596744 58046 596800 58102
rect 596868 58046 596924 58102
rect 596496 57922 596552 57978
rect 596620 57922 596676 57978
rect 596744 57922 596800 57978
rect 596868 57922 596924 57978
rect 596496 40294 596552 40350
rect 596620 40294 596676 40350
rect 596744 40294 596800 40350
rect 596868 40294 596924 40350
rect 596496 40170 596552 40226
rect 596620 40170 596676 40226
rect 596744 40170 596800 40226
rect 596868 40170 596924 40226
rect 596496 40046 596552 40102
rect 596620 40046 596676 40102
rect 596744 40046 596800 40102
rect 596868 40046 596924 40102
rect 596496 39922 596552 39978
rect 596620 39922 596676 39978
rect 596744 39922 596800 39978
rect 596868 39922 596924 39978
rect 596496 22294 596552 22350
rect 596620 22294 596676 22350
rect 596744 22294 596800 22350
rect 596868 22294 596924 22350
rect 596496 22170 596552 22226
rect 596620 22170 596676 22226
rect 596744 22170 596800 22226
rect 596868 22170 596924 22226
rect 596496 22046 596552 22102
rect 596620 22046 596676 22102
rect 596744 22046 596800 22102
rect 596868 22046 596924 22102
rect 596496 21922 596552 21978
rect 596620 21922 596676 21978
rect 596744 21922 596800 21978
rect 596868 21922 596924 21978
rect 596496 4294 596552 4350
rect 596620 4294 596676 4350
rect 596744 4294 596800 4350
rect 596868 4294 596924 4350
rect 596496 4170 596552 4226
rect 596620 4170 596676 4226
rect 596744 4170 596800 4226
rect 596868 4170 596924 4226
rect 596496 4046 596552 4102
rect 596620 4046 596676 4102
rect 596744 4046 596800 4102
rect 596868 4046 596924 4102
rect 596496 3922 596552 3978
rect 596620 3922 596676 3978
rect 596744 3922 596800 3978
rect 596868 3922 596924 3978
rect 596496 -216 596552 -160
rect 596620 -216 596676 -160
rect 596744 -216 596800 -160
rect 596868 -216 596924 -160
rect 596496 -340 596552 -284
rect 596620 -340 596676 -284
rect 596744 -340 596800 -284
rect 596868 -340 596924 -284
rect 596496 -464 596552 -408
rect 596620 -464 596676 -408
rect 596744 -464 596800 -408
rect 596868 -464 596924 -408
rect 596496 -588 596552 -532
rect 596620 -588 596676 -532
rect 596744 -588 596800 -532
rect 596868 -588 596924 -532
rect 597456 586294 597512 586350
rect 597580 586294 597636 586350
rect 597704 586294 597760 586350
rect 597828 586294 597884 586350
rect 597456 586170 597512 586226
rect 597580 586170 597636 586226
rect 597704 586170 597760 586226
rect 597828 586170 597884 586226
rect 597456 586046 597512 586102
rect 597580 586046 597636 586102
rect 597704 586046 597760 586102
rect 597828 586046 597884 586102
rect 597456 585922 597512 585978
rect 597580 585922 597636 585978
rect 597704 585922 597760 585978
rect 597828 585922 597884 585978
rect 597456 568294 597512 568350
rect 597580 568294 597636 568350
rect 597704 568294 597760 568350
rect 597828 568294 597884 568350
rect 597456 568170 597512 568226
rect 597580 568170 597636 568226
rect 597704 568170 597760 568226
rect 597828 568170 597884 568226
rect 597456 568046 597512 568102
rect 597580 568046 597636 568102
rect 597704 568046 597760 568102
rect 597828 568046 597884 568102
rect 597456 567922 597512 567978
rect 597580 567922 597636 567978
rect 597704 567922 597760 567978
rect 597828 567922 597884 567978
rect 597456 550294 597512 550350
rect 597580 550294 597636 550350
rect 597704 550294 597760 550350
rect 597828 550294 597884 550350
rect 597456 550170 597512 550226
rect 597580 550170 597636 550226
rect 597704 550170 597760 550226
rect 597828 550170 597884 550226
rect 597456 550046 597512 550102
rect 597580 550046 597636 550102
rect 597704 550046 597760 550102
rect 597828 550046 597884 550102
rect 597456 549922 597512 549978
rect 597580 549922 597636 549978
rect 597704 549922 597760 549978
rect 597828 549922 597884 549978
rect 597456 532294 597512 532350
rect 597580 532294 597636 532350
rect 597704 532294 597760 532350
rect 597828 532294 597884 532350
rect 597456 532170 597512 532226
rect 597580 532170 597636 532226
rect 597704 532170 597760 532226
rect 597828 532170 597884 532226
rect 597456 532046 597512 532102
rect 597580 532046 597636 532102
rect 597704 532046 597760 532102
rect 597828 532046 597884 532102
rect 597456 531922 597512 531978
rect 597580 531922 597636 531978
rect 597704 531922 597760 531978
rect 597828 531922 597884 531978
rect 597456 514294 597512 514350
rect 597580 514294 597636 514350
rect 597704 514294 597760 514350
rect 597828 514294 597884 514350
rect 597456 514170 597512 514226
rect 597580 514170 597636 514226
rect 597704 514170 597760 514226
rect 597828 514170 597884 514226
rect 597456 514046 597512 514102
rect 597580 514046 597636 514102
rect 597704 514046 597760 514102
rect 597828 514046 597884 514102
rect 597456 513922 597512 513978
rect 597580 513922 597636 513978
rect 597704 513922 597760 513978
rect 597828 513922 597884 513978
rect 597456 496294 597512 496350
rect 597580 496294 597636 496350
rect 597704 496294 597760 496350
rect 597828 496294 597884 496350
rect 597456 496170 597512 496226
rect 597580 496170 597636 496226
rect 597704 496170 597760 496226
rect 597828 496170 597884 496226
rect 597456 496046 597512 496102
rect 597580 496046 597636 496102
rect 597704 496046 597760 496102
rect 597828 496046 597884 496102
rect 597456 495922 597512 495978
rect 597580 495922 597636 495978
rect 597704 495922 597760 495978
rect 597828 495922 597884 495978
rect 597456 478294 597512 478350
rect 597580 478294 597636 478350
rect 597704 478294 597760 478350
rect 597828 478294 597884 478350
rect 597456 478170 597512 478226
rect 597580 478170 597636 478226
rect 597704 478170 597760 478226
rect 597828 478170 597884 478226
rect 597456 478046 597512 478102
rect 597580 478046 597636 478102
rect 597704 478046 597760 478102
rect 597828 478046 597884 478102
rect 597456 477922 597512 477978
rect 597580 477922 597636 477978
rect 597704 477922 597760 477978
rect 597828 477922 597884 477978
rect 597456 460294 597512 460350
rect 597580 460294 597636 460350
rect 597704 460294 597760 460350
rect 597828 460294 597884 460350
rect 597456 460170 597512 460226
rect 597580 460170 597636 460226
rect 597704 460170 597760 460226
rect 597828 460170 597884 460226
rect 597456 460046 597512 460102
rect 597580 460046 597636 460102
rect 597704 460046 597760 460102
rect 597828 460046 597884 460102
rect 597456 459922 597512 459978
rect 597580 459922 597636 459978
rect 597704 459922 597760 459978
rect 597828 459922 597884 459978
rect 597456 442294 597512 442350
rect 597580 442294 597636 442350
rect 597704 442294 597760 442350
rect 597828 442294 597884 442350
rect 597456 442170 597512 442226
rect 597580 442170 597636 442226
rect 597704 442170 597760 442226
rect 597828 442170 597884 442226
rect 597456 442046 597512 442102
rect 597580 442046 597636 442102
rect 597704 442046 597760 442102
rect 597828 442046 597884 442102
rect 597456 441922 597512 441978
rect 597580 441922 597636 441978
rect 597704 441922 597760 441978
rect 597828 441922 597884 441978
rect 597456 424294 597512 424350
rect 597580 424294 597636 424350
rect 597704 424294 597760 424350
rect 597828 424294 597884 424350
rect 597456 424170 597512 424226
rect 597580 424170 597636 424226
rect 597704 424170 597760 424226
rect 597828 424170 597884 424226
rect 597456 424046 597512 424102
rect 597580 424046 597636 424102
rect 597704 424046 597760 424102
rect 597828 424046 597884 424102
rect 597456 423922 597512 423978
rect 597580 423922 597636 423978
rect 597704 423922 597760 423978
rect 597828 423922 597884 423978
rect 597456 406294 597512 406350
rect 597580 406294 597636 406350
rect 597704 406294 597760 406350
rect 597828 406294 597884 406350
rect 597456 406170 597512 406226
rect 597580 406170 597636 406226
rect 597704 406170 597760 406226
rect 597828 406170 597884 406226
rect 597456 406046 597512 406102
rect 597580 406046 597636 406102
rect 597704 406046 597760 406102
rect 597828 406046 597884 406102
rect 597456 405922 597512 405978
rect 597580 405922 597636 405978
rect 597704 405922 597760 405978
rect 597828 405922 597884 405978
rect 597456 388294 597512 388350
rect 597580 388294 597636 388350
rect 597704 388294 597760 388350
rect 597828 388294 597884 388350
rect 597456 388170 597512 388226
rect 597580 388170 597636 388226
rect 597704 388170 597760 388226
rect 597828 388170 597884 388226
rect 597456 388046 597512 388102
rect 597580 388046 597636 388102
rect 597704 388046 597760 388102
rect 597828 388046 597884 388102
rect 597456 387922 597512 387978
rect 597580 387922 597636 387978
rect 597704 387922 597760 387978
rect 597828 387922 597884 387978
rect 597456 370294 597512 370350
rect 597580 370294 597636 370350
rect 597704 370294 597760 370350
rect 597828 370294 597884 370350
rect 597456 370170 597512 370226
rect 597580 370170 597636 370226
rect 597704 370170 597760 370226
rect 597828 370170 597884 370226
rect 597456 370046 597512 370102
rect 597580 370046 597636 370102
rect 597704 370046 597760 370102
rect 597828 370046 597884 370102
rect 597456 369922 597512 369978
rect 597580 369922 597636 369978
rect 597704 369922 597760 369978
rect 597828 369922 597884 369978
rect 597456 352294 597512 352350
rect 597580 352294 597636 352350
rect 597704 352294 597760 352350
rect 597828 352294 597884 352350
rect 597456 352170 597512 352226
rect 597580 352170 597636 352226
rect 597704 352170 597760 352226
rect 597828 352170 597884 352226
rect 597456 352046 597512 352102
rect 597580 352046 597636 352102
rect 597704 352046 597760 352102
rect 597828 352046 597884 352102
rect 597456 351922 597512 351978
rect 597580 351922 597636 351978
rect 597704 351922 597760 351978
rect 597828 351922 597884 351978
rect 597456 334294 597512 334350
rect 597580 334294 597636 334350
rect 597704 334294 597760 334350
rect 597828 334294 597884 334350
rect 597456 334170 597512 334226
rect 597580 334170 597636 334226
rect 597704 334170 597760 334226
rect 597828 334170 597884 334226
rect 597456 334046 597512 334102
rect 597580 334046 597636 334102
rect 597704 334046 597760 334102
rect 597828 334046 597884 334102
rect 597456 333922 597512 333978
rect 597580 333922 597636 333978
rect 597704 333922 597760 333978
rect 597828 333922 597884 333978
rect 597456 316294 597512 316350
rect 597580 316294 597636 316350
rect 597704 316294 597760 316350
rect 597828 316294 597884 316350
rect 597456 316170 597512 316226
rect 597580 316170 597636 316226
rect 597704 316170 597760 316226
rect 597828 316170 597884 316226
rect 597456 316046 597512 316102
rect 597580 316046 597636 316102
rect 597704 316046 597760 316102
rect 597828 316046 597884 316102
rect 597456 315922 597512 315978
rect 597580 315922 597636 315978
rect 597704 315922 597760 315978
rect 597828 315922 597884 315978
rect 597456 298294 597512 298350
rect 597580 298294 597636 298350
rect 597704 298294 597760 298350
rect 597828 298294 597884 298350
rect 597456 298170 597512 298226
rect 597580 298170 597636 298226
rect 597704 298170 597760 298226
rect 597828 298170 597884 298226
rect 597456 298046 597512 298102
rect 597580 298046 597636 298102
rect 597704 298046 597760 298102
rect 597828 298046 597884 298102
rect 597456 297922 597512 297978
rect 597580 297922 597636 297978
rect 597704 297922 597760 297978
rect 597828 297922 597884 297978
rect 597456 280294 597512 280350
rect 597580 280294 597636 280350
rect 597704 280294 597760 280350
rect 597828 280294 597884 280350
rect 597456 280170 597512 280226
rect 597580 280170 597636 280226
rect 597704 280170 597760 280226
rect 597828 280170 597884 280226
rect 597456 280046 597512 280102
rect 597580 280046 597636 280102
rect 597704 280046 597760 280102
rect 597828 280046 597884 280102
rect 597456 279922 597512 279978
rect 597580 279922 597636 279978
rect 597704 279922 597760 279978
rect 597828 279922 597884 279978
rect 597456 262294 597512 262350
rect 597580 262294 597636 262350
rect 597704 262294 597760 262350
rect 597828 262294 597884 262350
rect 597456 262170 597512 262226
rect 597580 262170 597636 262226
rect 597704 262170 597760 262226
rect 597828 262170 597884 262226
rect 597456 262046 597512 262102
rect 597580 262046 597636 262102
rect 597704 262046 597760 262102
rect 597828 262046 597884 262102
rect 597456 261922 597512 261978
rect 597580 261922 597636 261978
rect 597704 261922 597760 261978
rect 597828 261922 597884 261978
rect 597456 244294 597512 244350
rect 597580 244294 597636 244350
rect 597704 244294 597760 244350
rect 597828 244294 597884 244350
rect 597456 244170 597512 244226
rect 597580 244170 597636 244226
rect 597704 244170 597760 244226
rect 597828 244170 597884 244226
rect 597456 244046 597512 244102
rect 597580 244046 597636 244102
rect 597704 244046 597760 244102
rect 597828 244046 597884 244102
rect 597456 243922 597512 243978
rect 597580 243922 597636 243978
rect 597704 243922 597760 243978
rect 597828 243922 597884 243978
rect 597456 226294 597512 226350
rect 597580 226294 597636 226350
rect 597704 226294 597760 226350
rect 597828 226294 597884 226350
rect 597456 226170 597512 226226
rect 597580 226170 597636 226226
rect 597704 226170 597760 226226
rect 597828 226170 597884 226226
rect 597456 226046 597512 226102
rect 597580 226046 597636 226102
rect 597704 226046 597760 226102
rect 597828 226046 597884 226102
rect 597456 225922 597512 225978
rect 597580 225922 597636 225978
rect 597704 225922 597760 225978
rect 597828 225922 597884 225978
rect 597456 208294 597512 208350
rect 597580 208294 597636 208350
rect 597704 208294 597760 208350
rect 597828 208294 597884 208350
rect 597456 208170 597512 208226
rect 597580 208170 597636 208226
rect 597704 208170 597760 208226
rect 597828 208170 597884 208226
rect 597456 208046 597512 208102
rect 597580 208046 597636 208102
rect 597704 208046 597760 208102
rect 597828 208046 597884 208102
rect 597456 207922 597512 207978
rect 597580 207922 597636 207978
rect 597704 207922 597760 207978
rect 597828 207922 597884 207978
rect 597456 190294 597512 190350
rect 597580 190294 597636 190350
rect 597704 190294 597760 190350
rect 597828 190294 597884 190350
rect 597456 190170 597512 190226
rect 597580 190170 597636 190226
rect 597704 190170 597760 190226
rect 597828 190170 597884 190226
rect 597456 190046 597512 190102
rect 597580 190046 597636 190102
rect 597704 190046 597760 190102
rect 597828 190046 597884 190102
rect 597456 189922 597512 189978
rect 597580 189922 597636 189978
rect 597704 189922 597760 189978
rect 597828 189922 597884 189978
rect 597456 172294 597512 172350
rect 597580 172294 597636 172350
rect 597704 172294 597760 172350
rect 597828 172294 597884 172350
rect 597456 172170 597512 172226
rect 597580 172170 597636 172226
rect 597704 172170 597760 172226
rect 597828 172170 597884 172226
rect 597456 172046 597512 172102
rect 597580 172046 597636 172102
rect 597704 172046 597760 172102
rect 597828 172046 597884 172102
rect 597456 171922 597512 171978
rect 597580 171922 597636 171978
rect 597704 171922 597760 171978
rect 597828 171922 597884 171978
rect 597456 154294 597512 154350
rect 597580 154294 597636 154350
rect 597704 154294 597760 154350
rect 597828 154294 597884 154350
rect 597456 154170 597512 154226
rect 597580 154170 597636 154226
rect 597704 154170 597760 154226
rect 597828 154170 597884 154226
rect 597456 154046 597512 154102
rect 597580 154046 597636 154102
rect 597704 154046 597760 154102
rect 597828 154046 597884 154102
rect 597456 153922 597512 153978
rect 597580 153922 597636 153978
rect 597704 153922 597760 153978
rect 597828 153922 597884 153978
rect 597456 136294 597512 136350
rect 597580 136294 597636 136350
rect 597704 136294 597760 136350
rect 597828 136294 597884 136350
rect 597456 136170 597512 136226
rect 597580 136170 597636 136226
rect 597704 136170 597760 136226
rect 597828 136170 597884 136226
rect 597456 136046 597512 136102
rect 597580 136046 597636 136102
rect 597704 136046 597760 136102
rect 597828 136046 597884 136102
rect 597456 135922 597512 135978
rect 597580 135922 597636 135978
rect 597704 135922 597760 135978
rect 597828 135922 597884 135978
rect 597456 118294 597512 118350
rect 597580 118294 597636 118350
rect 597704 118294 597760 118350
rect 597828 118294 597884 118350
rect 597456 118170 597512 118226
rect 597580 118170 597636 118226
rect 597704 118170 597760 118226
rect 597828 118170 597884 118226
rect 597456 118046 597512 118102
rect 597580 118046 597636 118102
rect 597704 118046 597760 118102
rect 597828 118046 597884 118102
rect 597456 117922 597512 117978
rect 597580 117922 597636 117978
rect 597704 117922 597760 117978
rect 597828 117922 597884 117978
rect 597456 100294 597512 100350
rect 597580 100294 597636 100350
rect 597704 100294 597760 100350
rect 597828 100294 597884 100350
rect 597456 100170 597512 100226
rect 597580 100170 597636 100226
rect 597704 100170 597760 100226
rect 597828 100170 597884 100226
rect 597456 100046 597512 100102
rect 597580 100046 597636 100102
rect 597704 100046 597760 100102
rect 597828 100046 597884 100102
rect 597456 99922 597512 99978
rect 597580 99922 597636 99978
rect 597704 99922 597760 99978
rect 597828 99922 597884 99978
rect 597456 82294 597512 82350
rect 597580 82294 597636 82350
rect 597704 82294 597760 82350
rect 597828 82294 597884 82350
rect 597456 82170 597512 82226
rect 597580 82170 597636 82226
rect 597704 82170 597760 82226
rect 597828 82170 597884 82226
rect 597456 82046 597512 82102
rect 597580 82046 597636 82102
rect 597704 82046 597760 82102
rect 597828 82046 597884 82102
rect 597456 81922 597512 81978
rect 597580 81922 597636 81978
rect 597704 81922 597760 81978
rect 597828 81922 597884 81978
rect 597456 64294 597512 64350
rect 597580 64294 597636 64350
rect 597704 64294 597760 64350
rect 597828 64294 597884 64350
rect 597456 64170 597512 64226
rect 597580 64170 597636 64226
rect 597704 64170 597760 64226
rect 597828 64170 597884 64226
rect 597456 64046 597512 64102
rect 597580 64046 597636 64102
rect 597704 64046 597760 64102
rect 597828 64046 597884 64102
rect 597456 63922 597512 63978
rect 597580 63922 597636 63978
rect 597704 63922 597760 63978
rect 597828 63922 597884 63978
rect 597456 46294 597512 46350
rect 597580 46294 597636 46350
rect 597704 46294 597760 46350
rect 597828 46294 597884 46350
rect 597456 46170 597512 46226
rect 597580 46170 597636 46226
rect 597704 46170 597760 46226
rect 597828 46170 597884 46226
rect 597456 46046 597512 46102
rect 597580 46046 597636 46102
rect 597704 46046 597760 46102
rect 597828 46046 597884 46102
rect 597456 45922 597512 45978
rect 597580 45922 597636 45978
rect 597704 45922 597760 45978
rect 597828 45922 597884 45978
rect 597456 28294 597512 28350
rect 597580 28294 597636 28350
rect 597704 28294 597760 28350
rect 597828 28294 597884 28350
rect 597456 28170 597512 28226
rect 597580 28170 597636 28226
rect 597704 28170 597760 28226
rect 597828 28170 597884 28226
rect 597456 28046 597512 28102
rect 597580 28046 597636 28102
rect 597704 28046 597760 28102
rect 597828 28046 597884 28102
rect 597456 27922 597512 27978
rect 597580 27922 597636 27978
rect 597704 27922 597760 27978
rect 597828 27922 597884 27978
rect 597456 10294 597512 10350
rect 597580 10294 597636 10350
rect 597704 10294 597760 10350
rect 597828 10294 597884 10350
rect 597456 10170 597512 10226
rect 597580 10170 597636 10226
rect 597704 10170 597760 10226
rect 597828 10170 597884 10226
rect 597456 10046 597512 10102
rect 597580 10046 597636 10102
rect 597704 10046 597760 10102
rect 597828 10046 597884 10102
rect 597456 9922 597512 9978
rect 597580 9922 597636 9978
rect 597704 9922 597760 9978
rect 597828 9922 597884 9978
rect 582970 -1176 583026 -1120
rect 583094 -1176 583150 -1120
rect 583218 -1176 583274 -1120
rect 583342 -1176 583398 -1120
rect 582970 -1300 583026 -1244
rect 583094 -1300 583150 -1244
rect 583218 -1300 583274 -1244
rect 583342 -1300 583398 -1244
rect 582970 -1424 583026 -1368
rect 583094 -1424 583150 -1368
rect 583218 -1424 583274 -1368
rect 583342 -1424 583398 -1368
rect 582970 -1548 583026 -1492
rect 583094 -1548 583150 -1492
rect 583218 -1548 583274 -1492
rect 583342 -1548 583398 -1492
rect 597456 -1176 597512 -1120
rect 597580 -1176 597636 -1120
rect 597704 -1176 597760 -1120
rect 597828 -1176 597884 -1120
rect 597456 -1300 597512 -1244
rect 597580 -1300 597636 -1244
rect 597704 -1300 597760 -1244
rect 597828 -1300 597884 -1244
rect 597456 -1424 597512 -1368
rect 597580 -1424 597636 -1368
rect 597704 -1424 597760 -1368
rect 597828 -1424 597884 -1368
rect 597456 -1548 597512 -1492
rect 597580 -1548 597636 -1492
rect 597704 -1548 597760 -1492
rect 597828 -1548 597884 -1492
<< metal5 >>
rect -1916 598172 597980 598268
rect -1916 598116 -1820 598172
rect -1764 598116 -1696 598172
rect -1640 598116 -1572 598172
rect -1516 598116 -1448 598172
rect -1392 598116 6970 598172
rect 7026 598116 7094 598172
rect 7150 598116 7218 598172
rect 7274 598116 7342 598172
rect 7398 598116 24970 598172
rect 25026 598116 25094 598172
rect 25150 598116 25218 598172
rect 25274 598116 25342 598172
rect 25398 598116 42970 598172
rect 43026 598116 43094 598172
rect 43150 598116 43218 598172
rect 43274 598116 43342 598172
rect 43398 598116 60970 598172
rect 61026 598116 61094 598172
rect 61150 598116 61218 598172
rect 61274 598116 61342 598172
rect 61398 598116 78970 598172
rect 79026 598116 79094 598172
rect 79150 598116 79218 598172
rect 79274 598116 79342 598172
rect 79398 598116 96970 598172
rect 97026 598116 97094 598172
rect 97150 598116 97218 598172
rect 97274 598116 97342 598172
rect 97398 598116 114970 598172
rect 115026 598116 115094 598172
rect 115150 598116 115218 598172
rect 115274 598116 115342 598172
rect 115398 598116 132970 598172
rect 133026 598116 133094 598172
rect 133150 598116 133218 598172
rect 133274 598116 133342 598172
rect 133398 598116 150970 598172
rect 151026 598116 151094 598172
rect 151150 598116 151218 598172
rect 151274 598116 151342 598172
rect 151398 598116 168970 598172
rect 169026 598116 169094 598172
rect 169150 598116 169218 598172
rect 169274 598116 169342 598172
rect 169398 598116 186970 598172
rect 187026 598116 187094 598172
rect 187150 598116 187218 598172
rect 187274 598116 187342 598172
rect 187398 598116 204970 598172
rect 205026 598116 205094 598172
rect 205150 598116 205218 598172
rect 205274 598116 205342 598172
rect 205398 598116 222970 598172
rect 223026 598116 223094 598172
rect 223150 598116 223218 598172
rect 223274 598116 223342 598172
rect 223398 598116 240970 598172
rect 241026 598116 241094 598172
rect 241150 598116 241218 598172
rect 241274 598116 241342 598172
rect 241398 598116 258970 598172
rect 259026 598116 259094 598172
rect 259150 598116 259218 598172
rect 259274 598116 259342 598172
rect 259398 598116 276970 598172
rect 277026 598116 277094 598172
rect 277150 598116 277218 598172
rect 277274 598116 277342 598172
rect 277398 598116 294970 598172
rect 295026 598116 295094 598172
rect 295150 598116 295218 598172
rect 295274 598116 295342 598172
rect 295398 598116 312970 598172
rect 313026 598116 313094 598172
rect 313150 598116 313218 598172
rect 313274 598116 313342 598172
rect 313398 598116 330970 598172
rect 331026 598116 331094 598172
rect 331150 598116 331218 598172
rect 331274 598116 331342 598172
rect 331398 598116 348970 598172
rect 349026 598116 349094 598172
rect 349150 598116 349218 598172
rect 349274 598116 349342 598172
rect 349398 598116 366970 598172
rect 367026 598116 367094 598172
rect 367150 598116 367218 598172
rect 367274 598116 367342 598172
rect 367398 598116 384970 598172
rect 385026 598116 385094 598172
rect 385150 598116 385218 598172
rect 385274 598116 385342 598172
rect 385398 598116 402970 598172
rect 403026 598116 403094 598172
rect 403150 598116 403218 598172
rect 403274 598116 403342 598172
rect 403398 598116 420970 598172
rect 421026 598116 421094 598172
rect 421150 598116 421218 598172
rect 421274 598116 421342 598172
rect 421398 598116 438970 598172
rect 439026 598116 439094 598172
rect 439150 598116 439218 598172
rect 439274 598116 439342 598172
rect 439398 598116 456970 598172
rect 457026 598116 457094 598172
rect 457150 598116 457218 598172
rect 457274 598116 457342 598172
rect 457398 598116 474970 598172
rect 475026 598116 475094 598172
rect 475150 598116 475218 598172
rect 475274 598116 475342 598172
rect 475398 598116 492970 598172
rect 493026 598116 493094 598172
rect 493150 598116 493218 598172
rect 493274 598116 493342 598172
rect 493398 598116 510970 598172
rect 511026 598116 511094 598172
rect 511150 598116 511218 598172
rect 511274 598116 511342 598172
rect 511398 598116 528970 598172
rect 529026 598116 529094 598172
rect 529150 598116 529218 598172
rect 529274 598116 529342 598172
rect 529398 598116 546970 598172
rect 547026 598116 547094 598172
rect 547150 598116 547218 598172
rect 547274 598116 547342 598172
rect 547398 598116 564970 598172
rect 565026 598116 565094 598172
rect 565150 598116 565218 598172
rect 565274 598116 565342 598172
rect 565398 598116 582970 598172
rect 583026 598116 583094 598172
rect 583150 598116 583218 598172
rect 583274 598116 583342 598172
rect 583398 598116 597456 598172
rect 597512 598116 597580 598172
rect 597636 598116 597704 598172
rect 597760 598116 597828 598172
rect 597884 598116 597980 598172
rect -1916 598048 597980 598116
rect -1916 597992 -1820 598048
rect -1764 597992 -1696 598048
rect -1640 597992 -1572 598048
rect -1516 597992 -1448 598048
rect -1392 597992 6970 598048
rect 7026 597992 7094 598048
rect 7150 597992 7218 598048
rect 7274 597992 7342 598048
rect 7398 597992 24970 598048
rect 25026 597992 25094 598048
rect 25150 597992 25218 598048
rect 25274 597992 25342 598048
rect 25398 597992 42970 598048
rect 43026 597992 43094 598048
rect 43150 597992 43218 598048
rect 43274 597992 43342 598048
rect 43398 597992 60970 598048
rect 61026 597992 61094 598048
rect 61150 597992 61218 598048
rect 61274 597992 61342 598048
rect 61398 597992 78970 598048
rect 79026 597992 79094 598048
rect 79150 597992 79218 598048
rect 79274 597992 79342 598048
rect 79398 597992 96970 598048
rect 97026 597992 97094 598048
rect 97150 597992 97218 598048
rect 97274 597992 97342 598048
rect 97398 597992 114970 598048
rect 115026 597992 115094 598048
rect 115150 597992 115218 598048
rect 115274 597992 115342 598048
rect 115398 597992 132970 598048
rect 133026 597992 133094 598048
rect 133150 597992 133218 598048
rect 133274 597992 133342 598048
rect 133398 597992 150970 598048
rect 151026 597992 151094 598048
rect 151150 597992 151218 598048
rect 151274 597992 151342 598048
rect 151398 597992 168970 598048
rect 169026 597992 169094 598048
rect 169150 597992 169218 598048
rect 169274 597992 169342 598048
rect 169398 597992 186970 598048
rect 187026 597992 187094 598048
rect 187150 597992 187218 598048
rect 187274 597992 187342 598048
rect 187398 597992 204970 598048
rect 205026 597992 205094 598048
rect 205150 597992 205218 598048
rect 205274 597992 205342 598048
rect 205398 597992 222970 598048
rect 223026 597992 223094 598048
rect 223150 597992 223218 598048
rect 223274 597992 223342 598048
rect 223398 597992 240970 598048
rect 241026 597992 241094 598048
rect 241150 597992 241218 598048
rect 241274 597992 241342 598048
rect 241398 597992 258970 598048
rect 259026 597992 259094 598048
rect 259150 597992 259218 598048
rect 259274 597992 259342 598048
rect 259398 597992 276970 598048
rect 277026 597992 277094 598048
rect 277150 597992 277218 598048
rect 277274 597992 277342 598048
rect 277398 597992 294970 598048
rect 295026 597992 295094 598048
rect 295150 597992 295218 598048
rect 295274 597992 295342 598048
rect 295398 597992 312970 598048
rect 313026 597992 313094 598048
rect 313150 597992 313218 598048
rect 313274 597992 313342 598048
rect 313398 597992 330970 598048
rect 331026 597992 331094 598048
rect 331150 597992 331218 598048
rect 331274 597992 331342 598048
rect 331398 597992 348970 598048
rect 349026 597992 349094 598048
rect 349150 597992 349218 598048
rect 349274 597992 349342 598048
rect 349398 597992 366970 598048
rect 367026 597992 367094 598048
rect 367150 597992 367218 598048
rect 367274 597992 367342 598048
rect 367398 597992 384970 598048
rect 385026 597992 385094 598048
rect 385150 597992 385218 598048
rect 385274 597992 385342 598048
rect 385398 597992 402970 598048
rect 403026 597992 403094 598048
rect 403150 597992 403218 598048
rect 403274 597992 403342 598048
rect 403398 597992 420970 598048
rect 421026 597992 421094 598048
rect 421150 597992 421218 598048
rect 421274 597992 421342 598048
rect 421398 597992 438970 598048
rect 439026 597992 439094 598048
rect 439150 597992 439218 598048
rect 439274 597992 439342 598048
rect 439398 597992 456970 598048
rect 457026 597992 457094 598048
rect 457150 597992 457218 598048
rect 457274 597992 457342 598048
rect 457398 597992 474970 598048
rect 475026 597992 475094 598048
rect 475150 597992 475218 598048
rect 475274 597992 475342 598048
rect 475398 597992 492970 598048
rect 493026 597992 493094 598048
rect 493150 597992 493218 598048
rect 493274 597992 493342 598048
rect 493398 597992 510970 598048
rect 511026 597992 511094 598048
rect 511150 597992 511218 598048
rect 511274 597992 511342 598048
rect 511398 597992 528970 598048
rect 529026 597992 529094 598048
rect 529150 597992 529218 598048
rect 529274 597992 529342 598048
rect 529398 597992 546970 598048
rect 547026 597992 547094 598048
rect 547150 597992 547218 598048
rect 547274 597992 547342 598048
rect 547398 597992 564970 598048
rect 565026 597992 565094 598048
rect 565150 597992 565218 598048
rect 565274 597992 565342 598048
rect 565398 597992 582970 598048
rect 583026 597992 583094 598048
rect 583150 597992 583218 598048
rect 583274 597992 583342 598048
rect 583398 597992 597456 598048
rect 597512 597992 597580 598048
rect 597636 597992 597704 598048
rect 597760 597992 597828 598048
rect 597884 597992 597980 598048
rect -1916 597924 597980 597992
rect -1916 597868 -1820 597924
rect -1764 597868 -1696 597924
rect -1640 597868 -1572 597924
rect -1516 597868 -1448 597924
rect -1392 597868 6970 597924
rect 7026 597868 7094 597924
rect 7150 597868 7218 597924
rect 7274 597868 7342 597924
rect 7398 597868 24970 597924
rect 25026 597868 25094 597924
rect 25150 597868 25218 597924
rect 25274 597868 25342 597924
rect 25398 597868 42970 597924
rect 43026 597868 43094 597924
rect 43150 597868 43218 597924
rect 43274 597868 43342 597924
rect 43398 597868 60970 597924
rect 61026 597868 61094 597924
rect 61150 597868 61218 597924
rect 61274 597868 61342 597924
rect 61398 597868 78970 597924
rect 79026 597868 79094 597924
rect 79150 597868 79218 597924
rect 79274 597868 79342 597924
rect 79398 597868 96970 597924
rect 97026 597868 97094 597924
rect 97150 597868 97218 597924
rect 97274 597868 97342 597924
rect 97398 597868 114970 597924
rect 115026 597868 115094 597924
rect 115150 597868 115218 597924
rect 115274 597868 115342 597924
rect 115398 597868 132970 597924
rect 133026 597868 133094 597924
rect 133150 597868 133218 597924
rect 133274 597868 133342 597924
rect 133398 597868 150970 597924
rect 151026 597868 151094 597924
rect 151150 597868 151218 597924
rect 151274 597868 151342 597924
rect 151398 597868 168970 597924
rect 169026 597868 169094 597924
rect 169150 597868 169218 597924
rect 169274 597868 169342 597924
rect 169398 597868 186970 597924
rect 187026 597868 187094 597924
rect 187150 597868 187218 597924
rect 187274 597868 187342 597924
rect 187398 597868 204970 597924
rect 205026 597868 205094 597924
rect 205150 597868 205218 597924
rect 205274 597868 205342 597924
rect 205398 597868 222970 597924
rect 223026 597868 223094 597924
rect 223150 597868 223218 597924
rect 223274 597868 223342 597924
rect 223398 597868 240970 597924
rect 241026 597868 241094 597924
rect 241150 597868 241218 597924
rect 241274 597868 241342 597924
rect 241398 597868 258970 597924
rect 259026 597868 259094 597924
rect 259150 597868 259218 597924
rect 259274 597868 259342 597924
rect 259398 597868 276970 597924
rect 277026 597868 277094 597924
rect 277150 597868 277218 597924
rect 277274 597868 277342 597924
rect 277398 597868 294970 597924
rect 295026 597868 295094 597924
rect 295150 597868 295218 597924
rect 295274 597868 295342 597924
rect 295398 597868 312970 597924
rect 313026 597868 313094 597924
rect 313150 597868 313218 597924
rect 313274 597868 313342 597924
rect 313398 597868 330970 597924
rect 331026 597868 331094 597924
rect 331150 597868 331218 597924
rect 331274 597868 331342 597924
rect 331398 597868 348970 597924
rect 349026 597868 349094 597924
rect 349150 597868 349218 597924
rect 349274 597868 349342 597924
rect 349398 597868 366970 597924
rect 367026 597868 367094 597924
rect 367150 597868 367218 597924
rect 367274 597868 367342 597924
rect 367398 597868 384970 597924
rect 385026 597868 385094 597924
rect 385150 597868 385218 597924
rect 385274 597868 385342 597924
rect 385398 597868 402970 597924
rect 403026 597868 403094 597924
rect 403150 597868 403218 597924
rect 403274 597868 403342 597924
rect 403398 597868 420970 597924
rect 421026 597868 421094 597924
rect 421150 597868 421218 597924
rect 421274 597868 421342 597924
rect 421398 597868 438970 597924
rect 439026 597868 439094 597924
rect 439150 597868 439218 597924
rect 439274 597868 439342 597924
rect 439398 597868 456970 597924
rect 457026 597868 457094 597924
rect 457150 597868 457218 597924
rect 457274 597868 457342 597924
rect 457398 597868 474970 597924
rect 475026 597868 475094 597924
rect 475150 597868 475218 597924
rect 475274 597868 475342 597924
rect 475398 597868 492970 597924
rect 493026 597868 493094 597924
rect 493150 597868 493218 597924
rect 493274 597868 493342 597924
rect 493398 597868 510970 597924
rect 511026 597868 511094 597924
rect 511150 597868 511218 597924
rect 511274 597868 511342 597924
rect 511398 597868 528970 597924
rect 529026 597868 529094 597924
rect 529150 597868 529218 597924
rect 529274 597868 529342 597924
rect 529398 597868 546970 597924
rect 547026 597868 547094 597924
rect 547150 597868 547218 597924
rect 547274 597868 547342 597924
rect 547398 597868 564970 597924
rect 565026 597868 565094 597924
rect 565150 597868 565218 597924
rect 565274 597868 565342 597924
rect 565398 597868 582970 597924
rect 583026 597868 583094 597924
rect 583150 597868 583218 597924
rect 583274 597868 583342 597924
rect 583398 597868 597456 597924
rect 597512 597868 597580 597924
rect 597636 597868 597704 597924
rect 597760 597868 597828 597924
rect 597884 597868 597980 597924
rect -1916 597800 597980 597868
rect -1916 597744 -1820 597800
rect -1764 597744 -1696 597800
rect -1640 597744 -1572 597800
rect -1516 597744 -1448 597800
rect -1392 597744 6970 597800
rect 7026 597744 7094 597800
rect 7150 597744 7218 597800
rect 7274 597744 7342 597800
rect 7398 597744 24970 597800
rect 25026 597744 25094 597800
rect 25150 597744 25218 597800
rect 25274 597744 25342 597800
rect 25398 597744 42970 597800
rect 43026 597744 43094 597800
rect 43150 597744 43218 597800
rect 43274 597744 43342 597800
rect 43398 597744 60970 597800
rect 61026 597744 61094 597800
rect 61150 597744 61218 597800
rect 61274 597744 61342 597800
rect 61398 597744 78970 597800
rect 79026 597744 79094 597800
rect 79150 597744 79218 597800
rect 79274 597744 79342 597800
rect 79398 597744 96970 597800
rect 97026 597744 97094 597800
rect 97150 597744 97218 597800
rect 97274 597744 97342 597800
rect 97398 597744 114970 597800
rect 115026 597744 115094 597800
rect 115150 597744 115218 597800
rect 115274 597744 115342 597800
rect 115398 597744 132970 597800
rect 133026 597744 133094 597800
rect 133150 597744 133218 597800
rect 133274 597744 133342 597800
rect 133398 597744 150970 597800
rect 151026 597744 151094 597800
rect 151150 597744 151218 597800
rect 151274 597744 151342 597800
rect 151398 597744 168970 597800
rect 169026 597744 169094 597800
rect 169150 597744 169218 597800
rect 169274 597744 169342 597800
rect 169398 597744 186970 597800
rect 187026 597744 187094 597800
rect 187150 597744 187218 597800
rect 187274 597744 187342 597800
rect 187398 597744 204970 597800
rect 205026 597744 205094 597800
rect 205150 597744 205218 597800
rect 205274 597744 205342 597800
rect 205398 597744 222970 597800
rect 223026 597744 223094 597800
rect 223150 597744 223218 597800
rect 223274 597744 223342 597800
rect 223398 597744 240970 597800
rect 241026 597744 241094 597800
rect 241150 597744 241218 597800
rect 241274 597744 241342 597800
rect 241398 597744 258970 597800
rect 259026 597744 259094 597800
rect 259150 597744 259218 597800
rect 259274 597744 259342 597800
rect 259398 597744 276970 597800
rect 277026 597744 277094 597800
rect 277150 597744 277218 597800
rect 277274 597744 277342 597800
rect 277398 597744 294970 597800
rect 295026 597744 295094 597800
rect 295150 597744 295218 597800
rect 295274 597744 295342 597800
rect 295398 597744 312970 597800
rect 313026 597744 313094 597800
rect 313150 597744 313218 597800
rect 313274 597744 313342 597800
rect 313398 597744 330970 597800
rect 331026 597744 331094 597800
rect 331150 597744 331218 597800
rect 331274 597744 331342 597800
rect 331398 597744 348970 597800
rect 349026 597744 349094 597800
rect 349150 597744 349218 597800
rect 349274 597744 349342 597800
rect 349398 597744 366970 597800
rect 367026 597744 367094 597800
rect 367150 597744 367218 597800
rect 367274 597744 367342 597800
rect 367398 597744 384970 597800
rect 385026 597744 385094 597800
rect 385150 597744 385218 597800
rect 385274 597744 385342 597800
rect 385398 597744 402970 597800
rect 403026 597744 403094 597800
rect 403150 597744 403218 597800
rect 403274 597744 403342 597800
rect 403398 597744 420970 597800
rect 421026 597744 421094 597800
rect 421150 597744 421218 597800
rect 421274 597744 421342 597800
rect 421398 597744 438970 597800
rect 439026 597744 439094 597800
rect 439150 597744 439218 597800
rect 439274 597744 439342 597800
rect 439398 597744 456970 597800
rect 457026 597744 457094 597800
rect 457150 597744 457218 597800
rect 457274 597744 457342 597800
rect 457398 597744 474970 597800
rect 475026 597744 475094 597800
rect 475150 597744 475218 597800
rect 475274 597744 475342 597800
rect 475398 597744 492970 597800
rect 493026 597744 493094 597800
rect 493150 597744 493218 597800
rect 493274 597744 493342 597800
rect 493398 597744 510970 597800
rect 511026 597744 511094 597800
rect 511150 597744 511218 597800
rect 511274 597744 511342 597800
rect 511398 597744 528970 597800
rect 529026 597744 529094 597800
rect 529150 597744 529218 597800
rect 529274 597744 529342 597800
rect 529398 597744 546970 597800
rect 547026 597744 547094 597800
rect 547150 597744 547218 597800
rect 547274 597744 547342 597800
rect 547398 597744 564970 597800
rect 565026 597744 565094 597800
rect 565150 597744 565218 597800
rect 565274 597744 565342 597800
rect 565398 597744 582970 597800
rect 583026 597744 583094 597800
rect 583150 597744 583218 597800
rect 583274 597744 583342 597800
rect 583398 597744 597456 597800
rect 597512 597744 597580 597800
rect 597636 597744 597704 597800
rect 597760 597744 597828 597800
rect 597884 597744 597980 597800
rect -1916 597648 597980 597744
rect -956 597212 597020 597308
rect -956 597156 -860 597212
rect -804 597156 -736 597212
rect -680 597156 -612 597212
rect -556 597156 -488 597212
rect -432 597156 3250 597212
rect 3306 597156 3374 597212
rect 3430 597156 3498 597212
rect 3554 597156 3622 597212
rect 3678 597156 21250 597212
rect 21306 597156 21374 597212
rect 21430 597156 21498 597212
rect 21554 597156 21622 597212
rect 21678 597156 39250 597212
rect 39306 597156 39374 597212
rect 39430 597156 39498 597212
rect 39554 597156 39622 597212
rect 39678 597156 57250 597212
rect 57306 597156 57374 597212
rect 57430 597156 57498 597212
rect 57554 597156 57622 597212
rect 57678 597156 75250 597212
rect 75306 597156 75374 597212
rect 75430 597156 75498 597212
rect 75554 597156 75622 597212
rect 75678 597156 93250 597212
rect 93306 597156 93374 597212
rect 93430 597156 93498 597212
rect 93554 597156 93622 597212
rect 93678 597156 111250 597212
rect 111306 597156 111374 597212
rect 111430 597156 111498 597212
rect 111554 597156 111622 597212
rect 111678 597156 129250 597212
rect 129306 597156 129374 597212
rect 129430 597156 129498 597212
rect 129554 597156 129622 597212
rect 129678 597156 147250 597212
rect 147306 597156 147374 597212
rect 147430 597156 147498 597212
rect 147554 597156 147622 597212
rect 147678 597156 165250 597212
rect 165306 597156 165374 597212
rect 165430 597156 165498 597212
rect 165554 597156 165622 597212
rect 165678 597156 183250 597212
rect 183306 597156 183374 597212
rect 183430 597156 183498 597212
rect 183554 597156 183622 597212
rect 183678 597156 201250 597212
rect 201306 597156 201374 597212
rect 201430 597156 201498 597212
rect 201554 597156 201622 597212
rect 201678 597156 219250 597212
rect 219306 597156 219374 597212
rect 219430 597156 219498 597212
rect 219554 597156 219622 597212
rect 219678 597156 237250 597212
rect 237306 597156 237374 597212
rect 237430 597156 237498 597212
rect 237554 597156 237622 597212
rect 237678 597156 255250 597212
rect 255306 597156 255374 597212
rect 255430 597156 255498 597212
rect 255554 597156 255622 597212
rect 255678 597156 273250 597212
rect 273306 597156 273374 597212
rect 273430 597156 273498 597212
rect 273554 597156 273622 597212
rect 273678 597156 291250 597212
rect 291306 597156 291374 597212
rect 291430 597156 291498 597212
rect 291554 597156 291622 597212
rect 291678 597156 309250 597212
rect 309306 597156 309374 597212
rect 309430 597156 309498 597212
rect 309554 597156 309622 597212
rect 309678 597156 327250 597212
rect 327306 597156 327374 597212
rect 327430 597156 327498 597212
rect 327554 597156 327622 597212
rect 327678 597156 345250 597212
rect 345306 597156 345374 597212
rect 345430 597156 345498 597212
rect 345554 597156 345622 597212
rect 345678 597156 363250 597212
rect 363306 597156 363374 597212
rect 363430 597156 363498 597212
rect 363554 597156 363622 597212
rect 363678 597156 381250 597212
rect 381306 597156 381374 597212
rect 381430 597156 381498 597212
rect 381554 597156 381622 597212
rect 381678 597156 399250 597212
rect 399306 597156 399374 597212
rect 399430 597156 399498 597212
rect 399554 597156 399622 597212
rect 399678 597156 417250 597212
rect 417306 597156 417374 597212
rect 417430 597156 417498 597212
rect 417554 597156 417622 597212
rect 417678 597156 435250 597212
rect 435306 597156 435374 597212
rect 435430 597156 435498 597212
rect 435554 597156 435622 597212
rect 435678 597156 453250 597212
rect 453306 597156 453374 597212
rect 453430 597156 453498 597212
rect 453554 597156 453622 597212
rect 453678 597156 471250 597212
rect 471306 597156 471374 597212
rect 471430 597156 471498 597212
rect 471554 597156 471622 597212
rect 471678 597156 489250 597212
rect 489306 597156 489374 597212
rect 489430 597156 489498 597212
rect 489554 597156 489622 597212
rect 489678 597156 507250 597212
rect 507306 597156 507374 597212
rect 507430 597156 507498 597212
rect 507554 597156 507622 597212
rect 507678 597156 525250 597212
rect 525306 597156 525374 597212
rect 525430 597156 525498 597212
rect 525554 597156 525622 597212
rect 525678 597156 543250 597212
rect 543306 597156 543374 597212
rect 543430 597156 543498 597212
rect 543554 597156 543622 597212
rect 543678 597156 561250 597212
rect 561306 597156 561374 597212
rect 561430 597156 561498 597212
rect 561554 597156 561622 597212
rect 561678 597156 579250 597212
rect 579306 597156 579374 597212
rect 579430 597156 579498 597212
rect 579554 597156 579622 597212
rect 579678 597156 596496 597212
rect 596552 597156 596620 597212
rect 596676 597156 596744 597212
rect 596800 597156 596868 597212
rect 596924 597156 597020 597212
rect -956 597088 597020 597156
rect -956 597032 -860 597088
rect -804 597032 -736 597088
rect -680 597032 -612 597088
rect -556 597032 -488 597088
rect -432 597032 3250 597088
rect 3306 597032 3374 597088
rect 3430 597032 3498 597088
rect 3554 597032 3622 597088
rect 3678 597032 21250 597088
rect 21306 597032 21374 597088
rect 21430 597032 21498 597088
rect 21554 597032 21622 597088
rect 21678 597032 39250 597088
rect 39306 597032 39374 597088
rect 39430 597032 39498 597088
rect 39554 597032 39622 597088
rect 39678 597032 57250 597088
rect 57306 597032 57374 597088
rect 57430 597032 57498 597088
rect 57554 597032 57622 597088
rect 57678 597032 75250 597088
rect 75306 597032 75374 597088
rect 75430 597032 75498 597088
rect 75554 597032 75622 597088
rect 75678 597032 93250 597088
rect 93306 597032 93374 597088
rect 93430 597032 93498 597088
rect 93554 597032 93622 597088
rect 93678 597032 111250 597088
rect 111306 597032 111374 597088
rect 111430 597032 111498 597088
rect 111554 597032 111622 597088
rect 111678 597032 129250 597088
rect 129306 597032 129374 597088
rect 129430 597032 129498 597088
rect 129554 597032 129622 597088
rect 129678 597032 147250 597088
rect 147306 597032 147374 597088
rect 147430 597032 147498 597088
rect 147554 597032 147622 597088
rect 147678 597032 165250 597088
rect 165306 597032 165374 597088
rect 165430 597032 165498 597088
rect 165554 597032 165622 597088
rect 165678 597032 183250 597088
rect 183306 597032 183374 597088
rect 183430 597032 183498 597088
rect 183554 597032 183622 597088
rect 183678 597032 201250 597088
rect 201306 597032 201374 597088
rect 201430 597032 201498 597088
rect 201554 597032 201622 597088
rect 201678 597032 219250 597088
rect 219306 597032 219374 597088
rect 219430 597032 219498 597088
rect 219554 597032 219622 597088
rect 219678 597032 237250 597088
rect 237306 597032 237374 597088
rect 237430 597032 237498 597088
rect 237554 597032 237622 597088
rect 237678 597032 255250 597088
rect 255306 597032 255374 597088
rect 255430 597032 255498 597088
rect 255554 597032 255622 597088
rect 255678 597032 273250 597088
rect 273306 597032 273374 597088
rect 273430 597032 273498 597088
rect 273554 597032 273622 597088
rect 273678 597032 291250 597088
rect 291306 597032 291374 597088
rect 291430 597032 291498 597088
rect 291554 597032 291622 597088
rect 291678 597032 309250 597088
rect 309306 597032 309374 597088
rect 309430 597032 309498 597088
rect 309554 597032 309622 597088
rect 309678 597032 327250 597088
rect 327306 597032 327374 597088
rect 327430 597032 327498 597088
rect 327554 597032 327622 597088
rect 327678 597032 345250 597088
rect 345306 597032 345374 597088
rect 345430 597032 345498 597088
rect 345554 597032 345622 597088
rect 345678 597032 363250 597088
rect 363306 597032 363374 597088
rect 363430 597032 363498 597088
rect 363554 597032 363622 597088
rect 363678 597032 381250 597088
rect 381306 597032 381374 597088
rect 381430 597032 381498 597088
rect 381554 597032 381622 597088
rect 381678 597032 399250 597088
rect 399306 597032 399374 597088
rect 399430 597032 399498 597088
rect 399554 597032 399622 597088
rect 399678 597032 417250 597088
rect 417306 597032 417374 597088
rect 417430 597032 417498 597088
rect 417554 597032 417622 597088
rect 417678 597032 435250 597088
rect 435306 597032 435374 597088
rect 435430 597032 435498 597088
rect 435554 597032 435622 597088
rect 435678 597032 453250 597088
rect 453306 597032 453374 597088
rect 453430 597032 453498 597088
rect 453554 597032 453622 597088
rect 453678 597032 471250 597088
rect 471306 597032 471374 597088
rect 471430 597032 471498 597088
rect 471554 597032 471622 597088
rect 471678 597032 489250 597088
rect 489306 597032 489374 597088
rect 489430 597032 489498 597088
rect 489554 597032 489622 597088
rect 489678 597032 507250 597088
rect 507306 597032 507374 597088
rect 507430 597032 507498 597088
rect 507554 597032 507622 597088
rect 507678 597032 525250 597088
rect 525306 597032 525374 597088
rect 525430 597032 525498 597088
rect 525554 597032 525622 597088
rect 525678 597032 543250 597088
rect 543306 597032 543374 597088
rect 543430 597032 543498 597088
rect 543554 597032 543622 597088
rect 543678 597032 561250 597088
rect 561306 597032 561374 597088
rect 561430 597032 561498 597088
rect 561554 597032 561622 597088
rect 561678 597032 579250 597088
rect 579306 597032 579374 597088
rect 579430 597032 579498 597088
rect 579554 597032 579622 597088
rect 579678 597032 596496 597088
rect 596552 597032 596620 597088
rect 596676 597032 596744 597088
rect 596800 597032 596868 597088
rect 596924 597032 597020 597088
rect -956 596964 597020 597032
rect -956 596908 -860 596964
rect -804 596908 -736 596964
rect -680 596908 -612 596964
rect -556 596908 -488 596964
rect -432 596908 3250 596964
rect 3306 596908 3374 596964
rect 3430 596908 3498 596964
rect 3554 596908 3622 596964
rect 3678 596908 21250 596964
rect 21306 596908 21374 596964
rect 21430 596908 21498 596964
rect 21554 596908 21622 596964
rect 21678 596908 39250 596964
rect 39306 596908 39374 596964
rect 39430 596908 39498 596964
rect 39554 596908 39622 596964
rect 39678 596908 57250 596964
rect 57306 596908 57374 596964
rect 57430 596908 57498 596964
rect 57554 596908 57622 596964
rect 57678 596908 75250 596964
rect 75306 596908 75374 596964
rect 75430 596908 75498 596964
rect 75554 596908 75622 596964
rect 75678 596908 93250 596964
rect 93306 596908 93374 596964
rect 93430 596908 93498 596964
rect 93554 596908 93622 596964
rect 93678 596908 111250 596964
rect 111306 596908 111374 596964
rect 111430 596908 111498 596964
rect 111554 596908 111622 596964
rect 111678 596908 129250 596964
rect 129306 596908 129374 596964
rect 129430 596908 129498 596964
rect 129554 596908 129622 596964
rect 129678 596908 147250 596964
rect 147306 596908 147374 596964
rect 147430 596908 147498 596964
rect 147554 596908 147622 596964
rect 147678 596908 165250 596964
rect 165306 596908 165374 596964
rect 165430 596908 165498 596964
rect 165554 596908 165622 596964
rect 165678 596908 183250 596964
rect 183306 596908 183374 596964
rect 183430 596908 183498 596964
rect 183554 596908 183622 596964
rect 183678 596908 201250 596964
rect 201306 596908 201374 596964
rect 201430 596908 201498 596964
rect 201554 596908 201622 596964
rect 201678 596908 219250 596964
rect 219306 596908 219374 596964
rect 219430 596908 219498 596964
rect 219554 596908 219622 596964
rect 219678 596908 237250 596964
rect 237306 596908 237374 596964
rect 237430 596908 237498 596964
rect 237554 596908 237622 596964
rect 237678 596908 255250 596964
rect 255306 596908 255374 596964
rect 255430 596908 255498 596964
rect 255554 596908 255622 596964
rect 255678 596908 273250 596964
rect 273306 596908 273374 596964
rect 273430 596908 273498 596964
rect 273554 596908 273622 596964
rect 273678 596908 291250 596964
rect 291306 596908 291374 596964
rect 291430 596908 291498 596964
rect 291554 596908 291622 596964
rect 291678 596908 309250 596964
rect 309306 596908 309374 596964
rect 309430 596908 309498 596964
rect 309554 596908 309622 596964
rect 309678 596908 327250 596964
rect 327306 596908 327374 596964
rect 327430 596908 327498 596964
rect 327554 596908 327622 596964
rect 327678 596908 345250 596964
rect 345306 596908 345374 596964
rect 345430 596908 345498 596964
rect 345554 596908 345622 596964
rect 345678 596908 363250 596964
rect 363306 596908 363374 596964
rect 363430 596908 363498 596964
rect 363554 596908 363622 596964
rect 363678 596908 381250 596964
rect 381306 596908 381374 596964
rect 381430 596908 381498 596964
rect 381554 596908 381622 596964
rect 381678 596908 399250 596964
rect 399306 596908 399374 596964
rect 399430 596908 399498 596964
rect 399554 596908 399622 596964
rect 399678 596908 417250 596964
rect 417306 596908 417374 596964
rect 417430 596908 417498 596964
rect 417554 596908 417622 596964
rect 417678 596908 435250 596964
rect 435306 596908 435374 596964
rect 435430 596908 435498 596964
rect 435554 596908 435622 596964
rect 435678 596908 453250 596964
rect 453306 596908 453374 596964
rect 453430 596908 453498 596964
rect 453554 596908 453622 596964
rect 453678 596908 471250 596964
rect 471306 596908 471374 596964
rect 471430 596908 471498 596964
rect 471554 596908 471622 596964
rect 471678 596908 489250 596964
rect 489306 596908 489374 596964
rect 489430 596908 489498 596964
rect 489554 596908 489622 596964
rect 489678 596908 507250 596964
rect 507306 596908 507374 596964
rect 507430 596908 507498 596964
rect 507554 596908 507622 596964
rect 507678 596908 525250 596964
rect 525306 596908 525374 596964
rect 525430 596908 525498 596964
rect 525554 596908 525622 596964
rect 525678 596908 543250 596964
rect 543306 596908 543374 596964
rect 543430 596908 543498 596964
rect 543554 596908 543622 596964
rect 543678 596908 561250 596964
rect 561306 596908 561374 596964
rect 561430 596908 561498 596964
rect 561554 596908 561622 596964
rect 561678 596908 579250 596964
rect 579306 596908 579374 596964
rect 579430 596908 579498 596964
rect 579554 596908 579622 596964
rect 579678 596908 596496 596964
rect 596552 596908 596620 596964
rect 596676 596908 596744 596964
rect 596800 596908 596868 596964
rect 596924 596908 597020 596964
rect -956 596840 597020 596908
rect -956 596784 -860 596840
rect -804 596784 -736 596840
rect -680 596784 -612 596840
rect -556 596784 -488 596840
rect -432 596784 3250 596840
rect 3306 596784 3374 596840
rect 3430 596784 3498 596840
rect 3554 596784 3622 596840
rect 3678 596784 21250 596840
rect 21306 596784 21374 596840
rect 21430 596784 21498 596840
rect 21554 596784 21622 596840
rect 21678 596784 39250 596840
rect 39306 596784 39374 596840
rect 39430 596784 39498 596840
rect 39554 596784 39622 596840
rect 39678 596784 57250 596840
rect 57306 596784 57374 596840
rect 57430 596784 57498 596840
rect 57554 596784 57622 596840
rect 57678 596784 75250 596840
rect 75306 596784 75374 596840
rect 75430 596784 75498 596840
rect 75554 596784 75622 596840
rect 75678 596784 93250 596840
rect 93306 596784 93374 596840
rect 93430 596784 93498 596840
rect 93554 596784 93622 596840
rect 93678 596784 111250 596840
rect 111306 596784 111374 596840
rect 111430 596784 111498 596840
rect 111554 596784 111622 596840
rect 111678 596784 129250 596840
rect 129306 596784 129374 596840
rect 129430 596784 129498 596840
rect 129554 596784 129622 596840
rect 129678 596784 147250 596840
rect 147306 596784 147374 596840
rect 147430 596784 147498 596840
rect 147554 596784 147622 596840
rect 147678 596784 165250 596840
rect 165306 596784 165374 596840
rect 165430 596784 165498 596840
rect 165554 596784 165622 596840
rect 165678 596784 183250 596840
rect 183306 596784 183374 596840
rect 183430 596784 183498 596840
rect 183554 596784 183622 596840
rect 183678 596784 201250 596840
rect 201306 596784 201374 596840
rect 201430 596784 201498 596840
rect 201554 596784 201622 596840
rect 201678 596784 219250 596840
rect 219306 596784 219374 596840
rect 219430 596784 219498 596840
rect 219554 596784 219622 596840
rect 219678 596784 237250 596840
rect 237306 596784 237374 596840
rect 237430 596784 237498 596840
rect 237554 596784 237622 596840
rect 237678 596784 255250 596840
rect 255306 596784 255374 596840
rect 255430 596784 255498 596840
rect 255554 596784 255622 596840
rect 255678 596784 273250 596840
rect 273306 596784 273374 596840
rect 273430 596784 273498 596840
rect 273554 596784 273622 596840
rect 273678 596784 291250 596840
rect 291306 596784 291374 596840
rect 291430 596784 291498 596840
rect 291554 596784 291622 596840
rect 291678 596784 309250 596840
rect 309306 596784 309374 596840
rect 309430 596784 309498 596840
rect 309554 596784 309622 596840
rect 309678 596784 327250 596840
rect 327306 596784 327374 596840
rect 327430 596784 327498 596840
rect 327554 596784 327622 596840
rect 327678 596784 345250 596840
rect 345306 596784 345374 596840
rect 345430 596784 345498 596840
rect 345554 596784 345622 596840
rect 345678 596784 363250 596840
rect 363306 596784 363374 596840
rect 363430 596784 363498 596840
rect 363554 596784 363622 596840
rect 363678 596784 381250 596840
rect 381306 596784 381374 596840
rect 381430 596784 381498 596840
rect 381554 596784 381622 596840
rect 381678 596784 399250 596840
rect 399306 596784 399374 596840
rect 399430 596784 399498 596840
rect 399554 596784 399622 596840
rect 399678 596784 417250 596840
rect 417306 596784 417374 596840
rect 417430 596784 417498 596840
rect 417554 596784 417622 596840
rect 417678 596784 435250 596840
rect 435306 596784 435374 596840
rect 435430 596784 435498 596840
rect 435554 596784 435622 596840
rect 435678 596784 453250 596840
rect 453306 596784 453374 596840
rect 453430 596784 453498 596840
rect 453554 596784 453622 596840
rect 453678 596784 471250 596840
rect 471306 596784 471374 596840
rect 471430 596784 471498 596840
rect 471554 596784 471622 596840
rect 471678 596784 489250 596840
rect 489306 596784 489374 596840
rect 489430 596784 489498 596840
rect 489554 596784 489622 596840
rect 489678 596784 507250 596840
rect 507306 596784 507374 596840
rect 507430 596784 507498 596840
rect 507554 596784 507622 596840
rect 507678 596784 525250 596840
rect 525306 596784 525374 596840
rect 525430 596784 525498 596840
rect 525554 596784 525622 596840
rect 525678 596784 543250 596840
rect 543306 596784 543374 596840
rect 543430 596784 543498 596840
rect 543554 596784 543622 596840
rect 543678 596784 561250 596840
rect 561306 596784 561374 596840
rect 561430 596784 561498 596840
rect 561554 596784 561622 596840
rect 561678 596784 579250 596840
rect 579306 596784 579374 596840
rect 579430 596784 579498 596840
rect 579554 596784 579622 596840
rect 579678 596784 596496 596840
rect 596552 596784 596620 596840
rect 596676 596784 596744 596840
rect 596800 596784 596868 596840
rect 596924 596784 597020 596840
rect -956 596688 597020 596784
rect -1916 586350 597980 586446
rect -1916 586294 -1820 586350
rect -1764 586294 -1696 586350
rect -1640 586294 -1572 586350
rect -1516 586294 -1448 586350
rect -1392 586294 6970 586350
rect 7026 586294 7094 586350
rect 7150 586294 7218 586350
rect 7274 586294 7342 586350
rect 7398 586294 24970 586350
rect 25026 586294 25094 586350
rect 25150 586294 25218 586350
rect 25274 586294 25342 586350
rect 25398 586294 42970 586350
rect 43026 586294 43094 586350
rect 43150 586294 43218 586350
rect 43274 586294 43342 586350
rect 43398 586294 60970 586350
rect 61026 586294 61094 586350
rect 61150 586294 61218 586350
rect 61274 586294 61342 586350
rect 61398 586294 78970 586350
rect 79026 586294 79094 586350
rect 79150 586294 79218 586350
rect 79274 586294 79342 586350
rect 79398 586294 96970 586350
rect 97026 586294 97094 586350
rect 97150 586294 97218 586350
rect 97274 586294 97342 586350
rect 97398 586294 114970 586350
rect 115026 586294 115094 586350
rect 115150 586294 115218 586350
rect 115274 586294 115342 586350
rect 115398 586294 132970 586350
rect 133026 586294 133094 586350
rect 133150 586294 133218 586350
rect 133274 586294 133342 586350
rect 133398 586294 150970 586350
rect 151026 586294 151094 586350
rect 151150 586294 151218 586350
rect 151274 586294 151342 586350
rect 151398 586294 168970 586350
rect 169026 586294 169094 586350
rect 169150 586294 169218 586350
rect 169274 586294 169342 586350
rect 169398 586294 186970 586350
rect 187026 586294 187094 586350
rect 187150 586294 187218 586350
rect 187274 586294 187342 586350
rect 187398 586294 204970 586350
rect 205026 586294 205094 586350
rect 205150 586294 205218 586350
rect 205274 586294 205342 586350
rect 205398 586294 222970 586350
rect 223026 586294 223094 586350
rect 223150 586294 223218 586350
rect 223274 586294 223342 586350
rect 223398 586294 240970 586350
rect 241026 586294 241094 586350
rect 241150 586294 241218 586350
rect 241274 586294 241342 586350
rect 241398 586294 258970 586350
rect 259026 586294 259094 586350
rect 259150 586294 259218 586350
rect 259274 586294 259342 586350
rect 259398 586294 276970 586350
rect 277026 586294 277094 586350
rect 277150 586294 277218 586350
rect 277274 586294 277342 586350
rect 277398 586294 294970 586350
rect 295026 586294 295094 586350
rect 295150 586294 295218 586350
rect 295274 586294 295342 586350
rect 295398 586294 312970 586350
rect 313026 586294 313094 586350
rect 313150 586294 313218 586350
rect 313274 586294 313342 586350
rect 313398 586294 330970 586350
rect 331026 586294 331094 586350
rect 331150 586294 331218 586350
rect 331274 586294 331342 586350
rect 331398 586294 348970 586350
rect 349026 586294 349094 586350
rect 349150 586294 349218 586350
rect 349274 586294 349342 586350
rect 349398 586294 366970 586350
rect 367026 586294 367094 586350
rect 367150 586294 367218 586350
rect 367274 586294 367342 586350
rect 367398 586294 384970 586350
rect 385026 586294 385094 586350
rect 385150 586294 385218 586350
rect 385274 586294 385342 586350
rect 385398 586294 402970 586350
rect 403026 586294 403094 586350
rect 403150 586294 403218 586350
rect 403274 586294 403342 586350
rect 403398 586294 420970 586350
rect 421026 586294 421094 586350
rect 421150 586294 421218 586350
rect 421274 586294 421342 586350
rect 421398 586294 438970 586350
rect 439026 586294 439094 586350
rect 439150 586294 439218 586350
rect 439274 586294 439342 586350
rect 439398 586294 456970 586350
rect 457026 586294 457094 586350
rect 457150 586294 457218 586350
rect 457274 586294 457342 586350
rect 457398 586294 474970 586350
rect 475026 586294 475094 586350
rect 475150 586294 475218 586350
rect 475274 586294 475342 586350
rect 475398 586294 492970 586350
rect 493026 586294 493094 586350
rect 493150 586294 493218 586350
rect 493274 586294 493342 586350
rect 493398 586294 510970 586350
rect 511026 586294 511094 586350
rect 511150 586294 511218 586350
rect 511274 586294 511342 586350
rect 511398 586294 528970 586350
rect 529026 586294 529094 586350
rect 529150 586294 529218 586350
rect 529274 586294 529342 586350
rect 529398 586294 546970 586350
rect 547026 586294 547094 586350
rect 547150 586294 547218 586350
rect 547274 586294 547342 586350
rect 547398 586294 564970 586350
rect 565026 586294 565094 586350
rect 565150 586294 565218 586350
rect 565274 586294 565342 586350
rect 565398 586294 582970 586350
rect 583026 586294 583094 586350
rect 583150 586294 583218 586350
rect 583274 586294 583342 586350
rect 583398 586294 597456 586350
rect 597512 586294 597580 586350
rect 597636 586294 597704 586350
rect 597760 586294 597828 586350
rect 597884 586294 597980 586350
rect -1916 586226 597980 586294
rect -1916 586170 -1820 586226
rect -1764 586170 -1696 586226
rect -1640 586170 -1572 586226
rect -1516 586170 -1448 586226
rect -1392 586170 6970 586226
rect 7026 586170 7094 586226
rect 7150 586170 7218 586226
rect 7274 586170 7342 586226
rect 7398 586170 24970 586226
rect 25026 586170 25094 586226
rect 25150 586170 25218 586226
rect 25274 586170 25342 586226
rect 25398 586170 42970 586226
rect 43026 586170 43094 586226
rect 43150 586170 43218 586226
rect 43274 586170 43342 586226
rect 43398 586170 60970 586226
rect 61026 586170 61094 586226
rect 61150 586170 61218 586226
rect 61274 586170 61342 586226
rect 61398 586170 78970 586226
rect 79026 586170 79094 586226
rect 79150 586170 79218 586226
rect 79274 586170 79342 586226
rect 79398 586170 96970 586226
rect 97026 586170 97094 586226
rect 97150 586170 97218 586226
rect 97274 586170 97342 586226
rect 97398 586170 114970 586226
rect 115026 586170 115094 586226
rect 115150 586170 115218 586226
rect 115274 586170 115342 586226
rect 115398 586170 132970 586226
rect 133026 586170 133094 586226
rect 133150 586170 133218 586226
rect 133274 586170 133342 586226
rect 133398 586170 150970 586226
rect 151026 586170 151094 586226
rect 151150 586170 151218 586226
rect 151274 586170 151342 586226
rect 151398 586170 168970 586226
rect 169026 586170 169094 586226
rect 169150 586170 169218 586226
rect 169274 586170 169342 586226
rect 169398 586170 186970 586226
rect 187026 586170 187094 586226
rect 187150 586170 187218 586226
rect 187274 586170 187342 586226
rect 187398 586170 204970 586226
rect 205026 586170 205094 586226
rect 205150 586170 205218 586226
rect 205274 586170 205342 586226
rect 205398 586170 222970 586226
rect 223026 586170 223094 586226
rect 223150 586170 223218 586226
rect 223274 586170 223342 586226
rect 223398 586170 240970 586226
rect 241026 586170 241094 586226
rect 241150 586170 241218 586226
rect 241274 586170 241342 586226
rect 241398 586170 258970 586226
rect 259026 586170 259094 586226
rect 259150 586170 259218 586226
rect 259274 586170 259342 586226
rect 259398 586170 276970 586226
rect 277026 586170 277094 586226
rect 277150 586170 277218 586226
rect 277274 586170 277342 586226
rect 277398 586170 294970 586226
rect 295026 586170 295094 586226
rect 295150 586170 295218 586226
rect 295274 586170 295342 586226
rect 295398 586170 312970 586226
rect 313026 586170 313094 586226
rect 313150 586170 313218 586226
rect 313274 586170 313342 586226
rect 313398 586170 330970 586226
rect 331026 586170 331094 586226
rect 331150 586170 331218 586226
rect 331274 586170 331342 586226
rect 331398 586170 348970 586226
rect 349026 586170 349094 586226
rect 349150 586170 349218 586226
rect 349274 586170 349342 586226
rect 349398 586170 366970 586226
rect 367026 586170 367094 586226
rect 367150 586170 367218 586226
rect 367274 586170 367342 586226
rect 367398 586170 384970 586226
rect 385026 586170 385094 586226
rect 385150 586170 385218 586226
rect 385274 586170 385342 586226
rect 385398 586170 402970 586226
rect 403026 586170 403094 586226
rect 403150 586170 403218 586226
rect 403274 586170 403342 586226
rect 403398 586170 420970 586226
rect 421026 586170 421094 586226
rect 421150 586170 421218 586226
rect 421274 586170 421342 586226
rect 421398 586170 438970 586226
rect 439026 586170 439094 586226
rect 439150 586170 439218 586226
rect 439274 586170 439342 586226
rect 439398 586170 456970 586226
rect 457026 586170 457094 586226
rect 457150 586170 457218 586226
rect 457274 586170 457342 586226
rect 457398 586170 474970 586226
rect 475026 586170 475094 586226
rect 475150 586170 475218 586226
rect 475274 586170 475342 586226
rect 475398 586170 492970 586226
rect 493026 586170 493094 586226
rect 493150 586170 493218 586226
rect 493274 586170 493342 586226
rect 493398 586170 510970 586226
rect 511026 586170 511094 586226
rect 511150 586170 511218 586226
rect 511274 586170 511342 586226
rect 511398 586170 528970 586226
rect 529026 586170 529094 586226
rect 529150 586170 529218 586226
rect 529274 586170 529342 586226
rect 529398 586170 546970 586226
rect 547026 586170 547094 586226
rect 547150 586170 547218 586226
rect 547274 586170 547342 586226
rect 547398 586170 564970 586226
rect 565026 586170 565094 586226
rect 565150 586170 565218 586226
rect 565274 586170 565342 586226
rect 565398 586170 582970 586226
rect 583026 586170 583094 586226
rect 583150 586170 583218 586226
rect 583274 586170 583342 586226
rect 583398 586170 597456 586226
rect 597512 586170 597580 586226
rect 597636 586170 597704 586226
rect 597760 586170 597828 586226
rect 597884 586170 597980 586226
rect -1916 586102 597980 586170
rect -1916 586046 -1820 586102
rect -1764 586046 -1696 586102
rect -1640 586046 -1572 586102
rect -1516 586046 -1448 586102
rect -1392 586046 6970 586102
rect 7026 586046 7094 586102
rect 7150 586046 7218 586102
rect 7274 586046 7342 586102
rect 7398 586046 24970 586102
rect 25026 586046 25094 586102
rect 25150 586046 25218 586102
rect 25274 586046 25342 586102
rect 25398 586046 42970 586102
rect 43026 586046 43094 586102
rect 43150 586046 43218 586102
rect 43274 586046 43342 586102
rect 43398 586046 60970 586102
rect 61026 586046 61094 586102
rect 61150 586046 61218 586102
rect 61274 586046 61342 586102
rect 61398 586046 78970 586102
rect 79026 586046 79094 586102
rect 79150 586046 79218 586102
rect 79274 586046 79342 586102
rect 79398 586046 96970 586102
rect 97026 586046 97094 586102
rect 97150 586046 97218 586102
rect 97274 586046 97342 586102
rect 97398 586046 114970 586102
rect 115026 586046 115094 586102
rect 115150 586046 115218 586102
rect 115274 586046 115342 586102
rect 115398 586046 132970 586102
rect 133026 586046 133094 586102
rect 133150 586046 133218 586102
rect 133274 586046 133342 586102
rect 133398 586046 150970 586102
rect 151026 586046 151094 586102
rect 151150 586046 151218 586102
rect 151274 586046 151342 586102
rect 151398 586046 168970 586102
rect 169026 586046 169094 586102
rect 169150 586046 169218 586102
rect 169274 586046 169342 586102
rect 169398 586046 186970 586102
rect 187026 586046 187094 586102
rect 187150 586046 187218 586102
rect 187274 586046 187342 586102
rect 187398 586046 204970 586102
rect 205026 586046 205094 586102
rect 205150 586046 205218 586102
rect 205274 586046 205342 586102
rect 205398 586046 222970 586102
rect 223026 586046 223094 586102
rect 223150 586046 223218 586102
rect 223274 586046 223342 586102
rect 223398 586046 240970 586102
rect 241026 586046 241094 586102
rect 241150 586046 241218 586102
rect 241274 586046 241342 586102
rect 241398 586046 258970 586102
rect 259026 586046 259094 586102
rect 259150 586046 259218 586102
rect 259274 586046 259342 586102
rect 259398 586046 276970 586102
rect 277026 586046 277094 586102
rect 277150 586046 277218 586102
rect 277274 586046 277342 586102
rect 277398 586046 294970 586102
rect 295026 586046 295094 586102
rect 295150 586046 295218 586102
rect 295274 586046 295342 586102
rect 295398 586046 312970 586102
rect 313026 586046 313094 586102
rect 313150 586046 313218 586102
rect 313274 586046 313342 586102
rect 313398 586046 330970 586102
rect 331026 586046 331094 586102
rect 331150 586046 331218 586102
rect 331274 586046 331342 586102
rect 331398 586046 348970 586102
rect 349026 586046 349094 586102
rect 349150 586046 349218 586102
rect 349274 586046 349342 586102
rect 349398 586046 366970 586102
rect 367026 586046 367094 586102
rect 367150 586046 367218 586102
rect 367274 586046 367342 586102
rect 367398 586046 384970 586102
rect 385026 586046 385094 586102
rect 385150 586046 385218 586102
rect 385274 586046 385342 586102
rect 385398 586046 402970 586102
rect 403026 586046 403094 586102
rect 403150 586046 403218 586102
rect 403274 586046 403342 586102
rect 403398 586046 420970 586102
rect 421026 586046 421094 586102
rect 421150 586046 421218 586102
rect 421274 586046 421342 586102
rect 421398 586046 438970 586102
rect 439026 586046 439094 586102
rect 439150 586046 439218 586102
rect 439274 586046 439342 586102
rect 439398 586046 456970 586102
rect 457026 586046 457094 586102
rect 457150 586046 457218 586102
rect 457274 586046 457342 586102
rect 457398 586046 474970 586102
rect 475026 586046 475094 586102
rect 475150 586046 475218 586102
rect 475274 586046 475342 586102
rect 475398 586046 492970 586102
rect 493026 586046 493094 586102
rect 493150 586046 493218 586102
rect 493274 586046 493342 586102
rect 493398 586046 510970 586102
rect 511026 586046 511094 586102
rect 511150 586046 511218 586102
rect 511274 586046 511342 586102
rect 511398 586046 528970 586102
rect 529026 586046 529094 586102
rect 529150 586046 529218 586102
rect 529274 586046 529342 586102
rect 529398 586046 546970 586102
rect 547026 586046 547094 586102
rect 547150 586046 547218 586102
rect 547274 586046 547342 586102
rect 547398 586046 564970 586102
rect 565026 586046 565094 586102
rect 565150 586046 565218 586102
rect 565274 586046 565342 586102
rect 565398 586046 582970 586102
rect 583026 586046 583094 586102
rect 583150 586046 583218 586102
rect 583274 586046 583342 586102
rect 583398 586046 597456 586102
rect 597512 586046 597580 586102
rect 597636 586046 597704 586102
rect 597760 586046 597828 586102
rect 597884 586046 597980 586102
rect -1916 585978 597980 586046
rect -1916 585922 -1820 585978
rect -1764 585922 -1696 585978
rect -1640 585922 -1572 585978
rect -1516 585922 -1448 585978
rect -1392 585922 6970 585978
rect 7026 585922 7094 585978
rect 7150 585922 7218 585978
rect 7274 585922 7342 585978
rect 7398 585922 24970 585978
rect 25026 585922 25094 585978
rect 25150 585922 25218 585978
rect 25274 585922 25342 585978
rect 25398 585922 42970 585978
rect 43026 585922 43094 585978
rect 43150 585922 43218 585978
rect 43274 585922 43342 585978
rect 43398 585922 60970 585978
rect 61026 585922 61094 585978
rect 61150 585922 61218 585978
rect 61274 585922 61342 585978
rect 61398 585922 78970 585978
rect 79026 585922 79094 585978
rect 79150 585922 79218 585978
rect 79274 585922 79342 585978
rect 79398 585922 96970 585978
rect 97026 585922 97094 585978
rect 97150 585922 97218 585978
rect 97274 585922 97342 585978
rect 97398 585922 114970 585978
rect 115026 585922 115094 585978
rect 115150 585922 115218 585978
rect 115274 585922 115342 585978
rect 115398 585922 132970 585978
rect 133026 585922 133094 585978
rect 133150 585922 133218 585978
rect 133274 585922 133342 585978
rect 133398 585922 150970 585978
rect 151026 585922 151094 585978
rect 151150 585922 151218 585978
rect 151274 585922 151342 585978
rect 151398 585922 168970 585978
rect 169026 585922 169094 585978
rect 169150 585922 169218 585978
rect 169274 585922 169342 585978
rect 169398 585922 186970 585978
rect 187026 585922 187094 585978
rect 187150 585922 187218 585978
rect 187274 585922 187342 585978
rect 187398 585922 204970 585978
rect 205026 585922 205094 585978
rect 205150 585922 205218 585978
rect 205274 585922 205342 585978
rect 205398 585922 222970 585978
rect 223026 585922 223094 585978
rect 223150 585922 223218 585978
rect 223274 585922 223342 585978
rect 223398 585922 240970 585978
rect 241026 585922 241094 585978
rect 241150 585922 241218 585978
rect 241274 585922 241342 585978
rect 241398 585922 258970 585978
rect 259026 585922 259094 585978
rect 259150 585922 259218 585978
rect 259274 585922 259342 585978
rect 259398 585922 276970 585978
rect 277026 585922 277094 585978
rect 277150 585922 277218 585978
rect 277274 585922 277342 585978
rect 277398 585922 294970 585978
rect 295026 585922 295094 585978
rect 295150 585922 295218 585978
rect 295274 585922 295342 585978
rect 295398 585922 312970 585978
rect 313026 585922 313094 585978
rect 313150 585922 313218 585978
rect 313274 585922 313342 585978
rect 313398 585922 330970 585978
rect 331026 585922 331094 585978
rect 331150 585922 331218 585978
rect 331274 585922 331342 585978
rect 331398 585922 348970 585978
rect 349026 585922 349094 585978
rect 349150 585922 349218 585978
rect 349274 585922 349342 585978
rect 349398 585922 366970 585978
rect 367026 585922 367094 585978
rect 367150 585922 367218 585978
rect 367274 585922 367342 585978
rect 367398 585922 384970 585978
rect 385026 585922 385094 585978
rect 385150 585922 385218 585978
rect 385274 585922 385342 585978
rect 385398 585922 402970 585978
rect 403026 585922 403094 585978
rect 403150 585922 403218 585978
rect 403274 585922 403342 585978
rect 403398 585922 420970 585978
rect 421026 585922 421094 585978
rect 421150 585922 421218 585978
rect 421274 585922 421342 585978
rect 421398 585922 438970 585978
rect 439026 585922 439094 585978
rect 439150 585922 439218 585978
rect 439274 585922 439342 585978
rect 439398 585922 456970 585978
rect 457026 585922 457094 585978
rect 457150 585922 457218 585978
rect 457274 585922 457342 585978
rect 457398 585922 474970 585978
rect 475026 585922 475094 585978
rect 475150 585922 475218 585978
rect 475274 585922 475342 585978
rect 475398 585922 492970 585978
rect 493026 585922 493094 585978
rect 493150 585922 493218 585978
rect 493274 585922 493342 585978
rect 493398 585922 510970 585978
rect 511026 585922 511094 585978
rect 511150 585922 511218 585978
rect 511274 585922 511342 585978
rect 511398 585922 528970 585978
rect 529026 585922 529094 585978
rect 529150 585922 529218 585978
rect 529274 585922 529342 585978
rect 529398 585922 546970 585978
rect 547026 585922 547094 585978
rect 547150 585922 547218 585978
rect 547274 585922 547342 585978
rect 547398 585922 564970 585978
rect 565026 585922 565094 585978
rect 565150 585922 565218 585978
rect 565274 585922 565342 585978
rect 565398 585922 582970 585978
rect 583026 585922 583094 585978
rect 583150 585922 583218 585978
rect 583274 585922 583342 585978
rect 583398 585922 597456 585978
rect 597512 585922 597580 585978
rect 597636 585922 597704 585978
rect 597760 585922 597828 585978
rect 597884 585922 597980 585978
rect -1916 585826 597980 585922
rect -1916 580350 597980 580446
rect -1916 580294 -860 580350
rect -804 580294 -736 580350
rect -680 580294 -612 580350
rect -556 580294 -488 580350
rect -432 580294 3250 580350
rect 3306 580294 3374 580350
rect 3430 580294 3498 580350
rect 3554 580294 3622 580350
rect 3678 580294 21250 580350
rect 21306 580294 21374 580350
rect 21430 580294 21498 580350
rect 21554 580294 21622 580350
rect 21678 580294 39250 580350
rect 39306 580294 39374 580350
rect 39430 580294 39498 580350
rect 39554 580294 39622 580350
rect 39678 580294 57250 580350
rect 57306 580294 57374 580350
rect 57430 580294 57498 580350
rect 57554 580294 57622 580350
rect 57678 580294 75250 580350
rect 75306 580294 75374 580350
rect 75430 580294 75498 580350
rect 75554 580294 75622 580350
rect 75678 580294 93250 580350
rect 93306 580294 93374 580350
rect 93430 580294 93498 580350
rect 93554 580294 93622 580350
rect 93678 580294 111250 580350
rect 111306 580294 111374 580350
rect 111430 580294 111498 580350
rect 111554 580294 111622 580350
rect 111678 580294 129250 580350
rect 129306 580294 129374 580350
rect 129430 580294 129498 580350
rect 129554 580294 129622 580350
rect 129678 580294 147250 580350
rect 147306 580294 147374 580350
rect 147430 580294 147498 580350
rect 147554 580294 147622 580350
rect 147678 580294 165250 580350
rect 165306 580294 165374 580350
rect 165430 580294 165498 580350
rect 165554 580294 165622 580350
rect 165678 580294 183250 580350
rect 183306 580294 183374 580350
rect 183430 580294 183498 580350
rect 183554 580294 183622 580350
rect 183678 580294 201250 580350
rect 201306 580294 201374 580350
rect 201430 580294 201498 580350
rect 201554 580294 201622 580350
rect 201678 580294 219250 580350
rect 219306 580294 219374 580350
rect 219430 580294 219498 580350
rect 219554 580294 219622 580350
rect 219678 580294 237250 580350
rect 237306 580294 237374 580350
rect 237430 580294 237498 580350
rect 237554 580294 237622 580350
rect 237678 580294 255250 580350
rect 255306 580294 255374 580350
rect 255430 580294 255498 580350
rect 255554 580294 255622 580350
rect 255678 580294 273250 580350
rect 273306 580294 273374 580350
rect 273430 580294 273498 580350
rect 273554 580294 273622 580350
rect 273678 580294 291250 580350
rect 291306 580294 291374 580350
rect 291430 580294 291498 580350
rect 291554 580294 291622 580350
rect 291678 580294 309250 580350
rect 309306 580294 309374 580350
rect 309430 580294 309498 580350
rect 309554 580294 309622 580350
rect 309678 580294 327250 580350
rect 327306 580294 327374 580350
rect 327430 580294 327498 580350
rect 327554 580294 327622 580350
rect 327678 580294 345250 580350
rect 345306 580294 345374 580350
rect 345430 580294 345498 580350
rect 345554 580294 345622 580350
rect 345678 580294 363250 580350
rect 363306 580294 363374 580350
rect 363430 580294 363498 580350
rect 363554 580294 363622 580350
rect 363678 580294 381250 580350
rect 381306 580294 381374 580350
rect 381430 580294 381498 580350
rect 381554 580294 381622 580350
rect 381678 580294 399250 580350
rect 399306 580294 399374 580350
rect 399430 580294 399498 580350
rect 399554 580294 399622 580350
rect 399678 580294 417250 580350
rect 417306 580294 417374 580350
rect 417430 580294 417498 580350
rect 417554 580294 417622 580350
rect 417678 580294 435250 580350
rect 435306 580294 435374 580350
rect 435430 580294 435498 580350
rect 435554 580294 435622 580350
rect 435678 580294 453250 580350
rect 453306 580294 453374 580350
rect 453430 580294 453498 580350
rect 453554 580294 453622 580350
rect 453678 580294 471250 580350
rect 471306 580294 471374 580350
rect 471430 580294 471498 580350
rect 471554 580294 471622 580350
rect 471678 580294 489250 580350
rect 489306 580294 489374 580350
rect 489430 580294 489498 580350
rect 489554 580294 489622 580350
rect 489678 580294 507250 580350
rect 507306 580294 507374 580350
rect 507430 580294 507498 580350
rect 507554 580294 507622 580350
rect 507678 580294 525250 580350
rect 525306 580294 525374 580350
rect 525430 580294 525498 580350
rect 525554 580294 525622 580350
rect 525678 580294 543250 580350
rect 543306 580294 543374 580350
rect 543430 580294 543498 580350
rect 543554 580294 543622 580350
rect 543678 580294 561250 580350
rect 561306 580294 561374 580350
rect 561430 580294 561498 580350
rect 561554 580294 561622 580350
rect 561678 580294 579250 580350
rect 579306 580294 579374 580350
rect 579430 580294 579498 580350
rect 579554 580294 579622 580350
rect 579678 580294 596496 580350
rect 596552 580294 596620 580350
rect 596676 580294 596744 580350
rect 596800 580294 596868 580350
rect 596924 580294 597980 580350
rect -1916 580226 597980 580294
rect -1916 580170 -860 580226
rect -804 580170 -736 580226
rect -680 580170 -612 580226
rect -556 580170 -488 580226
rect -432 580170 3250 580226
rect 3306 580170 3374 580226
rect 3430 580170 3498 580226
rect 3554 580170 3622 580226
rect 3678 580170 21250 580226
rect 21306 580170 21374 580226
rect 21430 580170 21498 580226
rect 21554 580170 21622 580226
rect 21678 580170 39250 580226
rect 39306 580170 39374 580226
rect 39430 580170 39498 580226
rect 39554 580170 39622 580226
rect 39678 580170 57250 580226
rect 57306 580170 57374 580226
rect 57430 580170 57498 580226
rect 57554 580170 57622 580226
rect 57678 580170 75250 580226
rect 75306 580170 75374 580226
rect 75430 580170 75498 580226
rect 75554 580170 75622 580226
rect 75678 580170 93250 580226
rect 93306 580170 93374 580226
rect 93430 580170 93498 580226
rect 93554 580170 93622 580226
rect 93678 580170 111250 580226
rect 111306 580170 111374 580226
rect 111430 580170 111498 580226
rect 111554 580170 111622 580226
rect 111678 580170 129250 580226
rect 129306 580170 129374 580226
rect 129430 580170 129498 580226
rect 129554 580170 129622 580226
rect 129678 580170 147250 580226
rect 147306 580170 147374 580226
rect 147430 580170 147498 580226
rect 147554 580170 147622 580226
rect 147678 580170 165250 580226
rect 165306 580170 165374 580226
rect 165430 580170 165498 580226
rect 165554 580170 165622 580226
rect 165678 580170 183250 580226
rect 183306 580170 183374 580226
rect 183430 580170 183498 580226
rect 183554 580170 183622 580226
rect 183678 580170 201250 580226
rect 201306 580170 201374 580226
rect 201430 580170 201498 580226
rect 201554 580170 201622 580226
rect 201678 580170 219250 580226
rect 219306 580170 219374 580226
rect 219430 580170 219498 580226
rect 219554 580170 219622 580226
rect 219678 580170 237250 580226
rect 237306 580170 237374 580226
rect 237430 580170 237498 580226
rect 237554 580170 237622 580226
rect 237678 580170 255250 580226
rect 255306 580170 255374 580226
rect 255430 580170 255498 580226
rect 255554 580170 255622 580226
rect 255678 580170 273250 580226
rect 273306 580170 273374 580226
rect 273430 580170 273498 580226
rect 273554 580170 273622 580226
rect 273678 580170 291250 580226
rect 291306 580170 291374 580226
rect 291430 580170 291498 580226
rect 291554 580170 291622 580226
rect 291678 580170 309250 580226
rect 309306 580170 309374 580226
rect 309430 580170 309498 580226
rect 309554 580170 309622 580226
rect 309678 580170 327250 580226
rect 327306 580170 327374 580226
rect 327430 580170 327498 580226
rect 327554 580170 327622 580226
rect 327678 580170 345250 580226
rect 345306 580170 345374 580226
rect 345430 580170 345498 580226
rect 345554 580170 345622 580226
rect 345678 580170 363250 580226
rect 363306 580170 363374 580226
rect 363430 580170 363498 580226
rect 363554 580170 363622 580226
rect 363678 580170 381250 580226
rect 381306 580170 381374 580226
rect 381430 580170 381498 580226
rect 381554 580170 381622 580226
rect 381678 580170 399250 580226
rect 399306 580170 399374 580226
rect 399430 580170 399498 580226
rect 399554 580170 399622 580226
rect 399678 580170 417250 580226
rect 417306 580170 417374 580226
rect 417430 580170 417498 580226
rect 417554 580170 417622 580226
rect 417678 580170 435250 580226
rect 435306 580170 435374 580226
rect 435430 580170 435498 580226
rect 435554 580170 435622 580226
rect 435678 580170 453250 580226
rect 453306 580170 453374 580226
rect 453430 580170 453498 580226
rect 453554 580170 453622 580226
rect 453678 580170 471250 580226
rect 471306 580170 471374 580226
rect 471430 580170 471498 580226
rect 471554 580170 471622 580226
rect 471678 580170 489250 580226
rect 489306 580170 489374 580226
rect 489430 580170 489498 580226
rect 489554 580170 489622 580226
rect 489678 580170 507250 580226
rect 507306 580170 507374 580226
rect 507430 580170 507498 580226
rect 507554 580170 507622 580226
rect 507678 580170 525250 580226
rect 525306 580170 525374 580226
rect 525430 580170 525498 580226
rect 525554 580170 525622 580226
rect 525678 580170 543250 580226
rect 543306 580170 543374 580226
rect 543430 580170 543498 580226
rect 543554 580170 543622 580226
rect 543678 580170 561250 580226
rect 561306 580170 561374 580226
rect 561430 580170 561498 580226
rect 561554 580170 561622 580226
rect 561678 580170 579250 580226
rect 579306 580170 579374 580226
rect 579430 580170 579498 580226
rect 579554 580170 579622 580226
rect 579678 580170 596496 580226
rect 596552 580170 596620 580226
rect 596676 580170 596744 580226
rect 596800 580170 596868 580226
rect 596924 580170 597980 580226
rect -1916 580102 597980 580170
rect -1916 580046 -860 580102
rect -804 580046 -736 580102
rect -680 580046 -612 580102
rect -556 580046 -488 580102
rect -432 580046 3250 580102
rect 3306 580046 3374 580102
rect 3430 580046 3498 580102
rect 3554 580046 3622 580102
rect 3678 580046 21250 580102
rect 21306 580046 21374 580102
rect 21430 580046 21498 580102
rect 21554 580046 21622 580102
rect 21678 580046 39250 580102
rect 39306 580046 39374 580102
rect 39430 580046 39498 580102
rect 39554 580046 39622 580102
rect 39678 580046 57250 580102
rect 57306 580046 57374 580102
rect 57430 580046 57498 580102
rect 57554 580046 57622 580102
rect 57678 580046 75250 580102
rect 75306 580046 75374 580102
rect 75430 580046 75498 580102
rect 75554 580046 75622 580102
rect 75678 580046 93250 580102
rect 93306 580046 93374 580102
rect 93430 580046 93498 580102
rect 93554 580046 93622 580102
rect 93678 580046 111250 580102
rect 111306 580046 111374 580102
rect 111430 580046 111498 580102
rect 111554 580046 111622 580102
rect 111678 580046 129250 580102
rect 129306 580046 129374 580102
rect 129430 580046 129498 580102
rect 129554 580046 129622 580102
rect 129678 580046 147250 580102
rect 147306 580046 147374 580102
rect 147430 580046 147498 580102
rect 147554 580046 147622 580102
rect 147678 580046 165250 580102
rect 165306 580046 165374 580102
rect 165430 580046 165498 580102
rect 165554 580046 165622 580102
rect 165678 580046 183250 580102
rect 183306 580046 183374 580102
rect 183430 580046 183498 580102
rect 183554 580046 183622 580102
rect 183678 580046 201250 580102
rect 201306 580046 201374 580102
rect 201430 580046 201498 580102
rect 201554 580046 201622 580102
rect 201678 580046 219250 580102
rect 219306 580046 219374 580102
rect 219430 580046 219498 580102
rect 219554 580046 219622 580102
rect 219678 580046 237250 580102
rect 237306 580046 237374 580102
rect 237430 580046 237498 580102
rect 237554 580046 237622 580102
rect 237678 580046 255250 580102
rect 255306 580046 255374 580102
rect 255430 580046 255498 580102
rect 255554 580046 255622 580102
rect 255678 580046 273250 580102
rect 273306 580046 273374 580102
rect 273430 580046 273498 580102
rect 273554 580046 273622 580102
rect 273678 580046 291250 580102
rect 291306 580046 291374 580102
rect 291430 580046 291498 580102
rect 291554 580046 291622 580102
rect 291678 580046 309250 580102
rect 309306 580046 309374 580102
rect 309430 580046 309498 580102
rect 309554 580046 309622 580102
rect 309678 580046 327250 580102
rect 327306 580046 327374 580102
rect 327430 580046 327498 580102
rect 327554 580046 327622 580102
rect 327678 580046 345250 580102
rect 345306 580046 345374 580102
rect 345430 580046 345498 580102
rect 345554 580046 345622 580102
rect 345678 580046 363250 580102
rect 363306 580046 363374 580102
rect 363430 580046 363498 580102
rect 363554 580046 363622 580102
rect 363678 580046 381250 580102
rect 381306 580046 381374 580102
rect 381430 580046 381498 580102
rect 381554 580046 381622 580102
rect 381678 580046 399250 580102
rect 399306 580046 399374 580102
rect 399430 580046 399498 580102
rect 399554 580046 399622 580102
rect 399678 580046 417250 580102
rect 417306 580046 417374 580102
rect 417430 580046 417498 580102
rect 417554 580046 417622 580102
rect 417678 580046 435250 580102
rect 435306 580046 435374 580102
rect 435430 580046 435498 580102
rect 435554 580046 435622 580102
rect 435678 580046 453250 580102
rect 453306 580046 453374 580102
rect 453430 580046 453498 580102
rect 453554 580046 453622 580102
rect 453678 580046 471250 580102
rect 471306 580046 471374 580102
rect 471430 580046 471498 580102
rect 471554 580046 471622 580102
rect 471678 580046 489250 580102
rect 489306 580046 489374 580102
rect 489430 580046 489498 580102
rect 489554 580046 489622 580102
rect 489678 580046 507250 580102
rect 507306 580046 507374 580102
rect 507430 580046 507498 580102
rect 507554 580046 507622 580102
rect 507678 580046 525250 580102
rect 525306 580046 525374 580102
rect 525430 580046 525498 580102
rect 525554 580046 525622 580102
rect 525678 580046 543250 580102
rect 543306 580046 543374 580102
rect 543430 580046 543498 580102
rect 543554 580046 543622 580102
rect 543678 580046 561250 580102
rect 561306 580046 561374 580102
rect 561430 580046 561498 580102
rect 561554 580046 561622 580102
rect 561678 580046 579250 580102
rect 579306 580046 579374 580102
rect 579430 580046 579498 580102
rect 579554 580046 579622 580102
rect 579678 580046 596496 580102
rect 596552 580046 596620 580102
rect 596676 580046 596744 580102
rect 596800 580046 596868 580102
rect 596924 580046 597980 580102
rect -1916 579978 597980 580046
rect -1916 579922 -860 579978
rect -804 579922 -736 579978
rect -680 579922 -612 579978
rect -556 579922 -488 579978
rect -432 579922 3250 579978
rect 3306 579922 3374 579978
rect 3430 579922 3498 579978
rect 3554 579922 3622 579978
rect 3678 579922 21250 579978
rect 21306 579922 21374 579978
rect 21430 579922 21498 579978
rect 21554 579922 21622 579978
rect 21678 579922 39250 579978
rect 39306 579922 39374 579978
rect 39430 579922 39498 579978
rect 39554 579922 39622 579978
rect 39678 579922 57250 579978
rect 57306 579922 57374 579978
rect 57430 579922 57498 579978
rect 57554 579922 57622 579978
rect 57678 579922 75250 579978
rect 75306 579922 75374 579978
rect 75430 579922 75498 579978
rect 75554 579922 75622 579978
rect 75678 579922 93250 579978
rect 93306 579922 93374 579978
rect 93430 579922 93498 579978
rect 93554 579922 93622 579978
rect 93678 579922 111250 579978
rect 111306 579922 111374 579978
rect 111430 579922 111498 579978
rect 111554 579922 111622 579978
rect 111678 579922 129250 579978
rect 129306 579922 129374 579978
rect 129430 579922 129498 579978
rect 129554 579922 129622 579978
rect 129678 579922 147250 579978
rect 147306 579922 147374 579978
rect 147430 579922 147498 579978
rect 147554 579922 147622 579978
rect 147678 579922 165250 579978
rect 165306 579922 165374 579978
rect 165430 579922 165498 579978
rect 165554 579922 165622 579978
rect 165678 579922 183250 579978
rect 183306 579922 183374 579978
rect 183430 579922 183498 579978
rect 183554 579922 183622 579978
rect 183678 579922 201250 579978
rect 201306 579922 201374 579978
rect 201430 579922 201498 579978
rect 201554 579922 201622 579978
rect 201678 579922 219250 579978
rect 219306 579922 219374 579978
rect 219430 579922 219498 579978
rect 219554 579922 219622 579978
rect 219678 579922 237250 579978
rect 237306 579922 237374 579978
rect 237430 579922 237498 579978
rect 237554 579922 237622 579978
rect 237678 579922 255250 579978
rect 255306 579922 255374 579978
rect 255430 579922 255498 579978
rect 255554 579922 255622 579978
rect 255678 579922 273250 579978
rect 273306 579922 273374 579978
rect 273430 579922 273498 579978
rect 273554 579922 273622 579978
rect 273678 579922 291250 579978
rect 291306 579922 291374 579978
rect 291430 579922 291498 579978
rect 291554 579922 291622 579978
rect 291678 579922 309250 579978
rect 309306 579922 309374 579978
rect 309430 579922 309498 579978
rect 309554 579922 309622 579978
rect 309678 579922 327250 579978
rect 327306 579922 327374 579978
rect 327430 579922 327498 579978
rect 327554 579922 327622 579978
rect 327678 579922 345250 579978
rect 345306 579922 345374 579978
rect 345430 579922 345498 579978
rect 345554 579922 345622 579978
rect 345678 579922 363250 579978
rect 363306 579922 363374 579978
rect 363430 579922 363498 579978
rect 363554 579922 363622 579978
rect 363678 579922 381250 579978
rect 381306 579922 381374 579978
rect 381430 579922 381498 579978
rect 381554 579922 381622 579978
rect 381678 579922 399250 579978
rect 399306 579922 399374 579978
rect 399430 579922 399498 579978
rect 399554 579922 399622 579978
rect 399678 579922 417250 579978
rect 417306 579922 417374 579978
rect 417430 579922 417498 579978
rect 417554 579922 417622 579978
rect 417678 579922 435250 579978
rect 435306 579922 435374 579978
rect 435430 579922 435498 579978
rect 435554 579922 435622 579978
rect 435678 579922 453250 579978
rect 453306 579922 453374 579978
rect 453430 579922 453498 579978
rect 453554 579922 453622 579978
rect 453678 579922 471250 579978
rect 471306 579922 471374 579978
rect 471430 579922 471498 579978
rect 471554 579922 471622 579978
rect 471678 579922 489250 579978
rect 489306 579922 489374 579978
rect 489430 579922 489498 579978
rect 489554 579922 489622 579978
rect 489678 579922 507250 579978
rect 507306 579922 507374 579978
rect 507430 579922 507498 579978
rect 507554 579922 507622 579978
rect 507678 579922 525250 579978
rect 525306 579922 525374 579978
rect 525430 579922 525498 579978
rect 525554 579922 525622 579978
rect 525678 579922 543250 579978
rect 543306 579922 543374 579978
rect 543430 579922 543498 579978
rect 543554 579922 543622 579978
rect 543678 579922 561250 579978
rect 561306 579922 561374 579978
rect 561430 579922 561498 579978
rect 561554 579922 561622 579978
rect 561678 579922 579250 579978
rect 579306 579922 579374 579978
rect 579430 579922 579498 579978
rect 579554 579922 579622 579978
rect 579678 579922 596496 579978
rect 596552 579922 596620 579978
rect 596676 579922 596744 579978
rect 596800 579922 596868 579978
rect 596924 579922 597980 579978
rect -1916 579826 597980 579922
rect -1916 568350 597980 568446
rect -1916 568294 -1820 568350
rect -1764 568294 -1696 568350
rect -1640 568294 -1572 568350
rect -1516 568294 -1448 568350
rect -1392 568294 6970 568350
rect 7026 568294 7094 568350
rect 7150 568294 7218 568350
rect 7274 568294 7342 568350
rect 7398 568294 24970 568350
rect 25026 568294 25094 568350
rect 25150 568294 25218 568350
rect 25274 568294 25342 568350
rect 25398 568294 42970 568350
rect 43026 568294 43094 568350
rect 43150 568294 43218 568350
rect 43274 568294 43342 568350
rect 43398 568294 60970 568350
rect 61026 568294 61094 568350
rect 61150 568294 61218 568350
rect 61274 568294 61342 568350
rect 61398 568294 78970 568350
rect 79026 568294 79094 568350
rect 79150 568294 79218 568350
rect 79274 568294 79342 568350
rect 79398 568294 96970 568350
rect 97026 568294 97094 568350
rect 97150 568294 97218 568350
rect 97274 568294 97342 568350
rect 97398 568294 114970 568350
rect 115026 568294 115094 568350
rect 115150 568294 115218 568350
rect 115274 568294 115342 568350
rect 115398 568294 132970 568350
rect 133026 568294 133094 568350
rect 133150 568294 133218 568350
rect 133274 568294 133342 568350
rect 133398 568294 150970 568350
rect 151026 568294 151094 568350
rect 151150 568294 151218 568350
rect 151274 568294 151342 568350
rect 151398 568294 168970 568350
rect 169026 568294 169094 568350
rect 169150 568294 169218 568350
rect 169274 568294 169342 568350
rect 169398 568294 186970 568350
rect 187026 568294 187094 568350
rect 187150 568294 187218 568350
rect 187274 568294 187342 568350
rect 187398 568294 204970 568350
rect 205026 568294 205094 568350
rect 205150 568294 205218 568350
rect 205274 568294 205342 568350
rect 205398 568294 222970 568350
rect 223026 568294 223094 568350
rect 223150 568294 223218 568350
rect 223274 568294 223342 568350
rect 223398 568294 240970 568350
rect 241026 568294 241094 568350
rect 241150 568294 241218 568350
rect 241274 568294 241342 568350
rect 241398 568294 258970 568350
rect 259026 568294 259094 568350
rect 259150 568294 259218 568350
rect 259274 568294 259342 568350
rect 259398 568294 276970 568350
rect 277026 568294 277094 568350
rect 277150 568294 277218 568350
rect 277274 568294 277342 568350
rect 277398 568294 294970 568350
rect 295026 568294 295094 568350
rect 295150 568294 295218 568350
rect 295274 568294 295342 568350
rect 295398 568294 312970 568350
rect 313026 568294 313094 568350
rect 313150 568294 313218 568350
rect 313274 568294 313342 568350
rect 313398 568294 330970 568350
rect 331026 568294 331094 568350
rect 331150 568294 331218 568350
rect 331274 568294 331342 568350
rect 331398 568294 348970 568350
rect 349026 568294 349094 568350
rect 349150 568294 349218 568350
rect 349274 568294 349342 568350
rect 349398 568294 366970 568350
rect 367026 568294 367094 568350
rect 367150 568294 367218 568350
rect 367274 568294 367342 568350
rect 367398 568294 384970 568350
rect 385026 568294 385094 568350
rect 385150 568294 385218 568350
rect 385274 568294 385342 568350
rect 385398 568294 402970 568350
rect 403026 568294 403094 568350
rect 403150 568294 403218 568350
rect 403274 568294 403342 568350
rect 403398 568294 420970 568350
rect 421026 568294 421094 568350
rect 421150 568294 421218 568350
rect 421274 568294 421342 568350
rect 421398 568294 438970 568350
rect 439026 568294 439094 568350
rect 439150 568294 439218 568350
rect 439274 568294 439342 568350
rect 439398 568294 456970 568350
rect 457026 568294 457094 568350
rect 457150 568294 457218 568350
rect 457274 568294 457342 568350
rect 457398 568294 474970 568350
rect 475026 568294 475094 568350
rect 475150 568294 475218 568350
rect 475274 568294 475342 568350
rect 475398 568294 492970 568350
rect 493026 568294 493094 568350
rect 493150 568294 493218 568350
rect 493274 568294 493342 568350
rect 493398 568294 510970 568350
rect 511026 568294 511094 568350
rect 511150 568294 511218 568350
rect 511274 568294 511342 568350
rect 511398 568294 528970 568350
rect 529026 568294 529094 568350
rect 529150 568294 529218 568350
rect 529274 568294 529342 568350
rect 529398 568294 546970 568350
rect 547026 568294 547094 568350
rect 547150 568294 547218 568350
rect 547274 568294 547342 568350
rect 547398 568294 564970 568350
rect 565026 568294 565094 568350
rect 565150 568294 565218 568350
rect 565274 568294 565342 568350
rect 565398 568294 582970 568350
rect 583026 568294 583094 568350
rect 583150 568294 583218 568350
rect 583274 568294 583342 568350
rect 583398 568294 597456 568350
rect 597512 568294 597580 568350
rect 597636 568294 597704 568350
rect 597760 568294 597828 568350
rect 597884 568294 597980 568350
rect -1916 568226 597980 568294
rect -1916 568170 -1820 568226
rect -1764 568170 -1696 568226
rect -1640 568170 -1572 568226
rect -1516 568170 -1448 568226
rect -1392 568170 6970 568226
rect 7026 568170 7094 568226
rect 7150 568170 7218 568226
rect 7274 568170 7342 568226
rect 7398 568170 24970 568226
rect 25026 568170 25094 568226
rect 25150 568170 25218 568226
rect 25274 568170 25342 568226
rect 25398 568170 42970 568226
rect 43026 568170 43094 568226
rect 43150 568170 43218 568226
rect 43274 568170 43342 568226
rect 43398 568170 60970 568226
rect 61026 568170 61094 568226
rect 61150 568170 61218 568226
rect 61274 568170 61342 568226
rect 61398 568170 78970 568226
rect 79026 568170 79094 568226
rect 79150 568170 79218 568226
rect 79274 568170 79342 568226
rect 79398 568170 96970 568226
rect 97026 568170 97094 568226
rect 97150 568170 97218 568226
rect 97274 568170 97342 568226
rect 97398 568170 114970 568226
rect 115026 568170 115094 568226
rect 115150 568170 115218 568226
rect 115274 568170 115342 568226
rect 115398 568170 132970 568226
rect 133026 568170 133094 568226
rect 133150 568170 133218 568226
rect 133274 568170 133342 568226
rect 133398 568170 150970 568226
rect 151026 568170 151094 568226
rect 151150 568170 151218 568226
rect 151274 568170 151342 568226
rect 151398 568170 168970 568226
rect 169026 568170 169094 568226
rect 169150 568170 169218 568226
rect 169274 568170 169342 568226
rect 169398 568170 186970 568226
rect 187026 568170 187094 568226
rect 187150 568170 187218 568226
rect 187274 568170 187342 568226
rect 187398 568170 204970 568226
rect 205026 568170 205094 568226
rect 205150 568170 205218 568226
rect 205274 568170 205342 568226
rect 205398 568170 222970 568226
rect 223026 568170 223094 568226
rect 223150 568170 223218 568226
rect 223274 568170 223342 568226
rect 223398 568170 240970 568226
rect 241026 568170 241094 568226
rect 241150 568170 241218 568226
rect 241274 568170 241342 568226
rect 241398 568170 258970 568226
rect 259026 568170 259094 568226
rect 259150 568170 259218 568226
rect 259274 568170 259342 568226
rect 259398 568170 276970 568226
rect 277026 568170 277094 568226
rect 277150 568170 277218 568226
rect 277274 568170 277342 568226
rect 277398 568170 294970 568226
rect 295026 568170 295094 568226
rect 295150 568170 295218 568226
rect 295274 568170 295342 568226
rect 295398 568170 312970 568226
rect 313026 568170 313094 568226
rect 313150 568170 313218 568226
rect 313274 568170 313342 568226
rect 313398 568170 330970 568226
rect 331026 568170 331094 568226
rect 331150 568170 331218 568226
rect 331274 568170 331342 568226
rect 331398 568170 348970 568226
rect 349026 568170 349094 568226
rect 349150 568170 349218 568226
rect 349274 568170 349342 568226
rect 349398 568170 366970 568226
rect 367026 568170 367094 568226
rect 367150 568170 367218 568226
rect 367274 568170 367342 568226
rect 367398 568170 384970 568226
rect 385026 568170 385094 568226
rect 385150 568170 385218 568226
rect 385274 568170 385342 568226
rect 385398 568170 402970 568226
rect 403026 568170 403094 568226
rect 403150 568170 403218 568226
rect 403274 568170 403342 568226
rect 403398 568170 420970 568226
rect 421026 568170 421094 568226
rect 421150 568170 421218 568226
rect 421274 568170 421342 568226
rect 421398 568170 438970 568226
rect 439026 568170 439094 568226
rect 439150 568170 439218 568226
rect 439274 568170 439342 568226
rect 439398 568170 456970 568226
rect 457026 568170 457094 568226
rect 457150 568170 457218 568226
rect 457274 568170 457342 568226
rect 457398 568170 474970 568226
rect 475026 568170 475094 568226
rect 475150 568170 475218 568226
rect 475274 568170 475342 568226
rect 475398 568170 492970 568226
rect 493026 568170 493094 568226
rect 493150 568170 493218 568226
rect 493274 568170 493342 568226
rect 493398 568170 510970 568226
rect 511026 568170 511094 568226
rect 511150 568170 511218 568226
rect 511274 568170 511342 568226
rect 511398 568170 528970 568226
rect 529026 568170 529094 568226
rect 529150 568170 529218 568226
rect 529274 568170 529342 568226
rect 529398 568170 546970 568226
rect 547026 568170 547094 568226
rect 547150 568170 547218 568226
rect 547274 568170 547342 568226
rect 547398 568170 564970 568226
rect 565026 568170 565094 568226
rect 565150 568170 565218 568226
rect 565274 568170 565342 568226
rect 565398 568170 582970 568226
rect 583026 568170 583094 568226
rect 583150 568170 583218 568226
rect 583274 568170 583342 568226
rect 583398 568170 597456 568226
rect 597512 568170 597580 568226
rect 597636 568170 597704 568226
rect 597760 568170 597828 568226
rect 597884 568170 597980 568226
rect -1916 568102 597980 568170
rect -1916 568046 -1820 568102
rect -1764 568046 -1696 568102
rect -1640 568046 -1572 568102
rect -1516 568046 -1448 568102
rect -1392 568046 6970 568102
rect 7026 568046 7094 568102
rect 7150 568046 7218 568102
rect 7274 568046 7342 568102
rect 7398 568046 24970 568102
rect 25026 568046 25094 568102
rect 25150 568046 25218 568102
rect 25274 568046 25342 568102
rect 25398 568046 42970 568102
rect 43026 568046 43094 568102
rect 43150 568046 43218 568102
rect 43274 568046 43342 568102
rect 43398 568046 60970 568102
rect 61026 568046 61094 568102
rect 61150 568046 61218 568102
rect 61274 568046 61342 568102
rect 61398 568046 78970 568102
rect 79026 568046 79094 568102
rect 79150 568046 79218 568102
rect 79274 568046 79342 568102
rect 79398 568046 96970 568102
rect 97026 568046 97094 568102
rect 97150 568046 97218 568102
rect 97274 568046 97342 568102
rect 97398 568046 114970 568102
rect 115026 568046 115094 568102
rect 115150 568046 115218 568102
rect 115274 568046 115342 568102
rect 115398 568046 132970 568102
rect 133026 568046 133094 568102
rect 133150 568046 133218 568102
rect 133274 568046 133342 568102
rect 133398 568046 150970 568102
rect 151026 568046 151094 568102
rect 151150 568046 151218 568102
rect 151274 568046 151342 568102
rect 151398 568046 168970 568102
rect 169026 568046 169094 568102
rect 169150 568046 169218 568102
rect 169274 568046 169342 568102
rect 169398 568046 186970 568102
rect 187026 568046 187094 568102
rect 187150 568046 187218 568102
rect 187274 568046 187342 568102
rect 187398 568046 204970 568102
rect 205026 568046 205094 568102
rect 205150 568046 205218 568102
rect 205274 568046 205342 568102
rect 205398 568046 222970 568102
rect 223026 568046 223094 568102
rect 223150 568046 223218 568102
rect 223274 568046 223342 568102
rect 223398 568046 240970 568102
rect 241026 568046 241094 568102
rect 241150 568046 241218 568102
rect 241274 568046 241342 568102
rect 241398 568046 258970 568102
rect 259026 568046 259094 568102
rect 259150 568046 259218 568102
rect 259274 568046 259342 568102
rect 259398 568046 276970 568102
rect 277026 568046 277094 568102
rect 277150 568046 277218 568102
rect 277274 568046 277342 568102
rect 277398 568046 294970 568102
rect 295026 568046 295094 568102
rect 295150 568046 295218 568102
rect 295274 568046 295342 568102
rect 295398 568046 312970 568102
rect 313026 568046 313094 568102
rect 313150 568046 313218 568102
rect 313274 568046 313342 568102
rect 313398 568046 330970 568102
rect 331026 568046 331094 568102
rect 331150 568046 331218 568102
rect 331274 568046 331342 568102
rect 331398 568046 348970 568102
rect 349026 568046 349094 568102
rect 349150 568046 349218 568102
rect 349274 568046 349342 568102
rect 349398 568046 366970 568102
rect 367026 568046 367094 568102
rect 367150 568046 367218 568102
rect 367274 568046 367342 568102
rect 367398 568046 384970 568102
rect 385026 568046 385094 568102
rect 385150 568046 385218 568102
rect 385274 568046 385342 568102
rect 385398 568046 402970 568102
rect 403026 568046 403094 568102
rect 403150 568046 403218 568102
rect 403274 568046 403342 568102
rect 403398 568046 420970 568102
rect 421026 568046 421094 568102
rect 421150 568046 421218 568102
rect 421274 568046 421342 568102
rect 421398 568046 438970 568102
rect 439026 568046 439094 568102
rect 439150 568046 439218 568102
rect 439274 568046 439342 568102
rect 439398 568046 456970 568102
rect 457026 568046 457094 568102
rect 457150 568046 457218 568102
rect 457274 568046 457342 568102
rect 457398 568046 474970 568102
rect 475026 568046 475094 568102
rect 475150 568046 475218 568102
rect 475274 568046 475342 568102
rect 475398 568046 492970 568102
rect 493026 568046 493094 568102
rect 493150 568046 493218 568102
rect 493274 568046 493342 568102
rect 493398 568046 510970 568102
rect 511026 568046 511094 568102
rect 511150 568046 511218 568102
rect 511274 568046 511342 568102
rect 511398 568046 528970 568102
rect 529026 568046 529094 568102
rect 529150 568046 529218 568102
rect 529274 568046 529342 568102
rect 529398 568046 546970 568102
rect 547026 568046 547094 568102
rect 547150 568046 547218 568102
rect 547274 568046 547342 568102
rect 547398 568046 564970 568102
rect 565026 568046 565094 568102
rect 565150 568046 565218 568102
rect 565274 568046 565342 568102
rect 565398 568046 582970 568102
rect 583026 568046 583094 568102
rect 583150 568046 583218 568102
rect 583274 568046 583342 568102
rect 583398 568046 597456 568102
rect 597512 568046 597580 568102
rect 597636 568046 597704 568102
rect 597760 568046 597828 568102
rect 597884 568046 597980 568102
rect -1916 567978 597980 568046
rect -1916 567922 -1820 567978
rect -1764 567922 -1696 567978
rect -1640 567922 -1572 567978
rect -1516 567922 -1448 567978
rect -1392 567922 6970 567978
rect 7026 567922 7094 567978
rect 7150 567922 7218 567978
rect 7274 567922 7342 567978
rect 7398 567922 24970 567978
rect 25026 567922 25094 567978
rect 25150 567922 25218 567978
rect 25274 567922 25342 567978
rect 25398 567922 42970 567978
rect 43026 567922 43094 567978
rect 43150 567922 43218 567978
rect 43274 567922 43342 567978
rect 43398 567922 60970 567978
rect 61026 567922 61094 567978
rect 61150 567922 61218 567978
rect 61274 567922 61342 567978
rect 61398 567922 78970 567978
rect 79026 567922 79094 567978
rect 79150 567922 79218 567978
rect 79274 567922 79342 567978
rect 79398 567922 96970 567978
rect 97026 567922 97094 567978
rect 97150 567922 97218 567978
rect 97274 567922 97342 567978
rect 97398 567922 114970 567978
rect 115026 567922 115094 567978
rect 115150 567922 115218 567978
rect 115274 567922 115342 567978
rect 115398 567922 132970 567978
rect 133026 567922 133094 567978
rect 133150 567922 133218 567978
rect 133274 567922 133342 567978
rect 133398 567922 150970 567978
rect 151026 567922 151094 567978
rect 151150 567922 151218 567978
rect 151274 567922 151342 567978
rect 151398 567922 168970 567978
rect 169026 567922 169094 567978
rect 169150 567922 169218 567978
rect 169274 567922 169342 567978
rect 169398 567922 186970 567978
rect 187026 567922 187094 567978
rect 187150 567922 187218 567978
rect 187274 567922 187342 567978
rect 187398 567922 204970 567978
rect 205026 567922 205094 567978
rect 205150 567922 205218 567978
rect 205274 567922 205342 567978
rect 205398 567922 222970 567978
rect 223026 567922 223094 567978
rect 223150 567922 223218 567978
rect 223274 567922 223342 567978
rect 223398 567922 240970 567978
rect 241026 567922 241094 567978
rect 241150 567922 241218 567978
rect 241274 567922 241342 567978
rect 241398 567922 258970 567978
rect 259026 567922 259094 567978
rect 259150 567922 259218 567978
rect 259274 567922 259342 567978
rect 259398 567922 276970 567978
rect 277026 567922 277094 567978
rect 277150 567922 277218 567978
rect 277274 567922 277342 567978
rect 277398 567922 294970 567978
rect 295026 567922 295094 567978
rect 295150 567922 295218 567978
rect 295274 567922 295342 567978
rect 295398 567922 312970 567978
rect 313026 567922 313094 567978
rect 313150 567922 313218 567978
rect 313274 567922 313342 567978
rect 313398 567922 330970 567978
rect 331026 567922 331094 567978
rect 331150 567922 331218 567978
rect 331274 567922 331342 567978
rect 331398 567922 348970 567978
rect 349026 567922 349094 567978
rect 349150 567922 349218 567978
rect 349274 567922 349342 567978
rect 349398 567922 366970 567978
rect 367026 567922 367094 567978
rect 367150 567922 367218 567978
rect 367274 567922 367342 567978
rect 367398 567922 384970 567978
rect 385026 567922 385094 567978
rect 385150 567922 385218 567978
rect 385274 567922 385342 567978
rect 385398 567922 402970 567978
rect 403026 567922 403094 567978
rect 403150 567922 403218 567978
rect 403274 567922 403342 567978
rect 403398 567922 420970 567978
rect 421026 567922 421094 567978
rect 421150 567922 421218 567978
rect 421274 567922 421342 567978
rect 421398 567922 438970 567978
rect 439026 567922 439094 567978
rect 439150 567922 439218 567978
rect 439274 567922 439342 567978
rect 439398 567922 456970 567978
rect 457026 567922 457094 567978
rect 457150 567922 457218 567978
rect 457274 567922 457342 567978
rect 457398 567922 474970 567978
rect 475026 567922 475094 567978
rect 475150 567922 475218 567978
rect 475274 567922 475342 567978
rect 475398 567922 492970 567978
rect 493026 567922 493094 567978
rect 493150 567922 493218 567978
rect 493274 567922 493342 567978
rect 493398 567922 510970 567978
rect 511026 567922 511094 567978
rect 511150 567922 511218 567978
rect 511274 567922 511342 567978
rect 511398 567922 528970 567978
rect 529026 567922 529094 567978
rect 529150 567922 529218 567978
rect 529274 567922 529342 567978
rect 529398 567922 546970 567978
rect 547026 567922 547094 567978
rect 547150 567922 547218 567978
rect 547274 567922 547342 567978
rect 547398 567922 564970 567978
rect 565026 567922 565094 567978
rect 565150 567922 565218 567978
rect 565274 567922 565342 567978
rect 565398 567922 582970 567978
rect 583026 567922 583094 567978
rect 583150 567922 583218 567978
rect 583274 567922 583342 567978
rect 583398 567922 597456 567978
rect 597512 567922 597580 567978
rect 597636 567922 597704 567978
rect 597760 567922 597828 567978
rect 597884 567922 597980 567978
rect -1916 567826 597980 567922
rect -1916 562350 597980 562446
rect -1916 562294 -860 562350
rect -804 562294 -736 562350
rect -680 562294 -612 562350
rect -556 562294 -488 562350
rect -432 562294 3250 562350
rect 3306 562294 3374 562350
rect 3430 562294 3498 562350
rect 3554 562294 3622 562350
rect 3678 562294 21250 562350
rect 21306 562294 21374 562350
rect 21430 562294 21498 562350
rect 21554 562294 21622 562350
rect 21678 562294 39250 562350
rect 39306 562294 39374 562350
rect 39430 562294 39498 562350
rect 39554 562294 39622 562350
rect 39678 562294 57250 562350
rect 57306 562294 57374 562350
rect 57430 562294 57498 562350
rect 57554 562294 57622 562350
rect 57678 562294 75250 562350
rect 75306 562294 75374 562350
rect 75430 562294 75498 562350
rect 75554 562294 75622 562350
rect 75678 562294 93250 562350
rect 93306 562294 93374 562350
rect 93430 562294 93498 562350
rect 93554 562294 93622 562350
rect 93678 562294 111250 562350
rect 111306 562294 111374 562350
rect 111430 562294 111498 562350
rect 111554 562294 111622 562350
rect 111678 562294 129250 562350
rect 129306 562294 129374 562350
rect 129430 562294 129498 562350
rect 129554 562294 129622 562350
rect 129678 562294 147250 562350
rect 147306 562294 147374 562350
rect 147430 562294 147498 562350
rect 147554 562294 147622 562350
rect 147678 562294 165250 562350
rect 165306 562294 165374 562350
rect 165430 562294 165498 562350
rect 165554 562294 165622 562350
rect 165678 562294 183250 562350
rect 183306 562294 183374 562350
rect 183430 562294 183498 562350
rect 183554 562294 183622 562350
rect 183678 562294 201250 562350
rect 201306 562294 201374 562350
rect 201430 562294 201498 562350
rect 201554 562294 201622 562350
rect 201678 562294 219250 562350
rect 219306 562294 219374 562350
rect 219430 562294 219498 562350
rect 219554 562294 219622 562350
rect 219678 562294 237250 562350
rect 237306 562294 237374 562350
rect 237430 562294 237498 562350
rect 237554 562294 237622 562350
rect 237678 562294 255250 562350
rect 255306 562294 255374 562350
rect 255430 562294 255498 562350
rect 255554 562294 255622 562350
rect 255678 562294 273250 562350
rect 273306 562294 273374 562350
rect 273430 562294 273498 562350
rect 273554 562294 273622 562350
rect 273678 562294 291250 562350
rect 291306 562294 291374 562350
rect 291430 562294 291498 562350
rect 291554 562294 291622 562350
rect 291678 562294 309250 562350
rect 309306 562294 309374 562350
rect 309430 562294 309498 562350
rect 309554 562294 309622 562350
rect 309678 562294 327250 562350
rect 327306 562294 327374 562350
rect 327430 562294 327498 562350
rect 327554 562294 327622 562350
rect 327678 562294 345250 562350
rect 345306 562294 345374 562350
rect 345430 562294 345498 562350
rect 345554 562294 345622 562350
rect 345678 562294 363250 562350
rect 363306 562294 363374 562350
rect 363430 562294 363498 562350
rect 363554 562294 363622 562350
rect 363678 562294 381250 562350
rect 381306 562294 381374 562350
rect 381430 562294 381498 562350
rect 381554 562294 381622 562350
rect 381678 562294 399250 562350
rect 399306 562294 399374 562350
rect 399430 562294 399498 562350
rect 399554 562294 399622 562350
rect 399678 562294 417250 562350
rect 417306 562294 417374 562350
rect 417430 562294 417498 562350
rect 417554 562294 417622 562350
rect 417678 562294 435250 562350
rect 435306 562294 435374 562350
rect 435430 562294 435498 562350
rect 435554 562294 435622 562350
rect 435678 562294 453250 562350
rect 453306 562294 453374 562350
rect 453430 562294 453498 562350
rect 453554 562294 453622 562350
rect 453678 562294 471250 562350
rect 471306 562294 471374 562350
rect 471430 562294 471498 562350
rect 471554 562294 471622 562350
rect 471678 562294 489250 562350
rect 489306 562294 489374 562350
rect 489430 562294 489498 562350
rect 489554 562294 489622 562350
rect 489678 562294 507250 562350
rect 507306 562294 507374 562350
rect 507430 562294 507498 562350
rect 507554 562294 507622 562350
rect 507678 562294 525250 562350
rect 525306 562294 525374 562350
rect 525430 562294 525498 562350
rect 525554 562294 525622 562350
rect 525678 562294 543250 562350
rect 543306 562294 543374 562350
rect 543430 562294 543498 562350
rect 543554 562294 543622 562350
rect 543678 562294 561250 562350
rect 561306 562294 561374 562350
rect 561430 562294 561498 562350
rect 561554 562294 561622 562350
rect 561678 562294 579250 562350
rect 579306 562294 579374 562350
rect 579430 562294 579498 562350
rect 579554 562294 579622 562350
rect 579678 562294 596496 562350
rect 596552 562294 596620 562350
rect 596676 562294 596744 562350
rect 596800 562294 596868 562350
rect 596924 562294 597980 562350
rect -1916 562226 597980 562294
rect -1916 562170 -860 562226
rect -804 562170 -736 562226
rect -680 562170 -612 562226
rect -556 562170 -488 562226
rect -432 562170 3250 562226
rect 3306 562170 3374 562226
rect 3430 562170 3498 562226
rect 3554 562170 3622 562226
rect 3678 562170 21250 562226
rect 21306 562170 21374 562226
rect 21430 562170 21498 562226
rect 21554 562170 21622 562226
rect 21678 562170 39250 562226
rect 39306 562170 39374 562226
rect 39430 562170 39498 562226
rect 39554 562170 39622 562226
rect 39678 562170 57250 562226
rect 57306 562170 57374 562226
rect 57430 562170 57498 562226
rect 57554 562170 57622 562226
rect 57678 562170 75250 562226
rect 75306 562170 75374 562226
rect 75430 562170 75498 562226
rect 75554 562170 75622 562226
rect 75678 562170 93250 562226
rect 93306 562170 93374 562226
rect 93430 562170 93498 562226
rect 93554 562170 93622 562226
rect 93678 562170 111250 562226
rect 111306 562170 111374 562226
rect 111430 562170 111498 562226
rect 111554 562170 111622 562226
rect 111678 562170 129250 562226
rect 129306 562170 129374 562226
rect 129430 562170 129498 562226
rect 129554 562170 129622 562226
rect 129678 562170 147250 562226
rect 147306 562170 147374 562226
rect 147430 562170 147498 562226
rect 147554 562170 147622 562226
rect 147678 562170 165250 562226
rect 165306 562170 165374 562226
rect 165430 562170 165498 562226
rect 165554 562170 165622 562226
rect 165678 562170 183250 562226
rect 183306 562170 183374 562226
rect 183430 562170 183498 562226
rect 183554 562170 183622 562226
rect 183678 562170 201250 562226
rect 201306 562170 201374 562226
rect 201430 562170 201498 562226
rect 201554 562170 201622 562226
rect 201678 562170 219250 562226
rect 219306 562170 219374 562226
rect 219430 562170 219498 562226
rect 219554 562170 219622 562226
rect 219678 562170 237250 562226
rect 237306 562170 237374 562226
rect 237430 562170 237498 562226
rect 237554 562170 237622 562226
rect 237678 562170 255250 562226
rect 255306 562170 255374 562226
rect 255430 562170 255498 562226
rect 255554 562170 255622 562226
rect 255678 562170 273250 562226
rect 273306 562170 273374 562226
rect 273430 562170 273498 562226
rect 273554 562170 273622 562226
rect 273678 562170 291250 562226
rect 291306 562170 291374 562226
rect 291430 562170 291498 562226
rect 291554 562170 291622 562226
rect 291678 562170 309250 562226
rect 309306 562170 309374 562226
rect 309430 562170 309498 562226
rect 309554 562170 309622 562226
rect 309678 562170 327250 562226
rect 327306 562170 327374 562226
rect 327430 562170 327498 562226
rect 327554 562170 327622 562226
rect 327678 562170 345250 562226
rect 345306 562170 345374 562226
rect 345430 562170 345498 562226
rect 345554 562170 345622 562226
rect 345678 562170 363250 562226
rect 363306 562170 363374 562226
rect 363430 562170 363498 562226
rect 363554 562170 363622 562226
rect 363678 562170 381250 562226
rect 381306 562170 381374 562226
rect 381430 562170 381498 562226
rect 381554 562170 381622 562226
rect 381678 562170 399250 562226
rect 399306 562170 399374 562226
rect 399430 562170 399498 562226
rect 399554 562170 399622 562226
rect 399678 562170 417250 562226
rect 417306 562170 417374 562226
rect 417430 562170 417498 562226
rect 417554 562170 417622 562226
rect 417678 562170 435250 562226
rect 435306 562170 435374 562226
rect 435430 562170 435498 562226
rect 435554 562170 435622 562226
rect 435678 562170 453250 562226
rect 453306 562170 453374 562226
rect 453430 562170 453498 562226
rect 453554 562170 453622 562226
rect 453678 562170 471250 562226
rect 471306 562170 471374 562226
rect 471430 562170 471498 562226
rect 471554 562170 471622 562226
rect 471678 562170 489250 562226
rect 489306 562170 489374 562226
rect 489430 562170 489498 562226
rect 489554 562170 489622 562226
rect 489678 562170 507250 562226
rect 507306 562170 507374 562226
rect 507430 562170 507498 562226
rect 507554 562170 507622 562226
rect 507678 562170 525250 562226
rect 525306 562170 525374 562226
rect 525430 562170 525498 562226
rect 525554 562170 525622 562226
rect 525678 562170 543250 562226
rect 543306 562170 543374 562226
rect 543430 562170 543498 562226
rect 543554 562170 543622 562226
rect 543678 562170 561250 562226
rect 561306 562170 561374 562226
rect 561430 562170 561498 562226
rect 561554 562170 561622 562226
rect 561678 562170 579250 562226
rect 579306 562170 579374 562226
rect 579430 562170 579498 562226
rect 579554 562170 579622 562226
rect 579678 562170 596496 562226
rect 596552 562170 596620 562226
rect 596676 562170 596744 562226
rect 596800 562170 596868 562226
rect 596924 562170 597980 562226
rect -1916 562102 597980 562170
rect -1916 562046 -860 562102
rect -804 562046 -736 562102
rect -680 562046 -612 562102
rect -556 562046 -488 562102
rect -432 562046 3250 562102
rect 3306 562046 3374 562102
rect 3430 562046 3498 562102
rect 3554 562046 3622 562102
rect 3678 562046 21250 562102
rect 21306 562046 21374 562102
rect 21430 562046 21498 562102
rect 21554 562046 21622 562102
rect 21678 562046 39250 562102
rect 39306 562046 39374 562102
rect 39430 562046 39498 562102
rect 39554 562046 39622 562102
rect 39678 562046 57250 562102
rect 57306 562046 57374 562102
rect 57430 562046 57498 562102
rect 57554 562046 57622 562102
rect 57678 562046 75250 562102
rect 75306 562046 75374 562102
rect 75430 562046 75498 562102
rect 75554 562046 75622 562102
rect 75678 562046 93250 562102
rect 93306 562046 93374 562102
rect 93430 562046 93498 562102
rect 93554 562046 93622 562102
rect 93678 562046 111250 562102
rect 111306 562046 111374 562102
rect 111430 562046 111498 562102
rect 111554 562046 111622 562102
rect 111678 562046 129250 562102
rect 129306 562046 129374 562102
rect 129430 562046 129498 562102
rect 129554 562046 129622 562102
rect 129678 562046 147250 562102
rect 147306 562046 147374 562102
rect 147430 562046 147498 562102
rect 147554 562046 147622 562102
rect 147678 562046 165250 562102
rect 165306 562046 165374 562102
rect 165430 562046 165498 562102
rect 165554 562046 165622 562102
rect 165678 562046 183250 562102
rect 183306 562046 183374 562102
rect 183430 562046 183498 562102
rect 183554 562046 183622 562102
rect 183678 562046 201250 562102
rect 201306 562046 201374 562102
rect 201430 562046 201498 562102
rect 201554 562046 201622 562102
rect 201678 562046 219250 562102
rect 219306 562046 219374 562102
rect 219430 562046 219498 562102
rect 219554 562046 219622 562102
rect 219678 562046 237250 562102
rect 237306 562046 237374 562102
rect 237430 562046 237498 562102
rect 237554 562046 237622 562102
rect 237678 562046 255250 562102
rect 255306 562046 255374 562102
rect 255430 562046 255498 562102
rect 255554 562046 255622 562102
rect 255678 562046 273250 562102
rect 273306 562046 273374 562102
rect 273430 562046 273498 562102
rect 273554 562046 273622 562102
rect 273678 562046 291250 562102
rect 291306 562046 291374 562102
rect 291430 562046 291498 562102
rect 291554 562046 291622 562102
rect 291678 562046 309250 562102
rect 309306 562046 309374 562102
rect 309430 562046 309498 562102
rect 309554 562046 309622 562102
rect 309678 562046 327250 562102
rect 327306 562046 327374 562102
rect 327430 562046 327498 562102
rect 327554 562046 327622 562102
rect 327678 562046 345250 562102
rect 345306 562046 345374 562102
rect 345430 562046 345498 562102
rect 345554 562046 345622 562102
rect 345678 562046 363250 562102
rect 363306 562046 363374 562102
rect 363430 562046 363498 562102
rect 363554 562046 363622 562102
rect 363678 562046 381250 562102
rect 381306 562046 381374 562102
rect 381430 562046 381498 562102
rect 381554 562046 381622 562102
rect 381678 562046 399250 562102
rect 399306 562046 399374 562102
rect 399430 562046 399498 562102
rect 399554 562046 399622 562102
rect 399678 562046 417250 562102
rect 417306 562046 417374 562102
rect 417430 562046 417498 562102
rect 417554 562046 417622 562102
rect 417678 562046 435250 562102
rect 435306 562046 435374 562102
rect 435430 562046 435498 562102
rect 435554 562046 435622 562102
rect 435678 562046 453250 562102
rect 453306 562046 453374 562102
rect 453430 562046 453498 562102
rect 453554 562046 453622 562102
rect 453678 562046 471250 562102
rect 471306 562046 471374 562102
rect 471430 562046 471498 562102
rect 471554 562046 471622 562102
rect 471678 562046 489250 562102
rect 489306 562046 489374 562102
rect 489430 562046 489498 562102
rect 489554 562046 489622 562102
rect 489678 562046 507250 562102
rect 507306 562046 507374 562102
rect 507430 562046 507498 562102
rect 507554 562046 507622 562102
rect 507678 562046 525250 562102
rect 525306 562046 525374 562102
rect 525430 562046 525498 562102
rect 525554 562046 525622 562102
rect 525678 562046 543250 562102
rect 543306 562046 543374 562102
rect 543430 562046 543498 562102
rect 543554 562046 543622 562102
rect 543678 562046 561250 562102
rect 561306 562046 561374 562102
rect 561430 562046 561498 562102
rect 561554 562046 561622 562102
rect 561678 562046 579250 562102
rect 579306 562046 579374 562102
rect 579430 562046 579498 562102
rect 579554 562046 579622 562102
rect 579678 562046 596496 562102
rect 596552 562046 596620 562102
rect 596676 562046 596744 562102
rect 596800 562046 596868 562102
rect 596924 562046 597980 562102
rect -1916 561978 597980 562046
rect -1916 561922 -860 561978
rect -804 561922 -736 561978
rect -680 561922 -612 561978
rect -556 561922 -488 561978
rect -432 561922 3250 561978
rect 3306 561922 3374 561978
rect 3430 561922 3498 561978
rect 3554 561922 3622 561978
rect 3678 561922 21250 561978
rect 21306 561922 21374 561978
rect 21430 561922 21498 561978
rect 21554 561922 21622 561978
rect 21678 561922 39250 561978
rect 39306 561922 39374 561978
rect 39430 561922 39498 561978
rect 39554 561922 39622 561978
rect 39678 561922 57250 561978
rect 57306 561922 57374 561978
rect 57430 561922 57498 561978
rect 57554 561922 57622 561978
rect 57678 561922 75250 561978
rect 75306 561922 75374 561978
rect 75430 561922 75498 561978
rect 75554 561922 75622 561978
rect 75678 561922 93250 561978
rect 93306 561922 93374 561978
rect 93430 561922 93498 561978
rect 93554 561922 93622 561978
rect 93678 561922 111250 561978
rect 111306 561922 111374 561978
rect 111430 561922 111498 561978
rect 111554 561922 111622 561978
rect 111678 561922 129250 561978
rect 129306 561922 129374 561978
rect 129430 561922 129498 561978
rect 129554 561922 129622 561978
rect 129678 561922 147250 561978
rect 147306 561922 147374 561978
rect 147430 561922 147498 561978
rect 147554 561922 147622 561978
rect 147678 561922 165250 561978
rect 165306 561922 165374 561978
rect 165430 561922 165498 561978
rect 165554 561922 165622 561978
rect 165678 561922 183250 561978
rect 183306 561922 183374 561978
rect 183430 561922 183498 561978
rect 183554 561922 183622 561978
rect 183678 561922 201250 561978
rect 201306 561922 201374 561978
rect 201430 561922 201498 561978
rect 201554 561922 201622 561978
rect 201678 561922 219250 561978
rect 219306 561922 219374 561978
rect 219430 561922 219498 561978
rect 219554 561922 219622 561978
rect 219678 561922 237250 561978
rect 237306 561922 237374 561978
rect 237430 561922 237498 561978
rect 237554 561922 237622 561978
rect 237678 561922 255250 561978
rect 255306 561922 255374 561978
rect 255430 561922 255498 561978
rect 255554 561922 255622 561978
rect 255678 561922 273250 561978
rect 273306 561922 273374 561978
rect 273430 561922 273498 561978
rect 273554 561922 273622 561978
rect 273678 561922 291250 561978
rect 291306 561922 291374 561978
rect 291430 561922 291498 561978
rect 291554 561922 291622 561978
rect 291678 561922 309250 561978
rect 309306 561922 309374 561978
rect 309430 561922 309498 561978
rect 309554 561922 309622 561978
rect 309678 561922 327250 561978
rect 327306 561922 327374 561978
rect 327430 561922 327498 561978
rect 327554 561922 327622 561978
rect 327678 561922 345250 561978
rect 345306 561922 345374 561978
rect 345430 561922 345498 561978
rect 345554 561922 345622 561978
rect 345678 561922 363250 561978
rect 363306 561922 363374 561978
rect 363430 561922 363498 561978
rect 363554 561922 363622 561978
rect 363678 561922 381250 561978
rect 381306 561922 381374 561978
rect 381430 561922 381498 561978
rect 381554 561922 381622 561978
rect 381678 561922 399250 561978
rect 399306 561922 399374 561978
rect 399430 561922 399498 561978
rect 399554 561922 399622 561978
rect 399678 561922 417250 561978
rect 417306 561922 417374 561978
rect 417430 561922 417498 561978
rect 417554 561922 417622 561978
rect 417678 561922 435250 561978
rect 435306 561922 435374 561978
rect 435430 561922 435498 561978
rect 435554 561922 435622 561978
rect 435678 561922 453250 561978
rect 453306 561922 453374 561978
rect 453430 561922 453498 561978
rect 453554 561922 453622 561978
rect 453678 561922 471250 561978
rect 471306 561922 471374 561978
rect 471430 561922 471498 561978
rect 471554 561922 471622 561978
rect 471678 561922 489250 561978
rect 489306 561922 489374 561978
rect 489430 561922 489498 561978
rect 489554 561922 489622 561978
rect 489678 561922 507250 561978
rect 507306 561922 507374 561978
rect 507430 561922 507498 561978
rect 507554 561922 507622 561978
rect 507678 561922 525250 561978
rect 525306 561922 525374 561978
rect 525430 561922 525498 561978
rect 525554 561922 525622 561978
rect 525678 561922 543250 561978
rect 543306 561922 543374 561978
rect 543430 561922 543498 561978
rect 543554 561922 543622 561978
rect 543678 561922 561250 561978
rect 561306 561922 561374 561978
rect 561430 561922 561498 561978
rect 561554 561922 561622 561978
rect 561678 561922 579250 561978
rect 579306 561922 579374 561978
rect 579430 561922 579498 561978
rect 579554 561922 579622 561978
rect 579678 561922 596496 561978
rect 596552 561922 596620 561978
rect 596676 561922 596744 561978
rect 596800 561922 596868 561978
rect 596924 561922 597980 561978
rect -1916 561826 597980 561922
rect -1916 550350 597980 550446
rect -1916 550294 -1820 550350
rect -1764 550294 -1696 550350
rect -1640 550294 -1572 550350
rect -1516 550294 -1448 550350
rect -1392 550294 6970 550350
rect 7026 550294 7094 550350
rect 7150 550294 7218 550350
rect 7274 550294 7342 550350
rect 7398 550294 24970 550350
rect 25026 550294 25094 550350
rect 25150 550294 25218 550350
rect 25274 550294 25342 550350
rect 25398 550294 42970 550350
rect 43026 550294 43094 550350
rect 43150 550294 43218 550350
rect 43274 550294 43342 550350
rect 43398 550294 60970 550350
rect 61026 550294 61094 550350
rect 61150 550294 61218 550350
rect 61274 550294 61342 550350
rect 61398 550294 78970 550350
rect 79026 550294 79094 550350
rect 79150 550294 79218 550350
rect 79274 550294 79342 550350
rect 79398 550294 96970 550350
rect 97026 550294 97094 550350
rect 97150 550294 97218 550350
rect 97274 550294 97342 550350
rect 97398 550294 114970 550350
rect 115026 550294 115094 550350
rect 115150 550294 115218 550350
rect 115274 550294 115342 550350
rect 115398 550294 132970 550350
rect 133026 550294 133094 550350
rect 133150 550294 133218 550350
rect 133274 550294 133342 550350
rect 133398 550294 150970 550350
rect 151026 550294 151094 550350
rect 151150 550294 151218 550350
rect 151274 550294 151342 550350
rect 151398 550294 168970 550350
rect 169026 550294 169094 550350
rect 169150 550294 169218 550350
rect 169274 550294 169342 550350
rect 169398 550294 186970 550350
rect 187026 550294 187094 550350
rect 187150 550294 187218 550350
rect 187274 550294 187342 550350
rect 187398 550294 204970 550350
rect 205026 550294 205094 550350
rect 205150 550294 205218 550350
rect 205274 550294 205342 550350
rect 205398 550294 222970 550350
rect 223026 550294 223094 550350
rect 223150 550294 223218 550350
rect 223274 550294 223342 550350
rect 223398 550294 240970 550350
rect 241026 550294 241094 550350
rect 241150 550294 241218 550350
rect 241274 550294 241342 550350
rect 241398 550294 258970 550350
rect 259026 550294 259094 550350
rect 259150 550294 259218 550350
rect 259274 550294 259342 550350
rect 259398 550294 276970 550350
rect 277026 550294 277094 550350
rect 277150 550294 277218 550350
rect 277274 550294 277342 550350
rect 277398 550294 294970 550350
rect 295026 550294 295094 550350
rect 295150 550294 295218 550350
rect 295274 550294 295342 550350
rect 295398 550294 312970 550350
rect 313026 550294 313094 550350
rect 313150 550294 313218 550350
rect 313274 550294 313342 550350
rect 313398 550294 330970 550350
rect 331026 550294 331094 550350
rect 331150 550294 331218 550350
rect 331274 550294 331342 550350
rect 331398 550294 348970 550350
rect 349026 550294 349094 550350
rect 349150 550294 349218 550350
rect 349274 550294 349342 550350
rect 349398 550294 366970 550350
rect 367026 550294 367094 550350
rect 367150 550294 367218 550350
rect 367274 550294 367342 550350
rect 367398 550294 384970 550350
rect 385026 550294 385094 550350
rect 385150 550294 385218 550350
rect 385274 550294 385342 550350
rect 385398 550294 402970 550350
rect 403026 550294 403094 550350
rect 403150 550294 403218 550350
rect 403274 550294 403342 550350
rect 403398 550294 420970 550350
rect 421026 550294 421094 550350
rect 421150 550294 421218 550350
rect 421274 550294 421342 550350
rect 421398 550294 438970 550350
rect 439026 550294 439094 550350
rect 439150 550294 439218 550350
rect 439274 550294 439342 550350
rect 439398 550294 456970 550350
rect 457026 550294 457094 550350
rect 457150 550294 457218 550350
rect 457274 550294 457342 550350
rect 457398 550294 474970 550350
rect 475026 550294 475094 550350
rect 475150 550294 475218 550350
rect 475274 550294 475342 550350
rect 475398 550294 492970 550350
rect 493026 550294 493094 550350
rect 493150 550294 493218 550350
rect 493274 550294 493342 550350
rect 493398 550294 510970 550350
rect 511026 550294 511094 550350
rect 511150 550294 511218 550350
rect 511274 550294 511342 550350
rect 511398 550294 528970 550350
rect 529026 550294 529094 550350
rect 529150 550294 529218 550350
rect 529274 550294 529342 550350
rect 529398 550294 546970 550350
rect 547026 550294 547094 550350
rect 547150 550294 547218 550350
rect 547274 550294 547342 550350
rect 547398 550294 564970 550350
rect 565026 550294 565094 550350
rect 565150 550294 565218 550350
rect 565274 550294 565342 550350
rect 565398 550294 582970 550350
rect 583026 550294 583094 550350
rect 583150 550294 583218 550350
rect 583274 550294 583342 550350
rect 583398 550294 597456 550350
rect 597512 550294 597580 550350
rect 597636 550294 597704 550350
rect 597760 550294 597828 550350
rect 597884 550294 597980 550350
rect -1916 550226 597980 550294
rect -1916 550170 -1820 550226
rect -1764 550170 -1696 550226
rect -1640 550170 -1572 550226
rect -1516 550170 -1448 550226
rect -1392 550170 6970 550226
rect 7026 550170 7094 550226
rect 7150 550170 7218 550226
rect 7274 550170 7342 550226
rect 7398 550170 24970 550226
rect 25026 550170 25094 550226
rect 25150 550170 25218 550226
rect 25274 550170 25342 550226
rect 25398 550170 42970 550226
rect 43026 550170 43094 550226
rect 43150 550170 43218 550226
rect 43274 550170 43342 550226
rect 43398 550170 60970 550226
rect 61026 550170 61094 550226
rect 61150 550170 61218 550226
rect 61274 550170 61342 550226
rect 61398 550170 78970 550226
rect 79026 550170 79094 550226
rect 79150 550170 79218 550226
rect 79274 550170 79342 550226
rect 79398 550170 96970 550226
rect 97026 550170 97094 550226
rect 97150 550170 97218 550226
rect 97274 550170 97342 550226
rect 97398 550170 114970 550226
rect 115026 550170 115094 550226
rect 115150 550170 115218 550226
rect 115274 550170 115342 550226
rect 115398 550170 132970 550226
rect 133026 550170 133094 550226
rect 133150 550170 133218 550226
rect 133274 550170 133342 550226
rect 133398 550170 150970 550226
rect 151026 550170 151094 550226
rect 151150 550170 151218 550226
rect 151274 550170 151342 550226
rect 151398 550170 168970 550226
rect 169026 550170 169094 550226
rect 169150 550170 169218 550226
rect 169274 550170 169342 550226
rect 169398 550170 186970 550226
rect 187026 550170 187094 550226
rect 187150 550170 187218 550226
rect 187274 550170 187342 550226
rect 187398 550170 204970 550226
rect 205026 550170 205094 550226
rect 205150 550170 205218 550226
rect 205274 550170 205342 550226
rect 205398 550170 222970 550226
rect 223026 550170 223094 550226
rect 223150 550170 223218 550226
rect 223274 550170 223342 550226
rect 223398 550170 240970 550226
rect 241026 550170 241094 550226
rect 241150 550170 241218 550226
rect 241274 550170 241342 550226
rect 241398 550170 258970 550226
rect 259026 550170 259094 550226
rect 259150 550170 259218 550226
rect 259274 550170 259342 550226
rect 259398 550170 276970 550226
rect 277026 550170 277094 550226
rect 277150 550170 277218 550226
rect 277274 550170 277342 550226
rect 277398 550170 294970 550226
rect 295026 550170 295094 550226
rect 295150 550170 295218 550226
rect 295274 550170 295342 550226
rect 295398 550170 312970 550226
rect 313026 550170 313094 550226
rect 313150 550170 313218 550226
rect 313274 550170 313342 550226
rect 313398 550170 330970 550226
rect 331026 550170 331094 550226
rect 331150 550170 331218 550226
rect 331274 550170 331342 550226
rect 331398 550170 348970 550226
rect 349026 550170 349094 550226
rect 349150 550170 349218 550226
rect 349274 550170 349342 550226
rect 349398 550170 366970 550226
rect 367026 550170 367094 550226
rect 367150 550170 367218 550226
rect 367274 550170 367342 550226
rect 367398 550170 384970 550226
rect 385026 550170 385094 550226
rect 385150 550170 385218 550226
rect 385274 550170 385342 550226
rect 385398 550170 402970 550226
rect 403026 550170 403094 550226
rect 403150 550170 403218 550226
rect 403274 550170 403342 550226
rect 403398 550170 420970 550226
rect 421026 550170 421094 550226
rect 421150 550170 421218 550226
rect 421274 550170 421342 550226
rect 421398 550170 438970 550226
rect 439026 550170 439094 550226
rect 439150 550170 439218 550226
rect 439274 550170 439342 550226
rect 439398 550170 456970 550226
rect 457026 550170 457094 550226
rect 457150 550170 457218 550226
rect 457274 550170 457342 550226
rect 457398 550170 474970 550226
rect 475026 550170 475094 550226
rect 475150 550170 475218 550226
rect 475274 550170 475342 550226
rect 475398 550170 492970 550226
rect 493026 550170 493094 550226
rect 493150 550170 493218 550226
rect 493274 550170 493342 550226
rect 493398 550170 510970 550226
rect 511026 550170 511094 550226
rect 511150 550170 511218 550226
rect 511274 550170 511342 550226
rect 511398 550170 528970 550226
rect 529026 550170 529094 550226
rect 529150 550170 529218 550226
rect 529274 550170 529342 550226
rect 529398 550170 546970 550226
rect 547026 550170 547094 550226
rect 547150 550170 547218 550226
rect 547274 550170 547342 550226
rect 547398 550170 564970 550226
rect 565026 550170 565094 550226
rect 565150 550170 565218 550226
rect 565274 550170 565342 550226
rect 565398 550170 582970 550226
rect 583026 550170 583094 550226
rect 583150 550170 583218 550226
rect 583274 550170 583342 550226
rect 583398 550170 597456 550226
rect 597512 550170 597580 550226
rect 597636 550170 597704 550226
rect 597760 550170 597828 550226
rect 597884 550170 597980 550226
rect -1916 550102 597980 550170
rect -1916 550046 -1820 550102
rect -1764 550046 -1696 550102
rect -1640 550046 -1572 550102
rect -1516 550046 -1448 550102
rect -1392 550046 6970 550102
rect 7026 550046 7094 550102
rect 7150 550046 7218 550102
rect 7274 550046 7342 550102
rect 7398 550046 24970 550102
rect 25026 550046 25094 550102
rect 25150 550046 25218 550102
rect 25274 550046 25342 550102
rect 25398 550046 42970 550102
rect 43026 550046 43094 550102
rect 43150 550046 43218 550102
rect 43274 550046 43342 550102
rect 43398 550046 60970 550102
rect 61026 550046 61094 550102
rect 61150 550046 61218 550102
rect 61274 550046 61342 550102
rect 61398 550046 78970 550102
rect 79026 550046 79094 550102
rect 79150 550046 79218 550102
rect 79274 550046 79342 550102
rect 79398 550046 96970 550102
rect 97026 550046 97094 550102
rect 97150 550046 97218 550102
rect 97274 550046 97342 550102
rect 97398 550046 114970 550102
rect 115026 550046 115094 550102
rect 115150 550046 115218 550102
rect 115274 550046 115342 550102
rect 115398 550046 132970 550102
rect 133026 550046 133094 550102
rect 133150 550046 133218 550102
rect 133274 550046 133342 550102
rect 133398 550046 150970 550102
rect 151026 550046 151094 550102
rect 151150 550046 151218 550102
rect 151274 550046 151342 550102
rect 151398 550046 168970 550102
rect 169026 550046 169094 550102
rect 169150 550046 169218 550102
rect 169274 550046 169342 550102
rect 169398 550046 186970 550102
rect 187026 550046 187094 550102
rect 187150 550046 187218 550102
rect 187274 550046 187342 550102
rect 187398 550046 204970 550102
rect 205026 550046 205094 550102
rect 205150 550046 205218 550102
rect 205274 550046 205342 550102
rect 205398 550046 222970 550102
rect 223026 550046 223094 550102
rect 223150 550046 223218 550102
rect 223274 550046 223342 550102
rect 223398 550046 240970 550102
rect 241026 550046 241094 550102
rect 241150 550046 241218 550102
rect 241274 550046 241342 550102
rect 241398 550046 258970 550102
rect 259026 550046 259094 550102
rect 259150 550046 259218 550102
rect 259274 550046 259342 550102
rect 259398 550046 276970 550102
rect 277026 550046 277094 550102
rect 277150 550046 277218 550102
rect 277274 550046 277342 550102
rect 277398 550046 294970 550102
rect 295026 550046 295094 550102
rect 295150 550046 295218 550102
rect 295274 550046 295342 550102
rect 295398 550046 312970 550102
rect 313026 550046 313094 550102
rect 313150 550046 313218 550102
rect 313274 550046 313342 550102
rect 313398 550046 330970 550102
rect 331026 550046 331094 550102
rect 331150 550046 331218 550102
rect 331274 550046 331342 550102
rect 331398 550046 348970 550102
rect 349026 550046 349094 550102
rect 349150 550046 349218 550102
rect 349274 550046 349342 550102
rect 349398 550046 366970 550102
rect 367026 550046 367094 550102
rect 367150 550046 367218 550102
rect 367274 550046 367342 550102
rect 367398 550046 384970 550102
rect 385026 550046 385094 550102
rect 385150 550046 385218 550102
rect 385274 550046 385342 550102
rect 385398 550046 402970 550102
rect 403026 550046 403094 550102
rect 403150 550046 403218 550102
rect 403274 550046 403342 550102
rect 403398 550046 420970 550102
rect 421026 550046 421094 550102
rect 421150 550046 421218 550102
rect 421274 550046 421342 550102
rect 421398 550046 438970 550102
rect 439026 550046 439094 550102
rect 439150 550046 439218 550102
rect 439274 550046 439342 550102
rect 439398 550046 456970 550102
rect 457026 550046 457094 550102
rect 457150 550046 457218 550102
rect 457274 550046 457342 550102
rect 457398 550046 474970 550102
rect 475026 550046 475094 550102
rect 475150 550046 475218 550102
rect 475274 550046 475342 550102
rect 475398 550046 492970 550102
rect 493026 550046 493094 550102
rect 493150 550046 493218 550102
rect 493274 550046 493342 550102
rect 493398 550046 510970 550102
rect 511026 550046 511094 550102
rect 511150 550046 511218 550102
rect 511274 550046 511342 550102
rect 511398 550046 528970 550102
rect 529026 550046 529094 550102
rect 529150 550046 529218 550102
rect 529274 550046 529342 550102
rect 529398 550046 546970 550102
rect 547026 550046 547094 550102
rect 547150 550046 547218 550102
rect 547274 550046 547342 550102
rect 547398 550046 564970 550102
rect 565026 550046 565094 550102
rect 565150 550046 565218 550102
rect 565274 550046 565342 550102
rect 565398 550046 582970 550102
rect 583026 550046 583094 550102
rect 583150 550046 583218 550102
rect 583274 550046 583342 550102
rect 583398 550046 597456 550102
rect 597512 550046 597580 550102
rect 597636 550046 597704 550102
rect 597760 550046 597828 550102
rect 597884 550046 597980 550102
rect -1916 549978 597980 550046
rect -1916 549922 -1820 549978
rect -1764 549922 -1696 549978
rect -1640 549922 -1572 549978
rect -1516 549922 -1448 549978
rect -1392 549922 6970 549978
rect 7026 549922 7094 549978
rect 7150 549922 7218 549978
rect 7274 549922 7342 549978
rect 7398 549922 24970 549978
rect 25026 549922 25094 549978
rect 25150 549922 25218 549978
rect 25274 549922 25342 549978
rect 25398 549922 42970 549978
rect 43026 549922 43094 549978
rect 43150 549922 43218 549978
rect 43274 549922 43342 549978
rect 43398 549922 60970 549978
rect 61026 549922 61094 549978
rect 61150 549922 61218 549978
rect 61274 549922 61342 549978
rect 61398 549922 78970 549978
rect 79026 549922 79094 549978
rect 79150 549922 79218 549978
rect 79274 549922 79342 549978
rect 79398 549922 96970 549978
rect 97026 549922 97094 549978
rect 97150 549922 97218 549978
rect 97274 549922 97342 549978
rect 97398 549922 114970 549978
rect 115026 549922 115094 549978
rect 115150 549922 115218 549978
rect 115274 549922 115342 549978
rect 115398 549922 132970 549978
rect 133026 549922 133094 549978
rect 133150 549922 133218 549978
rect 133274 549922 133342 549978
rect 133398 549922 150970 549978
rect 151026 549922 151094 549978
rect 151150 549922 151218 549978
rect 151274 549922 151342 549978
rect 151398 549922 168970 549978
rect 169026 549922 169094 549978
rect 169150 549922 169218 549978
rect 169274 549922 169342 549978
rect 169398 549922 186970 549978
rect 187026 549922 187094 549978
rect 187150 549922 187218 549978
rect 187274 549922 187342 549978
rect 187398 549922 204970 549978
rect 205026 549922 205094 549978
rect 205150 549922 205218 549978
rect 205274 549922 205342 549978
rect 205398 549922 222970 549978
rect 223026 549922 223094 549978
rect 223150 549922 223218 549978
rect 223274 549922 223342 549978
rect 223398 549922 240970 549978
rect 241026 549922 241094 549978
rect 241150 549922 241218 549978
rect 241274 549922 241342 549978
rect 241398 549922 258970 549978
rect 259026 549922 259094 549978
rect 259150 549922 259218 549978
rect 259274 549922 259342 549978
rect 259398 549922 276970 549978
rect 277026 549922 277094 549978
rect 277150 549922 277218 549978
rect 277274 549922 277342 549978
rect 277398 549922 294970 549978
rect 295026 549922 295094 549978
rect 295150 549922 295218 549978
rect 295274 549922 295342 549978
rect 295398 549922 312970 549978
rect 313026 549922 313094 549978
rect 313150 549922 313218 549978
rect 313274 549922 313342 549978
rect 313398 549922 330970 549978
rect 331026 549922 331094 549978
rect 331150 549922 331218 549978
rect 331274 549922 331342 549978
rect 331398 549922 348970 549978
rect 349026 549922 349094 549978
rect 349150 549922 349218 549978
rect 349274 549922 349342 549978
rect 349398 549922 366970 549978
rect 367026 549922 367094 549978
rect 367150 549922 367218 549978
rect 367274 549922 367342 549978
rect 367398 549922 384970 549978
rect 385026 549922 385094 549978
rect 385150 549922 385218 549978
rect 385274 549922 385342 549978
rect 385398 549922 402970 549978
rect 403026 549922 403094 549978
rect 403150 549922 403218 549978
rect 403274 549922 403342 549978
rect 403398 549922 420970 549978
rect 421026 549922 421094 549978
rect 421150 549922 421218 549978
rect 421274 549922 421342 549978
rect 421398 549922 438970 549978
rect 439026 549922 439094 549978
rect 439150 549922 439218 549978
rect 439274 549922 439342 549978
rect 439398 549922 456970 549978
rect 457026 549922 457094 549978
rect 457150 549922 457218 549978
rect 457274 549922 457342 549978
rect 457398 549922 474970 549978
rect 475026 549922 475094 549978
rect 475150 549922 475218 549978
rect 475274 549922 475342 549978
rect 475398 549922 492970 549978
rect 493026 549922 493094 549978
rect 493150 549922 493218 549978
rect 493274 549922 493342 549978
rect 493398 549922 510970 549978
rect 511026 549922 511094 549978
rect 511150 549922 511218 549978
rect 511274 549922 511342 549978
rect 511398 549922 528970 549978
rect 529026 549922 529094 549978
rect 529150 549922 529218 549978
rect 529274 549922 529342 549978
rect 529398 549922 546970 549978
rect 547026 549922 547094 549978
rect 547150 549922 547218 549978
rect 547274 549922 547342 549978
rect 547398 549922 564970 549978
rect 565026 549922 565094 549978
rect 565150 549922 565218 549978
rect 565274 549922 565342 549978
rect 565398 549922 582970 549978
rect 583026 549922 583094 549978
rect 583150 549922 583218 549978
rect 583274 549922 583342 549978
rect 583398 549922 597456 549978
rect 597512 549922 597580 549978
rect 597636 549922 597704 549978
rect 597760 549922 597828 549978
rect 597884 549922 597980 549978
rect -1916 549826 597980 549922
rect -1916 544350 597980 544446
rect -1916 544294 -860 544350
rect -804 544294 -736 544350
rect -680 544294 -612 544350
rect -556 544294 -488 544350
rect -432 544294 3250 544350
rect 3306 544294 3374 544350
rect 3430 544294 3498 544350
rect 3554 544294 3622 544350
rect 3678 544294 21250 544350
rect 21306 544294 21374 544350
rect 21430 544294 21498 544350
rect 21554 544294 21622 544350
rect 21678 544294 39250 544350
rect 39306 544294 39374 544350
rect 39430 544294 39498 544350
rect 39554 544294 39622 544350
rect 39678 544294 57250 544350
rect 57306 544294 57374 544350
rect 57430 544294 57498 544350
rect 57554 544294 57622 544350
rect 57678 544294 75250 544350
rect 75306 544294 75374 544350
rect 75430 544294 75498 544350
rect 75554 544294 75622 544350
rect 75678 544294 93250 544350
rect 93306 544294 93374 544350
rect 93430 544294 93498 544350
rect 93554 544294 93622 544350
rect 93678 544294 111250 544350
rect 111306 544294 111374 544350
rect 111430 544294 111498 544350
rect 111554 544294 111622 544350
rect 111678 544294 129250 544350
rect 129306 544294 129374 544350
rect 129430 544294 129498 544350
rect 129554 544294 129622 544350
rect 129678 544294 147250 544350
rect 147306 544294 147374 544350
rect 147430 544294 147498 544350
rect 147554 544294 147622 544350
rect 147678 544294 165250 544350
rect 165306 544294 165374 544350
rect 165430 544294 165498 544350
rect 165554 544294 165622 544350
rect 165678 544294 183250 544350
rect 183306 544294 183374 544350
rect 183430 544294 183498 544350
rect 183554 544294 183622 544350
rect 183678 544294 201250 544350
rect 201306 544294 201374 544350
rect 201430 544294 201498 544350
rect 201554 544294 201622 544350
rect 201678 544294 219250 544350
rect 219306 544294 219374 544350
rect 219430 544294 219498 544350
rect 219554 544294 219622 544350
rect 219678 544294 237250 544350
rect 237306 544294 237374 544350
rect 237430 544294 237498 544350
rect 237554 544294 237622 544350
rect 237678 544294 255250 544350
rect 255306 544294 255374 544350
rect 255430 544294 255498 544350
rect 255554 544294 255622 544350
rect 255678 544294 273250 544350
rect 273306 544294 273374 544350
rect 273430 544294 273498 544350
rect 273554 544294 273622 544350
rect 273678 544294 291250 544350
rect 291306 544294 291374 544350
rect 291430 544294 291498 544350
rect 291554 544294 291622 544350
rect 291678 544294 309250 544350
rect 309306 544294 309374 544350
rect 309430 544294 309498 544350
rect 309554 544294 309622 544350
rect 309678 544294 327250 544350
rect 327306 544294 327374 544350
rect 327430 544294 327498 544350
rect 327554 544294 327622 544350
rect 327678 544294 345250 544350
rect 345306 544294 345374 544350
rect 345430 544294 345498 544350
rect 345554 544294 345622 544350
rect 345678 544294 363250 544350
rect 363306 544294 363374 544350
rect 363430 544294 363498 544350
rect 363554 544294 363622 544350
rect 363678 544294 381250 544350
rect 381306 544294 381374 544350
rect 381430 544294 381498 544350
rect 381554 544294 381622 544350
rect 381678 544294 399250 544350
rect 399306 544294 399374 544350
rect 399430 544294 399498 544350
rect 399554 544294 399622 544350
rect 399678 544294 417250 544350
rect 417306 544294 417374 544350
rect 417430 544294 417498 544350
rect 417554 544294 417622 544350
rect 417678 544294 435250 544350
rect 435306 544294 435374 544350
rect 435430 544294 435498 544350
rect 435554 544294 435622 544350
rect 435678 544294 453250 544350
rect 453306 544294 453374 544350
rect 453430 544294 453498 544350
rect 453554 544294 453622 544350
rect 453678 544294 471250 544350
rect 471306 544294 471374 544350
rect 471430 544294 471498 544350
rect 471554 544294 471622 544350
rect 471678 544294 489250 544350
rect 489306 544294 489374 544350
rect 489430 544294 489498 544350
rect 489554 544294 489622 544350
rect 489678 544294 507250 544350
rect 507306 544294 507374 544350
rect 507430 544294 507498 544350
rect 507554 544294 507622 544350
rect 507678 544294 525250 544350
rect 525306 544294 525374 544350
rect 525430 544294 525498 544350
rect 525554 544294 525622 544350
rect 525678 544294 543250 544350
rect 543306 544294 543374 544350
rect 543430 544294 543498 544350
rect 543554 544294 543622 544350
rect 543678 544294 561250 544350
rect 561306 544294 561374 544350
rect 561430 544294 561498 544350
rect 561554 544294 561622 544350
rect 561678 544294 579250 544350
rect 579306 544294 579374 544350
rect 579430 544294 579498 544350
rect 579554 544294 579622 544350
rect 579678 544294 596496 544350
rect 596552 544294 596620 544350
rect 596676 544294 596744 544350
rect 596800 544294 596868 544350
rect 596924 544294 597980 544350
rect -1916 544226 597980 544294
rect -1916 544170 -860 544226
rect -804 544170 -736 544226
rect -680 544170 -612 544226
rect -556 544170 -488 544226
rect -432 544170 3250 544226
rect 3306 544170 3374 544226
rect 3430 544170 3498 544226
rect 3554 544170 3622 544226
rect 3678 544170 21250 544226
rect 21306 544170 21374 544226
rect 21430 544170 21498 544226
rect 21554 544170 21622 544226
rect 21678 544170 39250 544226
rect 39306 544170 39374 544226
rect 39430 544170 39498 544226
rect 39554 544170 39622 544226
rect 39678 544170 57250 544226
rect 57306 544170 57374 544226
rect 57430 544170 57498 544226
rect 57554 544170 57622 544226
rect 57678 544170 75250 544226
rect 75306 544170 75374 544226
rect 75430 544170 75498 544226
rect 75554 544170 75622 544226
rect 75678 544170 93250 544226
rect 93306 544170 93374 544226
rect 93430 544170 93498 544226
rect 93554 544170 93622 544226
rect 93678 544170 111250 544226
rect 111306 544170 111374 544226
rect 111430 544170 111498 544226
rect 111554 544170 111622 544226
rect 111678 544170 129250 544226
rect 129306 544170 129374 544226
rect 129430 544170 129498 544226
rect 129554 544170 129622 544226
rect 129678 544170 147250 544226
rect 147306 544170 147374 544226
rect 147430 544170 147498 544226
rect 147554 544170 147622 544226
rect 147678 544170 165250 544226
rect 165306 544170 165374 544226
rect 165430 544170 165498 544226
rect 165554 544170 165622 544226
rect 165678 544170 183250 544226
rect 183306 544170 183374 544226
rect 183430 544170 183498 544226
rect 183554 544170 183622 544226
rect 183678 544170 201250 544226
rect 201306 544170 201374 544226
rect 201430 544170 201498 544226
rect 201554 544170 201622 544226
rect 201678 544170 219250 544226
rect 219306 544170 219374 544226
rect 219430 544170 219498 544226
rect 219554 544170 219622 544226
rect 219678 544170 237250 544226
rect 237306 544170 237374 544226
rect 237430 544170 237498 544226
rect 237554 544170 237622 544226
rect 237678 544170 255250 544226
rect 255306 544170 255374 544226
rect 255430 544170 255498 544226
rect 255554 544170 255622 544226
rect 255678 544170 273250 544226
rect 273306 544170 273374 544226
rect 273430 544170 273498 544226
rect 273554 544170 273622 544226
rect 273678 544170 291250 544226
rect 291306 544170 291374 544226
rect 291430 544170 291498 544226
rect 291554 544170 291622 544226
rect 291678 544170 309250 544226
rect 309306 544170 309374 544226
rect 309430 544170 309498 544226
rect 309554 544170 309622 544226
rect 309678 544170 327250 544226
rect 327306 544170 327374 544226
rect 327430 544170 327498 544226
rect 327554 544170 327622 544226
rect 327678 544170 345250 544226
rect 345306 544170 345374 544226
rect 345430 544170 345498 544226
rect 345554 544170 345622 544226
rect 345678 544170 363250 544226
rect 363306 544170 363374 544226
rect 363430 544170 363498 544226
rect 363554 544170 363622 544226
rect 363678 544170 381250 544226
rect 381306 544170 381374 544226
rect 381430 544170 381498 544226
rect 381554 544170 381622 544226
rect 381678 544170 399250 544226
rect 399306 544170 399374 544226
rect 399430 544170 399498 544226
rect 399554 544170 399622 544226
rect 399678 544170 417250 544226
rect 417306 544170 417374 544226
rect 417430 544170 417498 544226
rect 417554 544170 417622 544226
rect 417678 544170 435250 544226
rect 435306 544170 435374 544226
rect 435430 544170 435498 544226
rect 435554 544170 435622 544226
rect 435678 544170 453250 544226
rect 453306 544170 453374 544226
rect 453430 544170 453498 544226
rect 453554 544170 453622 544226
rect 453678 544170 471250 544226
rect 471306 544170 471374 544226
rect 471430 544170 471498 544226
rect 471554 544170 471622 544226
rect 471678 544170 489250 544226
rect 489306 544170 489374 544226
rect 489430 544170 489498 544226
rect 489554 544170 489622 544226
rect 489678 544170 507250 544226
rect 507306 544170 507374 544226
rect 507430 544170 507498 544226
rect 507554 544170 507622 544226
rect 507678 544170 525250 544226
rect 525306 544170 525374 544226
rect 525430 544170 525498 544226
rect 525554 544170 525622 544226
rect 525678 544170 543250 544226
rect 543306 544170 543374 544226
rect 543430 544170 543498 544226
rect 543554 544170 543622 544226
rect 543678 544170 561250 544226
rect 561306 544170 561374 544226
rect 561430 544170 561498 544226
rect 561554 544170 561622 544226
rect 561678 544170 579250 544226
rect 579306 544170 579374 544226
rect 579430 544170 579498 544226
rect 579554 544170 579622 544226
rect 579678 544170 596496 544226
rect 596552 544170 596620 544226
rect 596676 544170 596744 544226
rect 596800 544170 596868 544226
rect 596924 544170 597980 544226
rect -1916 544102 597980 544170
rect -1916 544046 -860 544102
rect -804 544046 -736 544102
rect -680 544046 -612 544102
rect -556 544046 -488 544102
rect -432 544046 3250 544102
rect 3306 544046 3374 544102
rect 3430 544046 3498 544102
rect 3554 544046 3622 544102
rect 3678 544046 21250 544102
rect 21306 544046 21374 544102
rect 21430 544046 21498 544102
rect 21554 544046 21622 544102
rect 21678 544046 39250 544102
rect 39306 544046 39374 544102
rect 39430 544046 39498 544102
rect 39554 544046 39622 544102
rect 39678 544046 57250 544102
rect 57306 544046 57374 544102
rect 57430 544046 57498 544102
rect 57554 544046 57622 544102
rect 57678 544046 75250 544102
rect 75306 544046 75374 544102
rect 75430 544046 75498 544102
rect 75554 544046 75622 544102
rect 75678 544046 93250 544102
rect 93306 544046 93374 544102
rect 93430 544046 93498 544102
rect 93554 544046 93622 544102
rect 93678 544046 111250 544102
rect 111306 544046 111374 544102
rect 111430 544046 111498 544102
rect 111554 544046 111622 544102
rect 111678 544046 129250 544102
rect 129306 544046 129374 544102
rect 129430 544046 129498 544102
rect 129554 544046 129622 544102
rect 129678 544046 147250 544102
rect 147306 544046 147374 544102
rect 147430 544046 147498 544102
rect 147554 544046 147622 544102
rect 147678 544046 165250 544102
rect 165306 544046 165374 544102
rect 165430 544046 165498 544102
rect 165554 544046 165622 544102
rect 165678 544046 183250 544102
rect 183306 544046 183374 544102
rect 183430 544046 183498 544102
rect 183554 544046 183622 544102
rect 183678 544046 201250 544102
rect 201306 544046 201374 544102
rect 201430 544046 201498 544102
rect 201554 544046 201622 544102
rect 201678 544046 219250 544102
rect 219306 544046 219374 544102
rect 219430 544046 219498 544102
rect 219554 544046 219622 544102
rect 219678 544046 237250 544102
rect 237306 544046 237374 544102
rect 237430 544046 237498 544102
rect 237554 544046 237622 544102
rect 237678 544046 255250 544102
rect 255306 544046 255374 544102
rect 255430 544046 255498 544102
rect 255554 544046 255622 544102
rect 255678 544046 273250 544102
rect 273306 544046 273374 544102
rect 273430 544046 273498 544102
rect 273554 544046 273622 544102
rect 273678 544046 291250 544102
rect 291306 544046 291374 544102
rect 291430 544046 291498 544102
rect 291554 544046 291622 544102
rect 291678 544046 309250 544102
rect 309306 544046 309374 544102
rect 309430 544046 309498 544102
rect 309554 544046 309622 544102
rect 309678 544046 327250 544102
rect 327306 544046 327374 544102
rect 327430 544046 327498 544102
rect 327554 544046 327622 544102
rect 327678 544046 345250 544102
rect 345306 544046 345374 544102
rect 345430 544046 345498 544102
rect 345554 544046 345622 544102
rect 345678 544046 363250 544102
rect 363306 544046 363374 544102
rect 363430 544046 363498 544102
rect 363554 544046 363622 544102
rect 363678 544046 381250 544102
rect 381306 544046 381374 544102
rect 381430 544046 381498 544102
rect 381554 544046 381622 544102
rect 381678 544046 399250 544102
rect 399306 544046 399374 544102
rect 399430 544046 399498 544102
rect 399554 544046 399622 544102
rect 399678 544046 417250 544102
rect 417306 544046 417374 544102
rect 417430 544046 417498 544102
rect 417554 544046 417622 544102
rect 417678 544046 435250 544102
rect 435306 544046 435374 544102
rect 435430 544046 435498 544102
rect 435554 544046 435622 544102
rect 435678 544046 453250 544102
rect 453306 544046 453374 544102
rect 453430 544046 453498 544102
rect 453554 544046 453622 544102
rect 453678 544046 471250 544102
rect 471306 544046 471374 544102
rect 471430 544046 471498 544102
rect 471554 544046 471622 544102
rect 471678 544046 489250 544102
rect 489306 544046 489374 544102
rect 489430 544046 489498 544102
rect 489554 544046 489622 544102
rect 489678 544046 507250 544102
rect 507306 544046 507374 544102
rect 507430 544046 507498 544102
rect 507554 544046 507622 544102
rect 507678 544046 525250 544102
rect 525306 544046 525374 544102
rect 525430 544046 525498 544102
rect 525554 544046 525622 544102
rect 525678 544046 543250 544102
rect 543306 544046 543374 544102
rect 543430 544046 543498 544102
rect 543554 544046 543622 544102
rect 543678 544046 561250 544102
rect 561306 544046 561374 544102
rect 561430 544046 561498 544102
rect 561554 544046 561622 544102
rect 561678 544046 579250 544102
rect 579306 544046 579374 544102
rect 579430 544046 579498 544102
rect 579554 544046 579622 544102
rect 579678 544046 596496 544102
rect 596552 544046 596620 544102
rect 596676 544046 596744 544102
rect 596800 544046 596868 544102
rect 596924 544046 597980 544102
rect -1916 543978 597980 544046
rect -1916 543922 -860 543978
rect -804 543922 -736 543978
rect -680 543922 -612 543978
rect -556 543922 -488 543978
rect -432 543922 3250 543978
rect 3306 543922 3374 543978
rect 3430 543922 3498 543978
rect 3554 543922 3622 543978
rect 3678 543922 21250 543978
rect 21306 543922 21374 543978
rect 21430 543922 21498 543978
rect 21554 543922 21622 543978
rect 21678 543922 39250 543978
rect 39306 543922 39374 543978
rect 39430 543922 39498 543978
rect 39554 543922 39622 543978
rect 39678 543922 57250 543978
rect 57306 543922 57374 543978
rect 57430 543922 57498 543978
rect 57554 543922 57622 543978
rect 57678 543922 75250 543978
rect 75306 543922 75374 543978
rect 75430 543922 75498 543978
rect 75554 543922 75622 543978
rect 75678 543922 93250 543978
rect 93306 543922 93374 543978
rect 93430 543922 93498 543978
rect 93554 543922 93622 543978
rect 93678 543922 111250 543978
rect 111306 543922 111374 543978
rect 111430 543922 111498 543978
rect 111554 543922 111622 543978
rect 111678 543922 129250 543978
rect 129306 543922 129374 543978
rect 129430 543922 129498 543978
rect 129554 543922 129622 543978
rect 129678 543922 147250 543978
rect 147306 543922 147374 543978
rect 147430 543922 147498 543978
rect 147554 543922 147622 543978
rect 147678 543922 165250 543978
rect 165306 543922 165374 543978
rect 165430 543922 165498 543978
rect 165554 543922 165622 543978
rect 165678 543922 183250 543978
rect 183306 543922 183374 543978
rect 183430 543922 183498 543978
rect 183554 543922 183622 543978
rect 183678 543922 201250 543978
rect 201306 543922 201374 543978
rect 201430 543922 201498 543978
rect 201554 543922 201622 543978
rect 201678 543922 219250 543978
rect 219306 543922 219374 543978
rect 219430 543922 219498 543978
rect 219554 543922 219622 543978
rect 219678 543922 237250 543978
rect 237306 543922 237374 543978
rect 237430 543922 237498 543978
rect 237554 543922 237622 543978
rect 237678 543922 255250 543978
rect 255306 543922 255374 543978
rect 255430 543922 255498 543978
rect 255554 543922 255622 543978
rect 255678 543922 273250 543978
rect 273306 543922 273374 543978
rect 273430 543922 273498 543978
rect 273554 543922 273622 543978
rect 273678 543922 291250 543978
rect 291306 543922 291374 543978
rect 291430 543922 291498 543978
rect 291554 543922 291622 543978
rect 291678 543922 309250 543978
rect 309306 543922 309374 543978
rect 309430 543922 309498 543978
rect 309554 543922 309622 543978
rect 309678 543922 327250 543978
rect 327306 543922 327374 543978
rect 327430 543922 327498 543978
rect 327554 543922 327622 543978
rect 327678 543922 345250 543978
rect 345306 543922 345374 543978
rect 345430 543922 345498 543978
rect 345554 543922 345622 543978
rect 345678 543922 363250 543978
rect 363306 543922 363374 543978
rect 363430 543922 363498 543978
rect 363554 543922 363622 543978
rect 363678 543922 381250 543978
rect 381306 543922 381374 543978
rect 381430 543922 381498 543978
rect 381554 543922 381622 543978
rect 381678 543922 399250 543978
rect 399306 543922 399374 543978
rect 399430 543922 399498 543978
rect 399554 543922 399622 543978
rect 399678 543922 417250 543978
rect 417306 543922 417374 543978
rect 417430 543922 417498 543978
rect 417554 543922 417622 543978
rect 417678 543922 435250 543978
rect 435306 543922 435374 543978
rect 435430 543922 435498 543978
rect 435554 543922 435622 543978
rect 435678 543922 453250 543978
rect 453306 543922 453374 543978
rect 453430 543922 453498 543978
rect 453554 543922 453622 543978
rect 453678 543922 471250 543978
rect 471306 543922 471374 543978
rect 471430 543922 471498 543978
rect 471554 543922 471622 543978
rect 471678 543922 489250 543978
rect 489306 543922 489374 543978
rect 489430 543922 489498 543978
rect 489554 543922 489622 543978
rect 489678 543922 507250 543978
rect 507306 543922 507374 543978
rect 507430 543922 507498 543978
rect 507554 543922 507622 543978
rect 507678 543922 525250 543978
rect 525306 543922 525374 543978
rect 525430 543922 525498 543978
rect 525554 543922 525622 543978
rect 525678 543922 543250 543978
rect 543306 543922 543374 543978
rect 543430 543922 543498 543978
rect 543554 543922 543622 543978
rect 543678 543922 561250 543978
rect 561306 543922 561374 543978
rect 561430 543922 561498 543978
rect 561554 543922 561622 543978
rect 561678 543922 579250 543978
rect 579306 543922 579374 543978
rect 579430 543922 579498 543978
rect 579554 543922 579622 543978
rect 579678 543922 596496 543978
rect 596552 543922 596620 543978
rect 596676 543922 596744 543978
rect 596800 543922 596868 543978
rect 596924 543922 597980 543978
rect -1916 543826 597980 543922
rect -1916 532350 597980 532446
rect -1916 532294 -1820 532350
rect -1764 532294 -1696 532350
rect -1640 532294 -1572 532350
rect -1516 532294 -1448 532350
rect -1392 532294 6970 532350
rect 7026 532294 7094 532350
rect 7150 532294 7218 532350
rect 7274 532294 7342 532350
rect 7398 532294 24970 532350
rect 25026 532294 25094 532350
rect 25150 532294 25218 532350
rect 25274 532294 25342 532350
rect 25398 532294 42970 532350
rect 43026 532294 43094 532350
rect 43150 532294 43218 532350
rect 43274 532294 43342 532350
rect 43398 532294 60970 532350
rect 61026 532294 61094 532350
rect 61150 532294 61218 532350
rect 61274 532294 61342 532350
rect 61398 532294 78970 532350
rect 79026 532294 79094 532350
rect 79150 532294 79218 532350
rect 79274 532294 79342 532350
rect 79398 532294 96970 532350
rect 97026 532294 97094 532350
rect 97150 532294 97218 532350
rect 97274 532294 97342 532350
rect 97398 532294 114970 532350
rect 115026 532294 115094 532350
rect 115150 532294 115218 532350
rect 115274 532294 115342 532350
rect 115398 532294 132970 532350
rect 133026 532294 133094 532350
rect 133150 532294 133218 532350
rect 133274 532294 133342 532350
rect 133398 532294 150970 532350
rect 151026 532294 151094 532350
rect 151150 532294 151218 532350
rect 151274 532294 151342 532350
rect 151398 532294 168970 532350
rect 169026 532294 169094 532350
rect 169150 532294 169218 532350
rect 169274 532294 169342 532350
rect 169398 532294 186970 532350
rect 187026 532294 187094 532350
rect 187150 532294 187218 532350
rect 187274 532294 187342 532350
rect 187398 532294 204970 532350
rect 205026 532294 205094 532350
rect 205150 532294 205218 532350
rect 205274 532294 205342 532350
rect 205398 532294 222970 532350
rect 223026 532294 223094 532350
rect 223150 532294 223218 532350
rect 223274 532294 223342 532350
rect 223398 532294 240970 532350
rect 241026 532294 241094 532350
rect 241150 532294 241218 532350
rect 241274 532294 241342 532350
rect 241398 532294 258970 532350
rect 259026 532294 259094 532350
rect 259150 532294 259218 532350
rect 259274 532294 259342 532350
rect 259398 532294 276970 532350
rect 277026 532294 277094 532350
rect 277150 532294 277218 532350
rect 277274 532294 277342 532350
rect 277398 532294 294970 532350
rect 295026 532294 295094 532350
rect 295150 532294 295218 532350
rect 295274 532294 295342 532350
rect 295398 532294 312970 532350
rect 313026 532294 313094 532350
rect 313150 532294 313218 532350
rect 313274 532294 313342 532350
rect 313398 532294 330970 532350
rect 331026 532294 331094 532350
rect 331150 532294 331218 532350
rect 331274 532294 331342 532350
rect 331398 532294 348970 532350
rect 349026 532294 349094 532350
rect 349150 532294 349218 532350
rect 349274 532294 349342 532350
rect 349398 532294 366970 532350
rect 367026 532294 367094 532350
rect 367150 532294 367218 532350
rect 367274 532294 367342 532350
rect 367398 532294 384970 532350
rect 385026 532294 385094 532350
rect 385150 532294 385218 532350
rect 385274 532294 385342 532350
rect 385398 532294 402970 532350
rect 403026 532294 403094 532350
rect 403150 532294 403218 532350
rect 403274 532294 403342 532350
rect 403398 532294 420970 532350
rect 421026 532294 421094 532350
rect 421150 532294 421218 532350
rect 421274 532294 421342 532350
rect 421398 532294 438970 532350
rect 439026 532294 439094 532350
rect 439150 532294 439218 532350
rect 439274 532294 439342 532350
rect 439398 532294 456970 532350
rect 457026 532294 457094 532350
rect 457150 532294 457218 532350
rect 457274 532294 457342 532350
rect 457398 532294 474970 532350
rect 475026 532294 475094 532350
rect 475150 532294 475218 532350
rect 475274 532294 475342 532350
rect 475398 532294 492970 532350
rect 493026 532294 493094 532350
rect 493150 532294 493218 532350
rect 493274 532294 493342 532350
rect 493398 532294 510970 532350
rect 511026 532294 511094 532350
rect 511150 532294 511218 532350
rect 511274 532294 511342 532350
rect 511398 532294 528970 532350
rect 529026 532294 529094 532350
rect 529150 532294 529218 532350
rect 529274 532294 529342 532350
rect 529398 532294 546970 532350
rect 547026 532294 547094 532350
rect 547150 532294 547218 532350
rect 547274 532294 547342 532350
rect 547398 532294 564970 532350
rect 565026 532294 565094 532350
rect 565150 532294 565218 532350
rect 565274 532294 565342 532350
rect 565398 532294 582970 532350
rect 583026 532294 583094 532350
rect 583150 532294 583218 532350
rect 583274 532294 583342 532350
rect 583398 532294 597456 532350
rect 597512 532294 597580 532350
rect 597636 532294 597704 532350
rect 597760 532294 597828 532350
rect 597884 532294 597980 532350
rect -1916 532226 597980 532294
rect -1916 532170 -1820 532226
rect -1764 532170 -1696 532226
rect -1640 532170 -1572 532226
rect -1516 532170 -1448 532226
rect -1392 532170 6970 532226
rect 7026 532170 7094 532226
rect 7150 532170 7218 532226
rect 7274 532170 7342 532226
rect 7398 532170 24970 532226
rect 25026 532170 25094 532226
rect 25150 532170 25218 532226
rect 25274 532170 25342 532226
rect 25398 532170 42970 532226
rect 43026 532170 43094 532226
rect 43150 532170 43218 532226
rect 43274 532170 43342 532226
rect 43398 532170 60970 532226
rect 61026 532170 61094 532226
rect 61150 532170 61218 532226
rect 61274 532170 61342 532226
rect 61398 532170 78970 532226
rect 79026 532170 79094 532226
rect 79150 532170 79218 532226
rect 79274 532170 79342 532226
rect 79398 532170 96970 532226
rect 97026 532170 97094 532226
rect 97150 532170 97218 532226
rect 97274 532170 97342 532226
rect 97398 532170 114970 532226
rect 115026 532170 115094 532226
rect 115150 532170 115218 532226
rect 115274 532170 115342 532226
rect 115398 532170 132970 532226
rect 133026 532170 133094 532226
rect 133150 532170 133218 532226
rect 133274 532170 133342 532226
rect 133398 532170 150970 532226
rect 151026 532170 151094 532226
rect 151150 532170 151218 532226
rect 151274 532170 151342 532226
rect 151398 532170 168970 532226
rect 169026 532170 169094 532226
rect 169150 532170 169218 532226
rect 169274 532170 169342 532226
rect 169398 532170 186970 532226
rect 187026 532170 187094 532226
rect 187150 532170 187218 532226
rect 187274 532170 187342 532226
rect 187398 532170 204970 532226
rect 205026 532170 205094 532226
rect 205150 532170 205218 532226
rect 205274 532170 205342 532226
rect 205398 532170 222970 532226
rect 223026 532170 223094 532226
rect 223150 532170 223218 532226
rect 223274 532170 223342 532226
rect 223398 532170 240970 532226
rect 241026 532170 241094 532226
rect 241150 532170 241218 532226
rect 241274 532170 241342 532226
rect 241398 532170 258970 532226
rect 259026 532170 259094 532226
rect 259150 532170 259218 532226
rect 259274 532170 259342 532226
rect 259398 532170 276970 532226
rect 277026 532170 277094 532226
rect 277150 532170 277218 532226
rect 277274 532170 277342 532226
rect 277398 532170 294970 532226
rect 295026 532170 295094 532226
rect 295150 532170 295218 532226
rect 295274 532170 295342 532226
rect 295398 532170 312970 532226
rect 313026 532170 313094 532226
rect 313150 532170 313218 532226
rect 313274 532170 313342 532226
rect 313398 532170 330970 532226
rect 331026 532170 331094 532226
rect 331150 532170 331218 532226
rect 331274 532170 331342 532226
rect 331398 532170 348970 532226
rect 349026 532170 349094 532226
rect 349150 532170 349218 532226
rect 349274 532170 349342 532226
rect 349398 532170 366970 532226
rect 367026 532170 367094 532226
rect 367150 532170 367218 532226
rect 367274 532170 367342 532226
rect 367398 532170 384970 532226
rect 385026 532170 385094 532226
rect 385150 532170 385218 532226
rect 385274 532170 385342 532226
rect 385398 532170 402970 532226
rect 403026 532170 403094 532226
rect 403150 532170 403218 532226
rect 403274 532170 403342 532226
rect 403398 532170 420970 532226
rect 421026 532170 421094 532226
rect 421150 532170 421218 532226
rect 421274 532170 421342 532226
rect 421398 532170 438970 532226
rect 439026 532170 439094 532226
rect 439150 532170 439218 532226
rect 439274 532170 439342 532226
rect 439398 532170 456970 532226
rect 457026 532170 457094 532226
rect 457150 532170 457218 532226
rect 457274 532170 457342 532226
rect 457398 532170 474970 532226
rect 475026 532170 475094 532226
rect 475150 532170 475218 532226
rect 475274 532170 475342 532226
rect 475398 532170 492970 532226
rect 493026 532170 493094 532226
rect 493150 532170 493218 532226
rect 493274 532170 493342 532226
rect 493398 532170 510970 532226
rect 511026 532170 511094 532226
rect 511150 532170 511218 532226
rect 511274 532170 511342 532226
rect 511398 532170 528970 532226
rect 529026 532170 529094 532226
rect 529150 532170 529218 532226
rect 529274 532170 529342 532226
rect 529398 532170 546970 532226
rect 547026 532170 547094 532226
rect 547150 532170 547218 532226
rect 547274 532170 547342 532226
rect 547398 532170 564970 532226
rect 565026 532170 565094 532226
rect 565150 532170 565218 532226
rect 565274 532170 565342 532226
rect 565398 532170 582970 532226
rect 583026 532170 583094 532226
rect 583150 532170 583218 532226
rect 583274 532170 583342 532226
rect 583398 532170 597456 532226
rect 597512 532170 597580 532226
rect 597636 532170 597704 532226
rect 597760 532170 597828 532226
rect 597884 532170 597980 532226
rect -1916 532102 597980 532170
rect -1916 532046 -1820 532102
rect -1764 532046 -1696 532102
rect -1640 532046 -1572 532102
rect -1516 532046 -1448 532102
rect -1392 532046 6970 532102
rect 7026 532046 7094 532102
rect 7150 532046 7218 532102
rect 7274 532046 7342 532102
rect 7398 532046 24970 532102
rect 25026 532046 25094 532102
rect 25150 532046 25218 532102
rect 25274 532046 25342 532102
rect 25398 532046 42970 532102
rect 43026 532046 43094 532102
rect 43150 532046 43218 532102
rect 43274 532046 43342 532102
rect 43398 532046 60970 532102
rect 61026 532046 61094 532102
rect 61150 532046 61218 532102
rect 61274 532046 61342 532102
rect 61398 532046 78970 532102
rect 79026 532046 79094 532102
rect 79150 532046 79218 532102
rect 79274 532046 79342 532102
rect 79398 532046 96970 532102
rect 97026 532046 97094 532102
rect 97150 532046 97218 532102
rect 97274 532046 97342 532102
rect 97398 532046 114970 532102
rect 115026 532046 115094 532102
rect 115150 532046 115218 532102
rect 115274 532046 115342 532102
rect 115398 532046 132970 532102
rect 133026 532046 133094 532102
rect 133150 532046 133218 532102
rect 133274 532046 133342 532102
rect 133398 532046 150970 532102
rect 151026 532046 151094 532102
rect 151150 532046 151218 532102
rect 151274 532046 151342 532102
rect 151398 532046 168970 532102
rect 169026 532046 169094 532102
rect 169150 532046 169218 532102
rect 169274 532046 169342 532102
rect 169398 532046 186970 532102
rect 187026 532046 187094 532102
rect 187150 532046 187218 532102
rect 187274 532046 187342 532102
rect 187398 532046 204970 532102
rect 205026 532046 205094 532102
rect 205150 532046 205218 532102
rect 205274 532046 205342 532102
rect 205398 532046 222970 532102
rect 223026 532046 223094 532102
rect 223150 532046 223218 532102
rect 223274 532046 223342 532102
rect 223398 532046 240970 532102
rect 241026 532046 241094 532102
rect 241150 532046 241218 532102
rect 241274 532046 241342 532102
rect 241398 532046 258970 532102
rect 259026 532046 259094 532102
rect 259150 532046 259218 532102
rect 259274 532046 259342 532102
rect 259398 532046 276970 532102
rect 277026 532046 277094 532102
rect 277150 532046 277218 532102
rect 277274 532046 277342 532102
rect 277398 532046 294970 532102
rect 295026 532046 295094 532102
rect 295150 532046 295218 532102
rect 295274 532046 295342 532102
rect 295398 532046 312970 532102
rect 313026 532046 313094 532102
rect 313150 532046 313218 532102
rect 313274 532046 313342 532102
rect 313398 532046 330970 532102
rect 331026 532046 331094 532102
rect 331150 532046 331218 532102
rect 331274 532046 331342 532102
rect 331398 532046 348970 532102
rect 349026 532046 349094 532102
rect 349150 532046 349218 532102
rect 349274 532046 349342 532102
rect 349398 532046 366970 532102
rect 367026 532046 367094 532102
rect 367150 532046 367218 532102
rect 367274 532046 367342 532102
rect 367398 532046 384970 532102
rect 385026 532046 385094 532102
rect 385150 532046 385218 532102
rect 385274 532046 385342 532102
rect 385398 532046 402970 532102
rect 403026 532046 403094 532102
rect 403150 532046 403218 532102
rect 403274 532046 403342 532102
rect 403398 532046 420970 532102
rect 421026 532046 421094 532102
rect 421150 532046 421218 532102
rect 421274 532046 421342 532102
rect 421398 532046 438970 532102
rect 439026 532046 439094 532102
rect 439150 532046 439218 532102
rect 439274 532046 439342 532102
rect 439398 532046 456970 532102
rect 457026 532046 457094 532102
rect 457150 532046 457218 532102
rect 457274 532046 457342 532102
rect 457398 532046 474970 532102
rect 475026 532046 475094 532102
rect 475150 532046 475218 532102
rect 475274 532046 475342 532102
rect 475398 532046 492970 532102
rect 493026 532046 493094 532102
rect 493150 532046 493218 532102
rect 493274 532046 493342 532102
rect 493398 532046 510970 532102
rect 511026 532046 511094 532102
rect 511150 532046 511218 532102
rect 511274 532046 511342 532102
rect 511398 532046 528970 532102
rect 529026 532046 529094 532102
rect 529150 532046 529218 532102
rect 529274 532046 529342 532102
rect 529398 532046 546970 532102
rect 547026 532046 547094 532102
rect 547150 532046 547218 532102
rect 547274 532046 547342 532102
rect 547398 532046 564970 532102
rect 565026 532046 565094 532102
rect 565150 532046 565218 532102
rect 565274 532046 565342 532102
rect 565398 532046 582970 532102
rect 583026 532046 583094 532102
rect 583150 532046 583218 532102
rect 583274 532046 583342 532102
rect 583398 532046 597456 532102
rect 597512 532046 597580 532102
rect 597636 532046 597704 532102
rect 597760 532046 597828 532102
rect 597884 532046 597980 532102
rect -1916 531978 597980 532046
rect -1916 531922 -1820 531978
rect -1764 531922 -1696 531978
rect -1640 531922 -1572 531978
rect -1516 531922 -1448 531978
rect -1392 531922 6970 531978
rect 7026 531922 7094 531978
rect 7150 531922 7218 531978
rect 7274 531922 7342 531978
rect 7398 531922 24970 531978
rect 25026 531922 25094 531978
rect 25150 531922 25218 531978
rect 25274 531922 25342 531978
rect 25398 531922 42970 531978
rect 43026 531922 43094 531978
rect 43150 531922 43218 531978
rect 43274 531922 43342 531978
rect 43398 531922 60970 531978
rect 61026 531922 61094 531978
rect 61150 531922 61218 531978
rect 61274 531922 61342 531978
rect 61398 531922 78970 531978
rect 79026 531922 79094 531978
rect 79150 531922 79218 531978
rect 79274 531922 79342 531978
rect 79398 531922 96970 531978
rect 97026 531922 97094 531978
rect 97150 531922 97218 531978
rect 97274 531922 97342 531978
rect 97398 531922 114970 531978
rect 115026 531922 115094 531978
rect 115150 531922 115218 531978
rect 115274 531922 115342 531978
rect 115398 531922 132970 531978
rect 133026 531922 133094 531978
rect 133150 531922 133218 531978
rect 133274 531922 133342 531978
rect 133398 531922 150970 531978
rect 151026 531922 151094 531978
rect 151150 531922 151218 531978
rect 151274 531922 151342 531978
rect 151398 531922 168970 531978
rect 169026 531922 169094 531978
rect 169150 531922 169218 531978
rect 169274 531922 169342 531978
rect 169398 531922 186970 531978
rect 187026 531922 187094 531978
rect 187150 531922 187218 531978
rect 187274 531922 187342 531978
rect 187398 531922 204970 531978
rect 205026 531922 205094 531978
rect 205150 531922 205218 531978
rect 205274 531922 205342 531978
rect 205398 531922 222970 531978
rect 223026 531922 223094 531978
rect 223150 531922 223218 531978
rect 223274 531922 223342 531978
rect 223398 531922 240970 531978
rect 241026 531922 241094 531978
rect 241150 531922 241218 531978
rect 241274 531922 241342 531978
rect 241398 531922 258970 531978
rect 259026 531922 259094 531978
rect 259150 531922 259218 531978
rect 259274 531922 259342 531978
rect 259398 531922 276970 531978
rect 277026 531922 277094 531978
rect 277150 531922 277218 531978
rect 277274 531922 277342 531978
rect 277398 531922 294970 531978
rect 295026 531922 295094 531978
rect 295150 531922 295218 531978
rect 295274 531922 295342 531978
rect 295398 531922 312970 531978
rect 313026 531922 313094 531978
rect 313150 531922 313218 531978
rect 313274 531922 313342 531978
rect 313398 531922 330970 531978
rect 331026 531922 331094 531978
rect 331150 531922 331218 531978
rect 331274 531922 331342 531978
rect 331398 531922 348970 531978
rect 349026 531922 349094 531978
rect 349150 531922 349218 531978
rect 349274 531922 349342 531978
rect 349398 531922 366970 531978
rect 367026 531922 367094 531978
rect 367150 531922 367218 531978
rect 367274 531922 367342 531978
rect 367398 531922 384970 531978
rect 385026 531922 385094 531978
rect 385150 531922 385218 531978
rect 385274 531922 385342 531978
rect 385398 531922 402970 531978
rect 403026 531922 403094 531978
rect 403150 531922 403218 531978
rect 403274 531922 403342 531978
rect 403398 531922 420970 531978
rect 421026 531922 421094 531978
rect 421150 531922 421218 531978
rect 421274 531922 421342 531978
rect 421398 531922 438970 531978
rect 439026 531922 439094 531978
rect 439150 531922 439218 531978
rect 439274 531922 439342 531978
rect 439398 531922 456970 531978
rect 457026 531922 457094 531978
rect 457150 531922 457218 531978
rect 457274 531922 457342 531978
rect 457398 531922 474970 531978
rect 475026 531922 475094 531978
rect 475150 531922 475218 531978
rect 475274 531922 475342 531978
rect 475398 531922 492970 531978
rect 493026 531922 493094 531978
rect 493150 531922 493218 531978
rect 493274 531922 493342 531978
rect 493398 531922 510970 531978
rect 511026 531922 511094 531978
rect 511150 531922 511218 531978
rect 511274 531922 511342 531978
rect 511398 531922 528970 531978
rect 529026 531922 529094 531978
rect 529150 531922 529218 531978
rect 529274 531922 529342 531978
rect 529398 531922 546970 531978
rect 547026 531922 547094 531978
rect 547150 531922 547218 531978
rect 547274 531922 547342 531978
rect 547398 531922 564970 531978
rect 565026 531922 565094 531978
rect 565150 531922 565218 531978
rect 565274 531922 565342 531978
rect 565398 531922 582970 531978
rect 583026 531922 583094 531978
rect 583150 531922 583218 531978
rect 583274 531922 583342 531978
rect 583398 531922 597456 531978
rect 597512 531922 597580 531978
rect 597636 531922 597704 531978
rect 597760 531922 597828 531978
rect 597884 531922 597980 531978
rect -1916 531826 597980 531922
rect -1916 526350 597980 526446
rect -1916 526294 -860 526350
rect -804 526294 -736 526350
rect -680 526294 -612 526350
rect -556 526294 -488 526350
rect -432 526294 3250 526350
rect 3306 526294 3374 526350
rect 3430 526294 3498 526350
rect 3554 526294 3622 526350
rect 3678 526294 21250 526350
rect 21306 526294 21374 526350
rect 21430 526294 21498 526350
rect 21554 526294 21622 526350
rect 21678 526294 39250 526350
rect 39306 526294 39374 526350
rect 39430 526294 39498 526350
rect 39554 526294 39622 526350
rect 39678 526294 57250 526350
rect 57306 526294 57374 526350
rect 57430 526294 57498 526350
rect 57554 526294 57622 526350
rect 57678 526294 75250 526350
rect 75306 526294 75374 526350
rect 75430 526294 75498 526350
rect 75554 526294 75622 526350
rect 75678 526294 93250 526350
rect 93306 526294 93374 526350
rect 93430 526294 93498 526350
rect 93554 526294 93622 526350
rect 93678 526294 111250 526350
rect 111306 526294 111374 526350
rect 111430 526294 111498 526350
rect 111554 526294 111622 526350
rect 111678 526294 129250 526350
rect 129306 526294 129374 526350
rect 129430 526294 129498 526350
rect 129554 526294 129622 526350
rect 129678 526294 147250 526350
rect 147306 526294 147374 526350
rect 147430 526294 147498 526350
rect 147554 526294 147622 526350
rect 147678 526294 165250 526350
rect 165306 526294 165374 526350
rect 165430 526294 165498 526350
rect 165554 526294 165622 526350
rect 165678 526294 183250 526350
rect 183306 526294 183374 526350
rect 183430 526294 183498 526350
rect 183554 526294 183622 526350
rect 183678 526294 201250 526350
rect 201306 526294 201374 526350
rect 201430 526294 201498 526350
rect 201554 526294 201622 526350
rect 201678 526294 219250 526350
rect 219306 526294 219374 526350
rect 219430 526294 219498 526350
rect 219554 526294 219622 526350
rect 219678 526294 237250 526350
rect 237306 526294 237374 526350
rect 237430 526294 237498 526350
rect 237554 526294 237622 526350
rect 237678 526294 255250 526350
rect 255306 526294 255374 526350
rect 255430 526294 255498 526350
rect 255554 526294 255622 526350
rect 255678 526294 273250 526350
rect 273306 526294 273374 526350
rect 273430 526294 273498 526350
rect 273554 526294 273622 526350
rect 273678 526294 291250 526350
rect 291306 526294 291374 526350
rect 291430 526294 291498 526350
rect 291554 526294 291622 526350
rect 291678 526294 309250 526350
rect 309306 526294 309374 526350
rect 309430 526294 309498 526350
rect 309554 526294 309622 526350
rect 309678 526294 327250 526350
rect 327306 526294 327374 526350
rect 327430 526294 327498 526350
rect 327554 526294 327622 526350
rect 327678 526294 345250 526350
rect 345306 526294 345374 526350
rect 345430 526294 345498 526350
rect 345554 526294 345622 526350
rect 345678 526294 363250 526350
rect 363306 526294 363374 526350
rect 363430 526294 363498 526350
rect 363554 526294 363622 526350
rect 363678 526294 381250 526350
rect 381306 526294 381374 526350
rect 381430 526294 381498 526350
rect 381554 526294 381622 526350
rect 381678 526294 399250 526350
rect 399306 526294 399374 526350
rect 399430 526294 399498 526350
rect 399554 526294 399622 526350
rect 399678 526294 417250 526350
rect 417306 526294 417374 526350
rect 417430 526294 417498 526350
rect 417554 526294 417622 526350
rect 417678 526294 435250 526350
rect 435306 526294 435374 526350
rect 435430 526294 435498 526350
rect 435554 526294 435622 526350
rect 435678 526294 453250 526350
rect 453306 526294 453374 526350
rect 453430 526294 453498 526350
rect 453554 526294 453622 526350
rect 453678 526294 471250 526350
rect 471306 526294 471374 526350
rect 471430 526294 471498 526350
rect 471554 526294 471622 526350
rect 471678 526294 489250 526350
rect 489306 526294 489374 526350
rect 489430 526294 489498 526350
rect 489554 526294 489622 526350
rect 489678 526294 507250 526350
rect 507306 526294 507374 526350
rect 507430 526294 507498 526350
rect 507554 526294 507622 526350
rect 507678 526294 525250 526350
rect 525306 526294 525374 526350
rect 525430 526294 525498 526350
rect 525554 526294 525622 526350
rect 525678 526294 543250 526350
rect 543306 526294 543374 526350
rect 543430 526294 543498 526350
rect 543554 526294 543622 526350
rect 543678 526294 561250 526350
rect 561306 526294 561374 526350
rect 561430 526294 561498 526350
rect 561554 526294 561622 526350
rect 561678 526294 579250 526350
rect 579306 526294 579374 526350
rect 579430 526294 579498 526350
rect 579554 526294 579622 526350
rect 579678 526294 596496 526350
rect 596552 526294 596620 526350
rect 596676 526294 596744 526350
rect 596800 526294 596868 526350
rect 596924 526294 597980 526350
rect -1916 526226 597980 526294
rect -1916 526170 -860 526226
rect -804 526170 -736 526226
rect -680 526170 -612 526226
rect -556 526170 -488 526226
rect -432 526170 3250 526226
rect 3306 526170 3374 526226
rect 3430 526170 3498 526226
rect 3554 526170 3622 526226
rect 3678 526170 21250 526226
rect 21306 526170 21374 526226
rect 21430 526170 21498 526226
rect 21554 526170 21622 526226
rect 21678 526170 39250 526226
rect 39306 526170 39374 526226
rect 39430 526170 39498 526226
rect 39554 526170 39622 526226
rect 39678 526170 57250 526226
rect 57306 526170 57374 526226
rect 57430 526170 57498 526226
rect 57554 526170 57622 526226
rect 57678 526170 75250 526226
rect 75306 526170 75374 526226
rect 75430 526170 75498 526226
rect 75554 526170 75622 526226
rect 75678 526170 93250 526226
rect 93306 526170 93374 526226
rect 93430 526170 93498 526226
rect 93554 526170 93622 526226
rect 93678 526170 111250 526226
rect 111306 526170 111374 526226
rect 111430 526170 111498 526226
rect 111554 526170 111622 526226
rect 111678 526170 129250 526226
rect 129306 526170 129374 526226
rect 129430 526170 129498 526226
rect 129554 526170 129622 526226
rect 129678 526170 147250 526226
rect 147306 526170 147374 526226
rect 147430 526170 147498 526226
rect 147554 526170 147622 526226
rect 147678 526170 165250 526226
rect 165306 526170 165374 526226
rect 165430 526170 165498 526226
rect 165554 526170 165622 526226
rect 165678 526170 183250 526226
rect 183306 526170 183374 526226
rect 183430 526170 183498 526226
rect 183554 526170 183622 526226
rect 183678 526170 201250 526226
rect 201306 526170 201374 526226
rect 201430 526170 201498 526226
rect 201554 526170 201622 526226
rect 201678 526170 219250 526226
rect 219306 526170 219374 526226
rect 219430 526170 219498 526226
rect 219554 526170 219622 526226
rect 219678 526170 237250 526226
rect 237306 526170 237374 526226
rect 237430 526170 237498 526226
rect 237554 526170 237622 526226
rect 237678 526170 255250 526226
rect 255306 526170 255374 526226
rect 255430 526170 255498 526226
rect 255554 526170 255622 526226
rect 255678 526170 273250 526226
rect 273306 526170 273374 526226
rect 273430 526170 273498 526226
rect 273554 526170 273622 526226
rect 273678 526170 291250 526226
rect 291306 526170 291374 526226
rect 291430 526170 291498 526226
rect 291554 526170 291622 526226
rect 291678 526170 309250 526226
rect 309306 526170 309374 526226
rect 309430 526170 309498 526226
rect 309554 526170 309622 526226
rect 309678 526170 327250 526226
rect 327306 526170 327374 526226
rect 327430 526170 327498 526226
rect 327554 526170 327622 526226
rect 327678 526170 345250 526226
rect 345306 526170 345374 526226
rect 345430 526170 345498 526226
rect 345554 526170 345622 526226
rect 345678 526170 363250 526226
rect 363306 526170 363374 526226
rect 363430 526170 363498 526226
rect 363554 526170 363622 526226
rect 363678 526170 381250 526226
rect 381306 526170 381374 526226
rect 381430 526170 381498 526226
rect 381554 526170 381622 526226
rect 381678 526170 399250 526226
rect 399306 526170 399374 526226
rect 399430 526170 399498 526226
rect 399554 526170 399622 526226
rect 399678 526170 417250 526226
rect 417306 526170 417374 526226
rect 417430 526170 417498 526226
rect 417554 526170 417622 526226
rect 417678 526170 435250 526226
rect 435306 526170 435374 526226
rect 435430 526170 435498 526226
rect 435554 526170 435622 526226
rect 435678 526170 453250 526226
rect 453306 526170 453374 526226
rect 453430 526170 453498 526226
rect 453554 526170 453622 526226
rect 453678 526170 471250 526226
rect 471306 526170 471374 526226
rect 471430 526170 471498 526226
rect 471554 526170 471622 526226
rect 471678 526170 489250 526226
rect 489306 526170 489374 526226
rect 489430 526170 489498 526226
rect 489554 526170 489622 526226
rect 489678 526170 507250 526226
rect 507306 526170 507374 526226
rect 507430 526170 507498 526226
rect 507554 526170 507622 526226
rect 507678 526170 525250 526226
rect 525306 526170 525374 526226
rect 525430 526170 525498 526226
rect 525554 526170 525622 526226
rect 525678 526170 543250 526226
rect 543306 526170 543374 526226
rect 543430 526170 543498 526226
rect 543554 526170 543622 526226
rect 543678 526170 561250 526226
rect 561306 526170 561374 526226
rect 561430 526170 561498 526226
rect 561554 526170 561622 526226
rect 561678 526170 579250 526226
rect 579306 526170 579374 526226
rect 579430 526170 579498 526226
rect 579554 526170 579622 526226
rect 579678 526170 596496 526226
rect 596552 526170 596620 526226
rect 596676 526170 596744 526226
rect 596800 526170 596868 526226
rect 596924 526170 597980 526226
rect -1916 526102 597980 526170
rect -1916 526046 -860 526102
rect -804 526046 -736 526102
rect -680 526046 -612 526102
rect -556 526046 -488 526102
rect -432 526046 3250 526102
rect 3306 526046 3374 526102
rect 3430 526046 3498 526102
rect 3554 526046 3622 526102
rect 3678 526046 21250 526102
rect 21306 526046 21374 526102
rect 21430 526046 21498 526102
rect 21554 526046 21622 526102
rect 21678 526046 39250 526102
rect 39306 526046 39374 526102
rect 39430 526046 39498 526102
rect 39554 526046 39622 526102
rect 39678 526046 57250 526102
rect 57306 526046 57374 526102
rect 57430 526046 57498 526102
rect 57554 526046 57622 526102
rect 57678 526046 75250 526102
rect 75306 526046 75374 526102
rect 75430 526046 75498 526102
rect 75554 526046 75622 526102
rect 75678 526046 93250 526102
rect 93306 526046 93374 526102
rect 93430 526046 93498 526102
rect 93554 526046 93622 526102
rect 93678 526046 111250 526102
rect 111306 526046 111374 526102
rect 111430 526046 111498 526102
rect 111554 526046 111622 526102
rect 111678 526046 129250 526102
rect 129306 526046 129374 526102
rect 129430 526046 129498 526102
rect 129554 526046 129622 526102
rect 129678 526046 147250 526102
rect 147306 526046 147374 526102
rect 147430 526046 147498 526102
rect 147554 526046 147622 526102
rect 147678 526046 165250 526102
rect 165306 526046 165374 526102
rect 165430 526046 165498 526102
rect 165554 526046 165622 526102
rect 165678 526046 183250 526102
rect 183306 526046 183374 526102
rect 183430 526046 183498 526102
rect 183554 526046 183622 526102
rect 183678 526046 201250 526102
rect 201306 526046 201374 526102
rect 201430 526046 201498 526102
rect 201554 526046 201622 526102
rect 201678 526046 219250 526102
rect 219306 526046 219374 526102
rect 219430 526046 219498 526102
rect 219554 526046 219622 526102
rect 219678 526046 237250 526102
rect 237306 526046 237374 526102
rect 237430 526046 237498 526102
rect 237554 526046 237622 526102
rect 237678 526046 255250 526102
rect 255306 526046 255374 526102
rect 255430 526046 255498 526102
rect 255554 526046 255622 526102
rect 255678 526046 273250 526102
rect 273306 526046 273374 526102
rect 273430 526046 273498 526102
rect 273554 526046 273622 526102
rect 273678 526046 291250 526102
rect 291306 526046 291374 526102
rect 291430 526046 291498 526102
rect 291554 526046 291622 526102
rect 291678 526046 309250 526102
rect 309306 526046 309374 526102
rect 309430 526046 309498 526102
rect 309554 526046 309622 526102
rect 309678 526046 327250 526102
rect 327306 526046 327374 526102
rect 327430 526046 327498 526102
rect 327554 526046 327622 526102
rect 327678 526046 345250 526102
rect 345306 526046 345374 526102
rect 345430 526046 345498 526102
rect 345554 526046 345622 526102
rect 345678 526046 363250 526102
rect 363306 526046 363374 526102
rect 363430 526046 363498 526102
rect 363554 526046 363622 526102
rect 363678 526046 381250 526102
rect 381306 526046 381374 526102
rect 381430 526046 381498 526102
rect 381554 526046 381622 526102
rect 381678 526046 399250 526102
rect 399306 526046 399374 526102
rect 399430 526046 399498 526102
rect 399554 526046 399622 526102
rect 399678 526046 417250 526102
rect 417306 526046 417374 526102
rect 417430 526046 417498 526102
rect 417554 526046 417622 526102
rect 417678 526046 435250 526102
rect 435306 526046 435374 526102
rect 435430 526046 435498 526102
rect 435554 526046 435622 526102
rect 435678 526046 453250 526102
rect 453306 526046 453374 526102
rect 453430 526046 453498 526102
rect 453554 526046 453622 526102
rect 453678 526046 471250 526102
rect 471306 526046 471374 526102
rect 471430 526046 471498 526102
rect 471554 526046 471622 526102
rect 471678 526046 489250 526102
rect 489306 526046 489374 526102
rect 489430 526046 489498 526102
rect 489554 526046 489622 526102
rect 489678 526046 507250 526102
rect 507306 526046 507374 526102
rect 507430 526046 507498 526102
rect 507554 526046 507622 526102
rect 507678 526046 525250 526102
rect 525306 526046 525374 526102
rect 525430 526046 525498 526102
rect 525554 526046 525622 526102
rect 525678 526046 543250 526102
rect 543306 526046 543374 526102
rect 543430 526046 543498 526102
rect 543554 526046 543622 526102
rect 543678 526046 561250 526102
rect 561306 526046 561374 526102
rect 561430 526046 561498 526102
rect 561554 526046 561622 526102
rect 561678 526046 579250 526102
rect 579306 526046 579374 526102
rect 579430 526046 579498 526102
rect 579554 526046 579622 526102
rect 579678 526046 596496 526102
rect 596552 526046 596620 526102
rect 596676 526046 596744 526102
rect 596800 526046 596868 526102
rect 596924 526046 597980 526102
rect -1916 525978 597980 526046
rect -1916 525922 -860 525978
rect -804 525922 -736 525978
rect -680 525922 -612 525978
rect -556 525922 -488 525978
rect -432 525922 3250 525978
rect 3306 525922 3374 525978
rect 3430 525922 3498 525978
rect 3554 525922 3622 525978
rect 3678 525922 21250 525978
rect 21306 525922 21374 525978
rect 21430 525922 21498 525978
rect 21554 525922 21622 525978
rect 21678 525922 39250 525978
rect 39306 525922 39374 525978
rect 39430 525922 39498 525978
rect 39554 525922 39622 525978
rect 39678 525922 57250 525978
rect 57306 525922 57374 525978
rect 57430 525922 57498 525978
rect 57554 525922 57622 525978
rect 57678 525922 75250 525978
rect 75306 525922 75374 525978
rect 75430 525922 75498 525978
rect 75554 525922 75622 525978
rect 75678 525922 93250 525978
rect 93306 525922 93374 525978
rect 93430 525922 93498 525978
rect 93554 525922 93622 525978
rect 93678 525922 111250 525978
rect 111306 525922 111374 525978
rect 111430 525922 111498 525978
rect 111554 525922 111622 525978
rect 111678 525922 129250 525978
rect 129306 525922 129374 525978
rect 129430 525922 129498 525978
rect 129554 525922 129622 525978
rect 129678 525922 147250 525978
rect 147306 525922 147374 525978
rect 147430 525922 147498 525978
rect 147554 525922 147622 525978
rect 147678 525922 165250 525978
rect 165306 525922 165374 525978
rect 165430 525922 165498 525978
rect 165554 525922 165622 525978
rect 165678 525922 183250 525978
rect 183306 525922 183374 525978
rect 183430 525922 183498 525978
rect 183554 525922 183622 525978
rect 183678 525922 201250 525978
rect 201306 525922 201374 525978
rect 201430 525922 201498 525978
rect 201554 525922 201622 525978
rect 201678 525922 219250 525978
rect 219306 525922 219374 525978
rect 219430 525922 219498 525978
rect 219554 525922 219622 525978
rect 219678 525922 237250 525978
rect 237306 525922 237374 525978
rect 237430 525922 237498 525978
rect 237554 525922 237622 525978
rect 237678 525922 255250 525978
rect 255306 525922 255374 525978
rect 255430 525922 255498 525978
rect 255554 525922 255622 525978
rect 255678 525922 273250 525978
rect 273306 525922 273374 525978
rect 273430 525922 273498 525978
rect 273554 525922 273622 525978
rect 273678 525922 291250 525978
rect 291306 525922 291374 525978
rect 291430 525922 291498 525978
rect 291554 525922 291622 525978
rect 291678 525922 309250 525978
rect 309306 525922 309374 525978
rect 309430 525922 309498 525978
rect 309554 525922 309622 525978
rect 309678 525922 327250 525978
rect 327306 525922 327374 525978
rect 327430 525922 327498 525978
rect 327554 525922 327622 525978
rect 327678 525922 345250 525978
rect 345306 525922 345374 525978
rect 345430 525922 345498 525978
rect 345554 525922 345622 525978
rect 345678 525922 363250 525978
rect 363306 525922 363374 525978
rect 363430 525922 363498 525978
rect 363554 525922 363622 525978
rect 363678 525922 381250 525978
rect 381306 525922 381374 525978
rect 381430 525922 381498 525978
rect 381554 525922 381622 525978
rect 381678 525922 399250 525978
rect 399306 525922 399374 525978
rect 399430 525922 399498 525978
rect 399554 525922 399622 525978
rect 399678 525922 417250 525978
rect 417306 525922 417374 525978
rect 417430 525922 417498 525978
rect 417554 525922 417622 525978
rect 417678 525922 435250 525978
rect 435306 525922 435374 525978
rect 435430 525922 435498 525978
rect 435554 525922 435622 525978
rect 435678 525922 453250 525978
rect 453306 525922 453374 525978
rect 453430 525922 453498 525978
rect 453554 525922 453622 525978
rect 453678 525922 471250 525978
rect 471306 525922 471374 525978
rect 471430 525922 471498 525978
rect 471554 525922 471622 525978
rect 471678 525922 489250 525978
rect 489306 525922 489374 525978
rect 489430 525922 489498 525978
rect 489554 525922 489622 525978
rect 489678 525922 507250 525978
rect 507306 525922 507374 525978
rect 507430 525922 507498 525978
rect 507554 525922 507622 525978
rect 507678 525922 525250 525978
rect 525306 525922 525374 525978
rect 525430 525922 525498 525978
rect 525554 525922 525622 525978
rect 525678 525922 543250 525978
rect 543306 525922 543374 525978
rect 543430 525922 543498 525978
rect 543554 525922 543622 525978
rect 543678 525922 561250 525978
rect 561306 525922 561374 525978
rect 561430 525922 561498 525978
rect 561554 525922 561622 525978
rect 561678 525922 579250 525978
rect 579306 525922 579374 525978
rect 579430 525922 579498 525978
rect 579554 525922 579622 525978
rect 579678 525922 596496 525978
rect 596552 525922 596620 525978
rect 596676 525922 596744 525978
rect 596800 525922 596868 525978
rect 596924 525922 597980 525978
rect -1916 525826 597980 525922
rect -1916 514350 597980 514446
rect -1916 514294 -1820 514350
rect -1764 514294 -1696 514350
rect -1640 514294 -1572 514350
rect -1516 514294 -1448 514350
rect -1392 514294 6970 514350
rect 7026 514294 7094 514350
rect 7150 514294 7218 514350
rect 7274 514294 7342 514350
rect 7398 514294 24970 514350
rect 25026 514294 25094 514350
rect 25150 514294 25218 514350
rect 25274 514294 25342 514350
rect 25398 514294 42970 514350
rect 43026 514294 43094 514350
rect 43150 514294 43218 514350
rect 43274 514294 43342 514350
rect 43398 514294 60970 514350
rect 61026 514294 61094 514350
rect 61150 514294 61218 514350
rect 61274 514294 61342 514350
rect 61398 514294 78970 514350
rect 79026 514294 79094 514350
rect 79150 514294 79218 514350
rect 79274 514294 79342 514350
rect 79398 514294 96970 514350
rect 97026 514294 97094 514350
rect 97150 514294 97218 514350
rect 97274 514294 97342 514350
rect 97398 514294 114970 514350
rect 115026 514294 115094 514350
rect 115150 514294 115218 514350
rect 115274 514294 115342 514350
rect 115398 514294 132970 514350
rect 133026 514294 133094 514350
rect 133150 514294 133218 514350
rect 133274 514294 133342 514350
rect 133398 514294 150970 514350
rect 151026 514294 151094 514350
rect 151150 514294 151218 514350
rect 151274 514294 151342 514350
rect 151398 514294 168970 514350
rect 169026 514294 169094 514350
rect 169150 514294 169218 514350
rect 169274 514294 169342 514350
rect 169398 514294 186970 514350
rect 187026 514294 187094 514350
rect 187150 514294 187218 514350
rect 187274 514294 187342 514350
rect 187398 514294 204970 514350
rect 205026 514294 205094 514350
rect 205150 514294 205218 514350
rect 205274 514294 205342 514350
rect 205398 514294 222970 514350
rect 223026 514294 223094 514350
rect 223150 514294 223218 514350
rect 223274 514294 223342 514350
rect 223398 514294 240970 514350
rect 241026 514294 241094 514350
rect 241150 514294 241218 514350
rect 241274 514294 241342 514350
rect 241398 514294 258970 514350
rect 259026 514294 259094 514350
rect 259150 514294 259218 514350
rect 259274 514294 259342 514350
rect 259398 514294 276970 514350
rect 277026 514294 277094 514350
rect 277150 514294 277218 514350
rect 277274 514294 277342 514350
rect 277398 514294 294970 514350
rect 295026 514294 295094 514350
rect 295150 514294 295218 514350
rect 295274 514294 295342 514350
rect 295398 514294 312970 514350
rect 313026 514294 313094 514350
rect 313150 514294 313218 514350
rect 313274 514294 313342 514350
rect 313398 514294 330970 514350
rect 331026 514294 331094 514350
rect 331150 514294 331218 514350
rect 331274 514294 331342 514350
rect 331398 514294 348970 514350
rect 349026 514294 349094 514350
rect 349150 514294 349218 514350
rect 349274 514294 349342 514350
rect 349398 514294 366970 514350
rect 367026 514294 367094 514350
rect 367150 514294 367218 514350
rect 367274 514294 367342 514350
rect 367398 514294 384970 514350
rect 385026 514294 385094 514350
rect 385150 514294 385218 514350
rect 385274 514294 385342 514350
rect 385398 514294 402970 514350
rect 403026 514294 403094 514350
rect 403150 514294 403218 514350
rect 403274 514294 403342 514350
rect 403398 514294 420970 514350
rect 421026 514294 421094 514350
rect 421150 514294 421218 514350
rect 421274 514294 421342 514350
rect 421398 514294 438970 514350
rect 439026 514294 439094 514350
rect 439150 514294 439218 514350
rect 439274 514294 439342 514350
rect 439398 514294 456970 514350
rect 457026 514294 457094 514350
rect 457150 514294 457218 514350
rect 457274 514294 457342 514350
rect 457398 514294 474970 514350
rect 475026 514294 475094 514350
rect 475150 514294 475218 514350
rect 475274 514294 475342 514350
rect 475398 514294 492970 514350
rect 493026 514294 493094 514350
rect 493150 514294 493218 514350
rect 493274 514294 493342 514350
rect 493398 514294 510970 514350
rect 511026 514294 511094 514350
rect 511150 514294 511218 514350
rect 511274 514294 511342 514350
rect 511398 514294 528970 514350
rect 529026 514294 529094 514350
rect 529150 514294 529218 514350
rect 529274 514294 529342 514350
rect 529398 514294 546970 514350
rect 547026 514294 547094 514350
rect 547150 514294 547218 514350
rect 547274 514294 547342 514350
rect 547398 514294 564970 514350
rect 565026 514294 565094 514350
rect 565150 514294 565218 514350
rect 565274 514294 565342 514350
rect 565398 514294 582970 514350
rect 583026 514294 583094 514350
rect 583150 514294 583218 514350
rect 583274 514294 583342 514350
rect 583398 514294 597456 514350
rect 597512 514294 597580 514350
rect 597636 514294 597704 514350
rect 597760 514294 597828 514350
rect 597884 514294 597980 514350
rect -1916 514226 597980 514294
rect -1916 514170 -1820 514226
rect -1764 514170 -1696 514226
rect -1640 514170 -1572 514226
rect -1516 514170 -1448 514226
rect -1392 514170 6970 514226
rect 7026 514170 7094 514226
rect 7150 514170 7218 514226
rect 7274 514170 7342 514226
rect 7398 514170 24970 514226
rect 25026 514170 25094 514226
rect 25150 514170 25218 514226
rect 25274 514170 25342 514226
rect 25398 514170 42970 514226
rect 43026 514170 43094 514226
rect 43150 514170 43218 514226
rect 43274 514170 43342 514226
rect 43398 514170 60970 514226
rect 61026 514170 61094 514226
rect 61150 514170 61218 514226
rect 61274 514170 61342 514226
rect 61398 514170 78970 514226
rect 79026 514170 79094 514226
rect 79150 514170 79218 514226
rect 79274 514170 79342 514226
rect 79398 514170 96970 514226
rect 97026 514170 97094 514226
rect 97150 514170 97218 514226
rect 97274 514170 97342 514226
rect 97398 514170 114970 514226
rect 115026 514170 115094 514226
rect 115150 514170 115218 514226
rect 115274 514170 115342 514226
rect 115398 514170 132970 514226
rect 133026 514170 133094 514226
rect 133150 514170 133218 514226
rect 133274 514170 133342 514226
rect 133398 514170 150970 514226
rect 151026 514170 151094 514226
rect 151150 514170 151218 514226
rect 151274 514170 151342 514226
rect 151398 514170 168970 514226
rect 169026 514170 169094 514226
rect 169150 514170 169218 514226
rect 169274 514170 169342 514226
rect 169398 514170 186970 514226
rect 187026 514170 187094 514226
rect 187150 514170 187218 514226
rect 187274 514170 187342 514226
rect 187398 514170 204970 514226
rect 205026 514170 205094 514226
rect 205150 514170 205218 514226
rect 205274 514170 205342 514226
rect 205398 514170 222970 514226
rect 223026 514170 223094 514226
rect 223150 514170 223218 514226
rect 223274 514170 223342 514226
rect 223398 514170 240970 514226
rect 241026 514170 241094 514226
rect 241150 514170 241218 514226
rect 241274 514170 241342 514226
rect 241398 514170 258970 514226
rect 259026 514170 259094 514226
rect 259150 514170 259218 514226
rect 259274 514170 259342 514226
rect 259398 514170 276970 514226
rect 277026 514170 277094 514226
rect 277150 514170 277218 514226
rect 277274 514170 277342 514226
rect 277398 514170 294970 514226
rect 295026 514170 295094 514226
rect 295150 514170 295218 514226
rect 295274 514170 295342 514226
rect 295398 514170 312970 514226
rect 313026 514170 313094 514226
rect 313150 514170 313218 514226
rect 313274 514170 313342 514226
rect 313398 514170 330970 514226
rect 331026 514170 331094 514226
rect 331150 514170 331218 514226
rect 331274 514170 331342 514226
rect 331398 514170 348970 514226
rect 349026 514170 349094 514226
rect 349150 514170 349218 514226
rect 349274 514170 349342 514226
rect 349398 514170 366970 514226
rect 367026 514170 367094 514226
rect 367150 514170 367218 514226
rect 367274 514170 367342 514226
rect 367398 514170 384970 514226
rect 385026 514170 385094 514226
rect 385150 514170 385218 514226
rect 385274 514170 385342 514226
rect 385398 514170 402970 514226
rect 403026 514170 403094 514226
rect 403150 514170 403218 514226
rect 403274 514170 403342 514226
rect 403398 514170 420970 514226
rect 421026 514170 421094 514226
rect 421150 514170 421218 514226
rect 421274 514170 421342 514226
rect 421398 514170 438970 514226
rect 439026 514170 439094 514226
rect 439150 514170 439218 514226
rect 439274 514170 439342 514226
rect 439398 514170 456970 514226
rect 457026 514170 457094 514226
rect 457150 514170 457218 514226
rect 457274 514170 457342 514226
rect 457398 514170 474970 514226
rect 475026 514170 475094 514226
rect 475150 514170 475218 514226
rect 475274 514170 475342 514226
rect 475398 514170 492970 514226
rect 493026 514170 493094 514226
rect 493150 514170 493218 514226
rect 493274 514170 493342 514226
rect 493398 514170 510970 514226
rect 511026 514170 511094 514226
rect 511150 514170 511218 514226
rect 511274 514170 511342 514226
rect 511398 514170 528970 514226
rect 529026 514170 529094 514226
rect 529150 514170 529218 514226
rect 529274 514170 529342 514226
rect 529398 514170 546970 514226
rect 547026 514170 547094 514226
rect 547150 514170 547218 514226
rect 547274 514170 547342 514226
rect 547398 514170 564970 514226
rect 565026 514170 565094 514226
rect 565150 514170 565218 514226
rect 565274 514170 565342 514226
rect 565398 514170 582970 514226
rect 583026 514170 583094 514226
rect 583150 514170 583218 514226
rect 583274 514170 583342 514226
rect 583398 514170 597456 514226
rect 597512 514170 597580 514226
rect 597636 514170 597704 514226
rect 597760 514170 597828 514226
rect 597884 514170 597980 514226
rect -1916 514102 597980 514170
rect -1916 514046 -1820 514102
rect -1764 514046 -1696 514102
rect -1640 514046 -1572 514102
rect -1516 514046 -1448 514102
rect -1392 514046 6970 514102
rect 7026 514046 7094 514102
rect 7150 514046 7218 514102
rect 7274 514046 7342 514102
rect 7398 514046 24970 514102
rect 25026 514046 25094 514102
rect 25150 514046 25218 514102
rect 25274 514046 25342 514102
rect 25398 514046 42970 514102
rect 43026 514046 43094 514102
rect 43150 514046 43218 514102
rect 43274 514046 43342 514102
rect 43398 514046 60970 514102
rect 61026 514046 61094 514102
rect 61150 514046 61218 514102
rect 61274 514046 61342 514102
rect 61398 514046 78970 514102
rect 79026 514046 79094 514102
rect 79150 514046 79218 514102
rect 79274 514046 79342 514102
rect 79398 514046 96970 514102
rect 97026 514046 97094 514102
rect 97150 514046 97218 514102
rect 97274 514046 97342 514102
rect 97398 514046 114970 514102
rect 115026 514046 115094 514102
rect 115150 514046 115218 514102
rect 115274 514046 115342 514102
rect 115398 514046 132970 514102
rect 133026 514046 133094 514102
rect 133150 514046 133218 514102
rect 133274 514046 133342 514102
rect 133398 514046 150970 514102
rect 151026 514046 151094 514102
rect 151150 514046 151218 514102
rect 151274 514046 151342 514102
rect 151398 514046 168970 514102
rect 169026 514046 169094 514102
rect 169150 514046 169218 514102
rect 169274 514046 169342 514102
rect 169398 514046 186970 514102
rect 187026 514046 187094 514102
rect 187150 514046 187218 514102
rect 187274 514046 187342 514102
rect 187398 514046 204970 514102
rect 205026 514046 205094 514102
rect 205150 514046 205218 514102
rect 205274 514046 205342 514102
rect 205398 514046 222970 514102
rect 223026 514046 223094 514102
rect 223150 514046 223218 514102
rect 223274 514046 223342 514102
rect 223398 514046 240970 514102
rect 241026 514046 241094 514102
rect 241150 514046 241218 514102
rect 241274 514046 241342 514102
rect 241398 514046 258970 514102
rect 259026 514046 259094 514102
rect 259150 514046 259218 514102
rect 259274 514046 259342 514102
rect 259398 514046 276970 514102
rect 277026 514046 277094 514102
rect 277150 514046 277218 514102
rect 277274 514046 277342 514102
rect 277398 514046 294970 514102
rect 295026 514046 295094 514102
rect 295150 514046 295218 514102
rect 295274 514046 295342 514102
rect 295398 514046 312970 514102
rect 313026 514046 313094 514102
rect 313150 514046 313218 514102
rect 313274 514046 313342 514102
rect 313398 514046 330970 514102
rect 331026 514046 331094 514102
rect 331150 514046 331218 514102
rect 331274 514046 331342 514102
rect 331398 514046 348970 514102
rect 349026 514046 349094 514102
rect 349150 514046 349218 514102
rect 349274 514046 349342 514102
rect 349398 514046 366970 514102
rect 367026 514046 367094 514102
rect 367150 514046 367218 514102
rect 367274 514046 367342 514102
rect 367398 514046 384970 514102
rect 385026 514046 385094 514102
rect 385150 514046 385218 514102
rect 385274 514046 385342 514102
rect 385398 514046 402970 514102
rect 403026 514046 403094 514102
rect 403150 514046 403218 514102
rect 403274 514046 403342 514102
rect 403398 514046 420970 514102
rect 421026 514046 421094 514102
rect 421150 514046 421218 514102
rect 421274 514046 421342 514102
rect 421398 514046 438970 514102
rect 439026 514046 439094 514102
rect 439150 514046 439218 514102
rect 439274 514046 439342 514102
rect 439398 514046 456970 514102
rect 457026 514046 457094 514102
rect 457150 514046 457218 514102
rect 457274 514046 457342 514102
rect 457398 514046 474970 514102
rect 475026 514046 475094 514102
rect 475150 514046 475218 514102
rect 475274 514046 475342 514102
rect 475398 514046 492970 514102
rect 493026 514046 493094 514102
rect 493150 514046 493218 514102
rect 493274 514046 493342 514102
rect 493398 514046 510970 514102
rect 511026 514046 511094 514102
rect 511150 514046 511218 514102
rect 511274 514046 511342 514102
rect 511398 514046 528970 514102
rect 529026 514046 529094 514102
rect 529150 514046 529218 514102
rect 529274 514046 529342 514102
rect 529398 514046 546970 514102
rect 547026 514046 547094 514102
rect 547150 514046 547218 514102
rect 547274 514046 547342 514102
rect 547398 514046 564970 514102
rect 565026 514046 565094 514102
rect 565150 514046 565218 514102
rect 565274 514046 565342 514102
rect 565398 514046 582970 514102
rect 583026 514046 583094 514102
rect 583150 514046 583218 514102
rect 583274 514046 583342 514102
rect 583398 514046 597456 514102
rect 597512 514046 597580 514102
rect 597636 514046 597704 514102
rect 597760 514046 597828 514102
rect 597884 514046 597980 514102
rect -1916 513978 597980 514046
rect -1916 513922 -1820 513978
rect -1764 513922 -1696 513978
rect -1640 513922 -1572 513978
rect -1516 513922 -1448 513978
rect -1392 513922 6970 513978
rect 7026 513922 7094 513978
rect 7150 513922 7218 513978
rect 7274 513922 7342 513978
rect 7398 513922 24970 513978
rect 25026 513922 25094 513978
rect 25150 513922 25218 513978
rect 25274 513922 25342 513978
rect 25398 513922 42970 513978
rect 43026 513922 43094 513978
rect 43150 513922 43218 513978
rect 43274 513922 43342 513978
rect 43398 513922 60970 513978
rect 61026 513922 61094 513978
rect 61150 513922 61218 513978
rect 61274 513922 61342 513978
rect 61398 513922 78970 513978
rect 79026 513922 79094 513978
rect 79150 513922 79218 513978
rect 79274 513922 79342 513978
rect 79398 513922 96970 513978
rect 97026 513922 97094 513978
rect 97150 513922 97218 513978
rect 97274 513922 97342 513978
rect 97398 513922 114970 513978
rect 115026 513922 115094 513978
rect 115150 513922 115218 513978
rect 115274 513922 115342 513978
rect 115398 513922 132970 513978
rect 133026 513922 133094 513978
rect 133150 513922 133218 513978
rect 133274 513922 133342 513978
rect 133398 513922 150970 513978
rect 151026 513922 151094 513978
rect 151150 513922 151218 513978
rect 151274 513922 151342 513978
rect 151398 513922 168970 513978
rect 169026 513922 169094 513978
rect 169150 513922 169218 513978
rect 169274 513922 169342 513978
rect 169398 513922 186970 513978
rect 187026 513922 187094 513978
rect 187150 513922 187218 513978
rect 187274 513922 187342 513978
rect 187398 513922 204970 513978
rect 205026 513922 205094 513978
rect 205150 513922 205218 513978
rect 205274 513922 205342 513978
rect 205398 513922 222970 513978
rect 223026 513922 223094 513978
rect 223150 513922 223218 513978
rect 223274 513922 223342 513978
rect 223398 513922 240970 513978
rect 241026 513922 241094 513978
rect 241150 513922 241218 513978
rect 241274 513922 241342 513978
rect 241398 513922 258970 513978
rect 259026 513922 259094 513978
rect 259150 513922 259218 513978
rect 259274 513922 259342 513978
rect 259398 513922 276970 513978
rect 277026 513922 277094 513978
rect 277150 513922 277218 513978
rect 277274 513922 277342 513978
rect 277398 513922 294970 513978
rect 295026 513922 295094 513978
rect 295150 513922 295218 513978
rect 295274 513922 295342 513978
rect 295398 513922 312970 513978
rect 313026 513922 313094 513978
rect 313150 513922 313218 513978
rect 313274 513922 313342 513978
rect 313398 513922 330970 513978
rect 331026 513922 331094 513978
rect 331150 513922 331218 513978
rect 331274 513922 331342 513978
rect 331398 513922 348970 513978
rect 349026 513922 349094 513978
rect 349150 513922 349218 513978
rect 349274 513922 349342 513978
rect 349398 513922 366970 513978
rect 367026 513922 367094 513978
rect 367150 513922 367218 513978
rect 367274 513922 367342 513978
rect 367398 513922 384970 513978
rect 385026 513922 385094 513978
rect 385150 513922 385218 513978
rect 385274 513922 385342 513978
rect 385398 513922 402970 513978
rect 403026 513922 403094 513978
rect 403150 513922 403218 513978
rect 403274 513922 403342 513978
rect 403398 513922 420970 513978
rect 421026 513922 421094 513978
rect 421150 513922 421218 513978
rect 421274 513922 421342 513978
rect 421398 513922 438970 513978
rect 439026 513922 439094 513978
rect 439150 513922 439218 513978
rect 439274 513922 439342 513978
rect 439398 513922 456970 513978
rect 457026 513922 457094 513978
rect 457150 513922 457218 513978
rect 457274 513922 457342 513978
rect 457398 513922 474970 513978
rect 475026 513922 475094 513978
rect 475150 513922 475218 513978
rect 475274 513922 475342 513978
rect 475398 513922 492970 513978
rect 493026 513922 493094 513978
rect 493150 513922 493218 513978
rect 493274 513922 493342 513978
rect 493398 513922 510970 513978
rect 511026 513922 511094 513978
rect 511150 513922 511218 513978
rect 511274 513922 511342 513978
rect 511398 513922 528970 513978
rect 529026 513922 529094 513978
rect 529150 513922 529218 513978
rect 529274 513922 529342 513978
rect 529398 513922 546970 513978
rect 547026 513922 547094 513978
rect 547150 513922 547218 513978
rect 547274 513922 547342 513978
rect 547398 513922 564970 513978
rect 565026 513922 565094 513978
rect 565150 513922 565218 513978
rect 565274 513922 565342 513978
rect 565398 513922 582970 513978
rect 583026 513922 583094 513978
rect 583150 513922 583218 513978
rect 583274 513922 583342 513978
rect 583398 513922 597456 513978
rect 597512 513922 597580 513978
rect 597636 513922 597704 513978
rect 597760 513922 597828 513978
rect 597884 513922 597980 513978
rect -1916 513826 597980 513922
rect -1916 508350 597980 508446
rect -1916 508294 -860 508350
rect -804 508294 -736 508350
rect -680 508294 -612 508350
rect -556 508294 -488 508350
rect -432 508294 3250 508350
rect 3306 508294 3374 508350
rect 3430 508294 3498 508350
rect 3554 508294 3622 508350
rect 3678 508294 21250 508350
rect 21306 508294 21374 508350
rect 21430 508294 21498 508350
rect 21554 508294 21622 508350
rect 21678 508294 39250 508350
rect 39306 508294 39374 508350
rect 39430 508294 39498 508350
rect 39554 508294 39622 508350
rect 39678 508294 57250 508350
rect 57306 508294 57374 508350
rect 57430 508294 57498 508350
rect 57554 508294 57622 508350
rect 57678 508294 75250 508350
rect 75306 508294 75374 508350
rect 75430 508294 75498 508350
rect 75554 508294 75622 508350
rect 75678 508294 93250 508350
rect 93306 508294 93374 508350
rect 93430 508294 93498 508350
rect 93554 508294 93622 508350
rect 93678 508294 111250 508350
rect 111306 508294 111374 508350
rect 111430 508294 111498 508350
rect 111554 508294 111622 508350
rect 111678 508294 129250 508350
rect 129306 508294 129374 508350
rect 129430 508294 129498 508350
rect 129554 508294 129622 508350
rect 129678 508294 147250 508350
rect 147306 508294 147374 508350
rect 147430 508294 147498 508350
rect 147554 508294 147622 508350
rect 147678 508294 165250 508350
rect 165306 508294 165374 508350
rect 165430 508294 165498 508350
rect 165554 508294 165622 508350
rect 165678 508294 183250 508350
rect 183306 508294 183374 508350
rect 183430 508294 183498 508350
rect 183554 508294 183622 508350
rect 183678 508294 201250 508350
rect 201306 508294 201374 508350
rect 201430 508294 201498 508350
rect 201554 508294 201622 508350
rect 201678 508294 219250 508350
rect 219306 508294 219374 508350
rect 219430 508294 219498 508350
rect 219554 508294 219622 508350
rect 219678 508294 237250 508350
rect 237306 508294 237374 508350
rect 237430 508294 237498 508350
rect 237554 508294 237622 508350
rect 237678 508294 255250 508350
rect 255306 508294 255374 508350
rect 255430 508294 255498 508350
rect 255554 508294 255622 508350
rect 255678 508294 273250 508350
rect 273306 508294 273374 508350
rect 273430 508294 273498 508350
rect 273554 508294 273622 508350
rect 273678 508294 291250 508350
rect 291306 508294 291374 508350
rect 291430 508294 291498 508350
rect 291554 508294 291622 508350
rect 291678 508294 309250 508350
rect 309306 508294 309374 508350
rect 309430 508294 309498 508350
rect 309554 508294 309622 508350
rect 309678 508294 327250 508350
rect 327306 508294 327374 508350
rect 327430 508294 327498 508350
rect 327554 508294 327622 508350
rect 327678 508294 345250 508350
rect 345306 508294 345374 508350
rect 345430 508294 345498 508350
rect 345554 508294 345622 508350
rect 345678 508294 363250 508350
rect 363306 508294 363374 508350
rect 363430 508294 363498 508350
rect 363554 508294 363622 508350
rect 363678 508294 381250 508350
rect 381306 508294 381374 508350
rect 381430 508294 381498 508350
rect 381554 508294 381622 508350
rect 381678 508294 399250 508350
rect 399306 508294 399374 508350
rect 399430 508294 399498 508350
rect 399554 508294 399622 508350
rect 399678 508294 417250 508350
rect 417306 508294 417374 508350
rect 417430 508294 417498 508350
rect 417554 508294 417622 508350
rect 417678 508294 435250 508350
rect 435306 508294 435374 508350
rect 435430 508294 435498 508350
rect 435554 508294 435622 508350
rect 435678 508294 453250 508350
rect 453306 508294 453374 508350
rect 453430 508294 453498 508350
rect 453554 508294 453622 508350
rect 453678 508294 471250 508350
rect 471306 508294 471374 508350
rect 471430 508294 471498 508350
rect 471554 508294 471622 508350
rect 471678 508294 489250 508350
rect 489306 508294 489374 508350
rect 489430 508294 489498 508350
rect 489554 508294 489622 508350
rect 489678 508294 507250 508350
rect 507306 508294 507374 508350
rect 507430 508294 507498 508350
rect 507554 508294 507622 508350
rect 507678 508294 525250 508350
rect 525306 508294 525374 508350
rect 525430 508294 525498 508350
rect 525554 508294 525622 508350
rect 525678 508294 543250 508350
rect 543306 508294 543374 508350
rect 543430 508294 543498 508350
rect 543554 508294 543622 508350
rect 543678 508294 561250 508350
rect 561306 508294 561374 508350
rect 561430 508294 561498 508350
rect 561554 508294 561622 508350
rect 561678 508294 579250 508350
rect 579306 508294 579374 508350
rect 579430 508294 579498 508350
rect 579554 508294 579622 508350
rect 579678 508294 596496 508350
rect 596552 508294 596620 508350
rect 596676 508294 596744 508350
rect 596800 508294 596868 508350
rect 596924 508294 597980 508350
rect -1916 508226 597980 508294
rect -1916 508170 -860 508226
rect -804 508170 -736 508226
rect -680 508170 -612 508226
rect -556 508170 -488 508226
rect -432 508170 3250 508226
rect 3306 508170 3374 508226
rect 3430 508170 3498 508226
rect 3554 508170 3622 508226
rect 3678 508170 21250 508226
rect 21306 508170 21374 508226
rect 21430 508170 21498 508226
rect 21554 508170 21622 508226
rect 21678 508170 39250 508226
rect 39306 508170 39374 508226
rect 39430 508170 39498 508226
rect 39554 508170 39622 508226
rect 39678 508170 57250 508226
rect 57306 508170 57374 508226
rect 57430 508170 57498 508226
rect 57554 508170 57622 508226
rect 57678 508170 75250 508226
rect 75306 508170 75374 508226
rect 75430 508170 75498 508226
rect 75554 508170 75622 508226
rect 75678 508170 93250 508226
rect 93306 508170 93374 508226
rect 93430 508170 93498 508226
rect 93554 508170 93622 508226
rect 93678 508170 111250 508226
rect 111306 508170 111374 508226
rect 111430 508170 111498 508226
rect 111554 508170 111622 508226
rect 111678 508170 129250 508226
rect 129306 508170 129374 508226
rect 129430 508170 129498 508226
rect 129554 508170 129622 508226
rect 129678 508170 147250 508226
rect 147306 508170 147374 508226
rect 147430 508170 147498 508226
rect 147554 508170 147622 508226
rect 147678 508170 165250 508226
rect 165306 508170 165374 508226
rect 165430 508170 165498 508226
rect 165554 508170 165622 508226
rect 165678 508170 183250 508226
rect 183306 508170 183374 508226
rect 183430 508170 183498 508226
rect 183554 508170 183622 508226
rect 183678 508170 201250 508226
rect 201306 508170 201374 508226
rect 201430 508170 201498 508226
rect 201554 508170 201622 508226
rect 201678 508170 219250 508226
rect 219306 508170 219374 508226
rect 219430 508170 219498 508226
rect 219554 508170 219622 508226
rect 219678 508170 237250 508226
rect 237306 508170 237374 508226
rect 237430 508170 237498 508226
rect 237554 508170 237622 508226
rect 237678 508170 255250 508226
rect 255306 508170 255374 508226
rect 255430 508170 255498 508226
rect 255554 508170 255622 508226
rect 255678 508170 273250 508226
rect 273306 508170 273374 508226
rect 273430 508170 273498 508226
rect 273554 508170 273622 508226
rect 273678 508170 291250 508226
rect 291306 508170 291374 508226
rect 291430 508170 291498 508226
rect 291554 508170 291622 508226
rect 291678 508170 309250 508226
rect 309306 508170 309374 508226
rect 309430 508170 309498 508226
rect 309554 508170 309622 508226
rect 309678 508170 327250 508226
rect 327306 508170 327374 508226
rect 327430 508170 327498 508226
rect 327554 508170 327622 508226
rect 327678 508170 345250 508226
rect 345306 508170 345374 508226
rect 345430 508170 345498 508226
rect 345554 508170 345622 508226
rect 345678 508170 363250 508226
rect 363306 508170 363374 508226
rect 363430 508170 363498 508226
rect 363554 508170 363622 508226
rect 363678 508170 381250 508226
rect 381306 508170 381374 508226
rect 381430 508170 381498 508226
rect 381554 508170 381622 508226
rect 381678 508170 399250 508226
rect 399306 508170 399374 508226
rect 399430 508170 399498 508226
rect 399554 508170 399622 508226
rect 399678 508170 417250 508226
rect 417306 508170 417374 508226
rect 417430 508170 417498 508226
rect 417554 508170 417622 508226
rect 417678 508170 435250 508226
rect 435306 508170 435374 508226
rect 435430 508170 435498 508226
rect 435554 508170 435622 508226
rect 435678 508170 453250 508226
rect 453306 508170 453374 508226
rect 453430 508170 453498 508226
rect 453554 508170 453622 508226
rect 453678 508170 471250 508226
rect 471306 508170 471374 508226
rect 471430 508170 471498 508226
rect 471554 508170 471622 508226
rect 471678 508170 489250 508226
rect 489306 508170 489374 508226
rect 489430 508170 489498 508226
rect 489554 508170 489622 508226
rect 489678 508170 507250 508226
rect 507306 508170 507374 508226
rect 507430 508170 507498 508226
rect 507554 508170 507622 508226
rect 507678 508170 525250 508226
rect 525306 508170 525374 508226
rect 525430 508170 525498 508226
rect 525554 508170 525622 508226
rect 525678 508170 543250 508226
rect 543306 508170 543374 508226
rect 543430 508170 543498 508226
rect 543554 508170 543622 508226
rect 543678 508170 561250 508226
rect 561306 508170 561374 508226
rect 561430 508170 561498 508226
rect 561554 508170 561622 508226
rect 561678 508170 579250 508226
rect 579306 508170 579374 508226
rect 579430 508170 579498 508226
rect 579554 508170 579622 508226
rect 579678 508170 596496 508226
rect 596552 508170 596620 508226
rect 596676 508170 596744 508226
rect 596800 508170 596868 508226
rect 596924 508170 597980 508226
rect -1916 508102 597980 508170
rect -1916 508046 -860 508102
rect -804 508046 -736 508102
rect -680 508046 -612 508102
rect -556 508046 -488 508102
rect -432 508046 3250 508102
rect 3306 508046 3374 508102
rect 3430 508046 3498 508102
rect 3554 508046 3622 508102
rect 3678 508046 21250 508102
rect 21306 508046 21374 508102
rect 21430 508046 21498 508102
rect 21554 508046 21622 508102
rect 21678 508046 39250 508102
rect 39306 508046 39374 508102
rect 39430 508046 39498 508102
rect 39554 508046 39622 508102
rect 39678 508046 57250 508102
rect 57306 508046 57374 508102
rect 57430 508046 57498 508102
rect 57554 508046 57622 508102
rect 57678 508046 75250 508102
rect 75306 508046 75374 508102
rect 75430 508046 75498 508102
rect 75554 508046 75622 508102
rect 75678 508046 93250 508102
rect 93306 508046 93374 508102
rect 93430 508046 93498 508102
rect 93554 508046 93622 508102
rect 93678 508046 111250 508102
rect 111306 508046 111374 508102
rect 111430 508046 111498 508102
rect 111554 508046 111622 508102
rect 111678 508046 129250 508102
rect 129306 508046 129374 508102
rect 129430 508046 129498 508102
rect 129554 508046 129622 508102
rect 129678 508046 147250 508102
rect 147306 508046 147374 508102
rect 147430 508046 147498 508102
rect 147554 508046 147622 508102
rect 147678 508046 165250 508102
rect 165306 508046 165374 508102
rect 165430 508046 165498 508102
rect 165554 508046 165622 508102
rect 165678 508046 183250 508102
rect 183306 508046 183374 508102
rect 183430 508046 183498 508102
rect 183554 508046 183622 508102
rect 183678 508046 201250 508102
rect 201306 508046 201374 508102
rect 201430 508046 201498 508102
rect 201554 508046 201622 508102
rect 201678 508046 219250 508102
rect 219306 508046 219374 508102
rect 219430 508046 219498 508102
rect 219554 508046 219622 508102
rect 219678 508046 237250 508102
rect 237306 508046 237374 508102
rect 237430 508046 237498 508102
rect 237554 508046 237622 508102
rect 237678 508046 255250 508102
rect 255306 508046 255374 508102
rect 255430 508046 255498 508102
rect 255554 508046 255622 508102
rect 255678 508046 273250 508102
rect 273306 508046 273374 508102
rect 273430 508046 273498 508102
rect 273554 508046 273622 508102
rect 273678 508046 291250 508102
rect 291306 508046 291374 508102
rect 291430 508046 291498 508102
rect 291554 508046 291622 508102
rect 291678 508046 309250 508102
rect 309306 508046 309374 508102
rect 309430 508046 309498 508102
rect 309554 508046 309622 508102
rect 309678 508046 327250 508102
rect 327306 508046 327374 508102
rect 327430 508046 327498 508102
rect 327554 508046 327622 508102
rect 327678 508046 345250 508102
rect 345306 508046 345374 508102
rect 345430 508046 345498 508102
rect 345554 508046 345622 508102
rect 345678 508046 363250 508102
rect 363306 508046 363374 508102
rect 363430 508046 363498 508102
rect 363554 508046 363622 508102
rect 363678 508046 381250 508102
rect 381306 508046 381374 508102
rect 381430 508046 381498 508102
rect 381554 508046 381622 508102
rect 381678 508046 399250 508102
rect 399306 508046 399374 508102
rect 399430 508046 399498 508102
rect 399554 508046 399622 508102
rect 399678 508046 417250 508102
rect 417306 508046 417374 508102
rect 417430 508046 417498 508102
rect 417554 508046 417622 508102
rect 417678 508046 435250 508102
rect 435306 508046 435374 508102
rect 435430 508046 435498 508102
rect 435554 508046 435622 508102
rect 435678 508046 453250 508102
rect 453306 508046 453374 508102
rect 453430 508046 453498 508102
rect 453554 508046 453622 508102
rect 453678 508046 471250 508102
rect 471306 508046 471374 508102
rect 471430 508046 471498 508102
rect 471554 508046 471622 508102
rect 471678 508046 489250 508102
rect 489306 508046 489374 508102
rect 489430 508046 489498 508102
rect 489554 508046 489622 508102
rect 489678 508046 507250 508102
rect 507306 508046 507374 508102
rect 507430 508046 507498 508102
rect 507554 508046 507622 508102
rect 507678 508046 525250 508102
rect 525306 508046 525374 508102
rect 525430 508046 525498 508102
rect 525554 508046 525622 508102
rect 525678 508046 543250 508102
rect 543306 508046 543374 508102
rect 543430 508046 543498 508102
rect 543554 508046 543622 508102
rect 543678 508046 561250 508102
rect 561306 508046 561374 508102
rect 561430 508046 561498 508102
rect 561554 508046 561622 508102
rect 561678 508046 579250 508102
rect 579306 508046 579374 508102
rect 579430 508046 579498 508102
rect 579554 508046 579622 508102
rect 579678 508046 596496 508102
rect 596552 508046 596620 508102
rect 596676 508046 596744 508102
rect 596800 508046 596868 508102
rect 596924 508046 597980 508102
rect -1916 507978 597980 508046
rect -1916 507922 -860 507978
rect -804 507922 -736 507978
rect -680 507922 -612 507978
rect -556 507922 -488 507978
rect -432 507922 3250 507978
rect 3306 507922 3374 507978
rect 3430 507922 3498 507978
rect 3554 507922 3622 507978
rect 3678 507922 21250 507978
rect 21306 507922 21374 507978
rect 21430 507922 21498 507978
rect 21554 507922 21622 507978
rect 21678 507922 39250 507978
rect 39306 507922 39374 507978
rect 39430 507922 39498 507978
rect 39554 507922 39622 507978
rect 39678 507922 57250 507978
rect 57306 507922 57374 507978
rect 57430 507922 57498 507978
rect 57554 507922 57622 507978
rect 57678 507922 75250 507978
rect 75306 507922 75374 507978
rect 75430 507922 75498 507978
rect 75554 507922 75622 507978
rect 75678 507922 93250 507978
rect 93306 507922 93374 507978
rect 93430 507922 93498 507978
rect 93554 507922 93622 507978
rect 93678 507922 111250 507978
rect 111306 507922 111374 507978
rect 111430 507922 111498 507978
rect 111554 507922 111622 507978
rect 111678 507922 129250 507978
rect 129306 507922 129374 507978
rect 129430 507922 129498 507978
rect 129554 507922 129622 507978
rect 129678 507922 147250 507978
rect 147306 507922 147374 507978
rect 147430 507922 147498 507978
rect 147554 507922 147622 507978
rect 147678 507922 165250 507978
rect 165306 507922 165374 507978
rect 165430 507922 165498 507978
rect 165554 507922 165622 507978
rect 165678 507922 183250 507978
rect 183306 507922 183374 507978
rect 183430 507922 183498 507978
rect 183554 507922 183622 507978
rect 183678 507922 201250 507978
rect 201306 507922 201374 507978
rect 201430 507922 201498 507978
rect 201554 507922 201622 507978
rect 201678 507922 219250 507978
rect 219306 507922 219374 507978
rect 219430 507922 219498 507978
rect 219554 507922 219622 507978
rect 219678 507922 237250 507978
rect 237306 507922 237374 507978
rect 237430 507922 237498 507978
rect 237554 507922 237622 507978
rect 237678 507922 255250 507978
rect 255306 507922 255374 507978
rect 255430 507922 255498 507978
rect 255554 507922 255622 507978
rect 255678 507922 273250 507978
rect 273306 507922 273374 507978
rect 273430 507922 273498 507978
rect 273554 507922 273622 507978
rect 273678 507922 291250 507978
rect 291306 507922 291374 507978
rect 291430 507922 291498 507978
rect 291554 507922 291622 507978
rect 291678 507922 309250 507978
rect 309306 507922 309374 507978
rect 309430 507922 309498 507978
rect 309554 507922 309622 507978
rect 309678 507922 327250 507978
rect 327306 507922 327374 507978
rect 327430 507922 327498 507978
rect 327554 507922 327622 507978
rect 327678 507922 345250 507978
rect 345306 507922 345374 507978
rect 345430 507922 345498 507978
rect 345554 507922 345622 507978
rect 345678 507922 363250 507978
rect 363306 507922 363374 507978
rect 363430 507922 363498 507978
rect 363554 507922 363622 507978
rect 363678 507922 381250 507978
rect 381306 507922 381374 507978
rect 381430 507922 381498 507978
rect 381554 507922 381622 507978
rect 381678 507922 399250 507978
rect 399306 507922 399374 507978
rect 399430 507922 399498 507978
rect 399554 507922 399622 507978
rect 399678 507922 417250 507978
rect 417306 507922 417374 507978
rect 417430 507922 417498 507978
rect 417554 507922 417622 507978
rect 417678 507922 435250 507978
rect 435306 507922 435374 507978
rect 435430 507922 435498 507978
rect 435554 507922 435622 507978
rect 435678 507922 453250 507978
rect 453306 507922 453374 507978
rect 453430 507922 453498 507978
rect 453554 507922 453622 507978
rect 453678 507922 471250 507978
rect 471306 507922 471374 507978
rect 471430 507922 471498 507978
rect 471554 507922 471622 507978
rect 471678 507922 489250 507978
rect 489306 507922 489374 507978
rect 489430 507922 489498 507978
rect 489554 507922 489622 507978
rect 489678 507922 507250 507978
rect 507306 507922 507374 507978
rect 507430 507922 507498 507978
rect 507554 507922 507622 507978
rect 507678 507922 525250 507978
rect 525306 507922 525374 507978
rect 525430 507922 525498 507978
rect 525554 507922 525622 507978
rect 525678 507922 543250 507978
rect 543306 507922 543374 507978
rect 543430 507922 543498 507978
rect 543554 507922 543622 507978
rect 543678 507922 561250 507978
rect 561306 507922 561374 507978
rect 561430 507922 561498 507978
rect 561554 507922 561622 507978
rect 561678 507922 579250 507978
rect 579306 507922 579374 507978
rect 579430 507922 579498 507978
rect 579554 507922 579622 507978
rect 579678 507922 596496 507978
rect 596552 507922 596620 507978
rect 596676 507922 596744 507978
rect 596800 507922 596868 507978
rect 596924 507922 597980 507978
rect -1916 507826 597980 507922
rect -1916 496350 597980 496446
rect -1916 496294 -1820 496350
rect -1764 496294 -1696 496350
rect -1640 496294 -1572 496350
rect -1516 496294 -1448 496350
rect -1392 496294 6970 496350
rect 7026 496294 7094 496350
rect 7150 496294 7218 496350
rect 7274 496294 7342 496350
rect 7398 496294 24970 496350
rect 25026 496294 25094 496350
rect 25150 496294 25218 496350
rect 25274 496294 25342 496350
rect 25398 496294 42970 496350
rect 43026 496294 43094 496350
rect 43150 496294 43218 496350
rect 43274 496294 43342 496350
rect 43398 496294 60970 496350
rect 61026 496294 61094 496350
rect 61150 496294 61218 496350
rect 61274 496294 61342 496350
rect 61398 496294 78970 496350
rect 79026 496294 79094 496350
rect 79150 496294 79218 496350
rect 79274 496294 79342 496350
rect 79398 496294 96970 496350
rect 97026 496294 97094 496350
rect 97150 496294 97218 496350
rect 97274 496294 97342 496350
rect 97398 496294 114970 496350
rect 115026 496294 115094 496350
rect 115150 496294 115218 496350
rect 115274 496294 115342 496350
rect 115398 496294 132970 496350
rect 133026 496294 133094 496350
rect 133150 496294 133218 496350
rect 133274 496294 133342 496350
rect 133398 496294 150970 496350
rect 151026 496294 151094 496350
rect 151150 496294 151218 496350
rect 151274 496294 151342 496350
rect 151398 496294 168970 496350
rect 169026 496294 169094 496350
rect 169150 496294 169218 496350
rect 169274 496294 169342 496350
rect 169398 496294 186970 496350
rect 187026 496294 187094 496350
rect 187150 496294 187218 496350
rect 187274 496294 187342 496350
rect 187398 496294 204970 496350
rect 205026 496294 205094 496350
rect 205150 496294 205218 496350
rect 205274 496294 205342 496350
rect 205398 496294 222970 496350
rect 223026 496294 223094 496350
rect 223150 496294 223218 496350
rect 223274 496294 223342 496350
rect 223398 496294 240970 496350
rect 241026 496294 241094 496350
rect 241150 496294 241218 496350
rect 241274 496294 241342 496350
rect 241398 496294 258970 496350
rect 259026 496294 259094 496350
rect 259150 496294 259218 496350
rect 259274 496294 259342 496350
rect 259398 496294 276970 496350
rect 277026 496294 277094 496350
rect 277150 496294 277218 496350
rect 277274 496294 277342 496350
rect 277398 496294 294970 496350
rect 295026 496294 295094 496350
rect 295150 496294 295218 496350
rect 295274 496294 295342 496350
rect 295398 496294 312970 496350
rect 313026 496294 313094 496350
rect 313150 496294 313218 496350
rect 313274 496294 313342 496350
rect 313398 496294 330970 496350
rect 331026 496294 331094 496350
rect 331150 496294 331218 496350
rect 331274 496294 331342 496350
rect 331398 496294 348970 496350
rect 349026 496294 349094 496350
rect 349150 496294 349218 496350
rect 349274 496294 349342 496350
rect 349398 496294 366970 496350
rect 367026 496294 367094 496350
rect 367150 496294 367218 496350
rect 367274 496294 367342 496350
rect 367398 496294 384970 496350
rect 385026 496294 385094 496350
rect 385150 496294 385218 496350
rect 385274 496294 385342 496350
rect 385398 496294 402970 496350
rect 403026 496294 403094 496350
rect 403150 496294 403218 496350
rect 403274 496294 403342 496350
rect 403398 496294 420970 496350
rect 421026 496294 421094 496350
rect 421150 496294 421218 496350
rect 421274 496294 421342 496350
rect 421398 496294 438970 496350
rect 439026 496294 439094 496350
rect 439150 496294 439218 496350
rect 439274 496294 439342 496350
rect 439398 496294 456970 496350
rect 457026 496294 457094 496350
rect 457150 496294 457218 496350
rect 457274 496294 457342 496350
rect 457398 496294 474970 496350
rect 475026 496294 475094 496350
rect 475150 496294 475218 496350
rect 475274 496294 475342 496350
rect 475398 496294 492970 496350
rect 493026 496294 493094 496350
rect 493150 496294 493218 496350
rect 493274 496294 493342 496350
rect 493398 496294 510970 496350
rect 511026 496294 511094 496350
rect 511150 496294 511218 496350
rect 511274 496294 511342 496350
rect 511398 496294 528970 496350
rect 529026 496294 529094 496350
rect 529150 496294 529218 496350
rect 529274 496294 529342 496350
rect 529398 496294 546970 496350
rect 547026 496294 547094 496350
rect 547150 496294 547218 496350
rect 547274 496294 547342 496350
rect 547398 496294 564970 496350
rect 565026 496294 565094 496350
rect 565150 496294 565218 496350
rect 565274 496294 565342 496350
rect 565398 496294 582970 496350
rect 583026 496294 583094 496350
rect 583150 496294 583218 496350
rect 583274 496294 583342 496350
rect 583398 496294 597456 496350
rect 597512 496294 597580 496350
rect 597636 496294 597704 496350
rect 597760 496294 597828 496350
rect 597884 496294 597980 496350
rect -1916 496226 597980 496294
rect -1916 496170 -1820 496226
rect -1764 496170 -1696 496226
rect -1640 496170 -1572 496226
rect -1516 496170 -1448 496226
rect -1392 496170 6970 496226
rect 7026 496170 7094 496226
rect 7150 496170 7218 496226
rect 7274 496170 7342 496226
rect 7398 496170 24970 496226
rect 25026 496170 25094 496226
rect 25150 496170 25218 496226
rect 25274 496170 25342 496226
rect 25398 496170 42970 496226
rect 43026 496170 43094 496226
rect 43150 496170 43218 496226
rect 43274 496170 43342 496226
rect 43398 496170 60970 496226
rect 61026 496170 61094 496226
rect 61150 496170 61218 496226
rect 61274 496170 61342 496226
rect 61398 496170 78970 496226
rect 79026 496170 79094 496226
rect 79150 496170 79218 496226
rect 79274 496170 79342 496226
rect 79398 496170 96970 496226
rect 97026 496170 97094 496226
rect 97150 496170 97218 496226
rect 97274 496170 97342 496226
rect 97398 496170 114970 496226
rect 115026 496170 115094 496226
rect 115150 496170 115218 496226
rect 115274 496170 115342 496226
rect 115398 496170 132970 496226
rect 133026 496170 133094 496226
rect 133150 496170 133218 496226
rect 133274 496170 133342 496226
rect 133398 496170 150970 496226
rect 151026 496170 151094 496226
rect 151150 496170 151218 496226
rect 151274 496170 151342 496226
rect 151398 496170 168970 496226
rect 169026 496170 169094 496226
rect 169150 496170 169218 496226
rect 169274 496170 169342 496226
rect 169398 496170 186970 496226
rect 187026 496170 187094 496226
rect 187150 496170 187218 496226
rect 187274 496170 187342 496226
rect 187398 496170 204970 496226
rect 205026 496170 205094 496226
rect 205150 496170 205218 496226
rect 205274 496170 205342 496226
rect 205398 496170 222970 496226
rect 223026 496170 223094 496226
rect 223150 496170 223218 496226
rect 223274 496170 223342 496226
rect 223398 496170 240970 496226
rect 241026 496170 241094 496226
rect 241150 496170 241218 496226
rect 241274 496170 241342 496226
rect 241398 496170 258970 496226
rect 259026 496170 259094 496226
rect 259150 496170 259218 496226
rect 259274 496170 259342 496226
rect 259398 496170 276970 496226
rect 277026 496170 277094 496226
rect 277150 496170 277218 496226
rect 277274 496170 277342 496226
rect 277398 496170 294970 496226
rect 295026 496170 295094 496226
rect 295150 496170 295218 496226
rect 295274 496170 295342 496226
rect 295398 496170 312970 496226
rect 313026 496170 313094 496226
rect 313150 496170 313218 496226
rect 313274 496170 313342 496226
rect 313398 496170 330970 496226
rect 331026 496170 331094 496226
rect 331150 496170 331218 496226
rect 331274 496170 331342 496226
rect 331398 496170 348970 496226
rect 349026 496170 349094 496226
rect 349150 496170 349218 496226
rect 349274 496170 349342 496226
rect 349398 496170 366970 496226
rect 367026 496170 367094 496226
rect 367150 496170 367218 496226
rect 367274 496170 367342 496226
rect 367398 496170 384970 496226
rect 385026 496170 385094 496226
rect 385150 496170 385218 496226
rect 385274 496170 385342 496226
rect 385398 496170 402970 496226
rect 403026 496170 403094 496226
rect 403150 496170 403218 496226
rect 403274 496170 403342 496226
rect 403398 496170 420970 496226
rect 421026 496170 421094 496226
rect 421150 496170 421218 496226
rect 421274 496170 421342 496226
rect 421398 496170 438970 496226
rect 439026 496170 439094 496226
rect 439150 496170 439218 496226
rect 439274 496170 439342 496226
rect 439398 496170 456970 496226
rect 457026 496170 457094 496226
rect 457150 496170 457218 496226
rect 457274 496170 457342 496226
rect 457398 496170 474970 496226
rect 475026 496170 475094 496226
rect 475150 496170 475218 496226
rect 475274 496170 475342 496226
rect 475398 496170 492970 496226
rect 493026 496170 493094 496226
rect 493150 496170 493218 496226
rect 493274 496170 493342 496226
rect 493398 496170 510970 496226
rect 511026 496170 511094 496226
rect 511150 496170 511218 496226
rect 511274 496170 511342 496226
rect 511398 496170 528970 496226
rect 529026 496170 529094 496226
rect 529150 496170 529218 496226
rect 529274 496170 529342 496226
rect 529398 496170 546970 496226
rect 547026 496170 547094 496226
rect 547150 496170 547218 496226
rect 547274 496170 547342 496226
rect 547398 496170 564970 496226
rect 565026 496170 565094 496226
rect 565150 496170 565218 496226
rect 565274 496170 565342 496226
rect 565398 496170 582970 496226
rect 583026 496170 583094 496226
rect 583150 496170 583218 496226
rect 583274 496170 583342 496226
rect 583398 496170 597456 496226
rect 597512 496170 597580 496226
rect 597636 496170 597704 496226
rect 597760 496170 597828 496226
rect 597884 496170 597980 496226
rect -1916 496102 597980 496170
rect -1916 496046 -1820 496102
rect -1764 496046 -1696 496102
rect -1640 496046 -1572 496102
rect -1516 496046 -1448 496102
rect -1392 496046 6970 496102
rect 7026 496046 7094 496102
rect 7150 496046 7218 496102
rect 7274 496046 7342 496102
rect 7398 496046 24970 496102
rect 25026 496046 25094 496102
rect 25150 496046 25218 496102
rect 25274 496046 25342 496102
rect 25398 496046 42970 496102
rect 43026 496046 43094 496102
rect 43150 496046 43218 496102
rect 43274 496046 43342 496102
rect 43398 496046 60970 496102
rect 61026 496046 61094 496102
rect 61150 496046 61218 496102
rect 61274 496046 61342 496102
rect 61398 496046 78970 496102
rect 79026 496046 79094 496102
rect 79150 496046 79218 496102
rect 79274 496046 79342 496102
rect 79398 496046 96970 496102
rect 97026 496046 97094 496102
rect 97150 496046 97218 496102
rect 97274 496046 97342 496102
rect 97398 496046 114970 496102
rect 115026 496046 115094 496102
rect 115150 496046 115218 496102
rect 115274 496046 115342 496102
rect 115398 496046 132970 496102
rect 133026 496046 133094 496102
rect 133150 496046 133218 496102
rect 133274 496046 133342 496102
rect 133398 496046 150970 496102
rect 151026 496046 151094 496102
rect 151150 496046 151218 496102
rect 151274 496046 151342 496102
rect 151398 496046 168970 496102
rect 169026 496046 169094 496102
rect 169150 496046 169218 496102
rect 169274 496046 169342 496102
rect 169398 496046 186970 496102
rect 187026 496046 187094 496102
rect 187150 496046 187218 496102
rect 187274 496046 187342 496102
rect 187398 496046 204970 496102
rect 205026 496046 205094 496102
rect 205150 496046 205218 496102
rect 205274 496046 205342 496102
rect 205398 496046 222970 496102
rect 223026 496046 223094 496102
rect 223150 496046 223218 496102
rect 223274 496046 223342 496102
rect 223398 496046 240970 496102
rect 241026 496046 241094 496102
rect 241150 496046 241218 496102
rect 241274 496046 241342 496102
rect 241398 496046 258970 496102
rect 259026 496046 259094 496102
rect 259150 496046 259218 496102
rect 259274 496046 259342 496102
rect 259398 496046 276970 496102
rect 277026 496046 277094 496102
rect 277150 496046 277218 496102
rect 277274 496046 277342 496102
rect 277398 496046 294970 496102
rect 295026 496046 295094 496102
rect 295150 496046 295218 496102
rect 295274 496046 295342 496102
rect 295398 496046 312970 496102
rect 313026 496046 313094 496102
rect 313150 496046 313218 496102
rect 313274 496046 313342 496102
rect 313398 496046 330970 496102
rect 331026 496046 331094 496102
rect 331150 496046 331218 496102
rect 331274 496046 331342 496102
rect 331398 496046 348970 496102
rect 349026 496046 349094 496102
rect 349150 496046 349218 496102
rect 349274 496046 349342 496102
rect 349398 496046 366970 496102
rect 367026 496046 367094 496102
rect 367150 496046 367218 496102
rect 367274 496046 367342 496102
rect 367398 496046 384970 496102
rect 385026 496046 385094 496102
rect 385150 496046 385218 496102
rect 385274 496046 385342 496102
rect 385398 496046 402970 496102
rect 403026 496046 403094 496102
rect 403150 496046 403218 496102
rect 403274 496046 403342 496102
rect 403398 496046 420970 496102
rect 421026 496046 421094 496102
rect 421150 496046 421218 496102
rect 421274 496046 421342 496102
rect 421398 496046 438970 496102
rect 439026 496046 439094 496102
rect 439150 496046 439218 496102
rect 439274 496046 439342 496102
rect 439398 496046 456970 496102
rect 457026 496046 457094 496102
rect 457150 496046 457218 496102
rect 457274 496046 457342 496102
rect 457398 496046 474970 496102
rect 475026 496046 475094 496102
rect 475150 496046 475218 496102
rect 475274 496046 475342 496102
rect 475398 496046 492970 496102
rect 493026 496046 493094 496102
rect 493150 496046 493218 496102
rect 493274 496046 493342 496102
rect 493398 496046 510970 496102
rect 511026 496046 511094 496102
rect 511150 496046 511218 496102
rect 511274 496046 511342 496102
rect 511398 496046 528970 496102
rect 529026 496046 529094 496102
rect 529150 496046 529218 496102
rect 529274 496046 529342 496102
rect 529398 496046 546970 496102
rect 547026 496046 547094 496102
rect 547150 496046 547218 496102
rect 547274 496046 547342 496102
rect 547398 496046 564970 496102
rect 565026 496046 565094 496102
rect 565150 496046 565218 496102
rect 565274 496046 565342 496102
rect 565398 496046 582970 496102
rect 583026 496046 583094 496102
rect 583150 496046 583218 496102
rect 583274 496046 583342 496102
rect 583398 496046 597456 496102
rect 597512 496046 597580 496102
rect 597636 496046 597704 496102
rect 597760 496046 597828 496102
rect 597884 496046 597980 496102
rect -1916 495978 597980 496046
rect -1916 495922 -1820 495978
rect -1764 495922 -1696 495978
rect -1640 495922 -1572 495978
rect -1516 495922 -1448 495978
rect -1392 495922 6970 495978
rect 7026 495922 7094 495978
rect 7150 495922 7218 495978
rect 7274 495922 7342 495978
rect 7398 495922 24970 495978
rect 25026 495922 25094 495978
rect 25150 495922 25218 495978
rect 25274 495922 25342 495978
rect 25398 495922 42970 495978
rect 43026 495922 43094 495978
rect 43150 495922 43218 495978
rect 43274 495922 43342 495978
rect 43398 495922 60970 495978
rect 61026 495922 61094 495978
rect 61150 495922 61218 495978
rect 61274 495922 61342 495978
rect 61398 495922 78970 495978
rect 79026 495922 79094 495978
rect 79150 495922 79218 495978
rect 79274 495922 79342 495978
rect 79398 495922 96970 495978
rect 97026 495922 97094 495978
rect 97150 495922 97218 495978
rect 97274 495922 97342 495978
rect 97398 495922 114970 495978
rect 115026 495922 115094 495978
rect 115150 495922 115218 495978
rect 115274 495922 115342 495978
rect 115398 495922 132970 495978
rect 133026 495922 133094 495978
rect 133150 495922 133218 495978
rect 133274 495922 133342 495978
rect 133398 495922 150970 495978
rect 151026 495922 151094 495978
rect 151150 495922 151218 495978
rect 151274 495922 151342 495978
rect 151398 495922 168970 495978
rect 169026 495922 169094 495978
rect 169150 495922 169218 495978
rect 169274 495922 169342 495978
rect 169398 495922 186970 495978
rect 187026 495922 187094 495978
rect 187150 495922 187218 495978
rect 187274 495922 187342 495978
rect 187398 495922 204970 495978
rect 205026 495922 205094 495978
rect 205150 495922 205218 495978
rect 205274 495922 205342 495978
rect 205398 495922 222970 495978
rect 223026 495922 223094 495978
rect 223150 495922 223218 495978
rect 223274 495922 223342 495978
rect 223398 495922 240970 495978
rect 241026 495922 241094 495978
rect 241150 495922 241218 495978
rect 241274 495922 241342 495978
rect 241398 495922 258970 495978
rect 259026 495922 259094 495978
rect 259150 495922 259218 495978
rect 259274 495922 259342 495978
rect 259398 495922 276970 495978
rect 277026 495922 277094 495978
rect 277150 495922 277218 495978
rect 277274 495922 277342 495978
rect 277398 495922 294970 495978
rect 295026 495922 295094 495978
rect 295150 495922 295218 495978
rect 295274 495922 295342 495978
rect 295398 495922 312970 495978
rect 313026 495922 313094 495978
rect 313150 495922 313218 495978
rect 313274 495922 313342 495978
rect 313398 495922 330970 495978
rect 331026 495922 331094 495978
rect 331150 495922 331218 495978
rect 331274 495922 331342 495978
rect 331398 495922 348970 495978
rect 349026 495922 349094 495978
rect 349150 495922 349218 495978
rect 349274 495922 349342 495978
rect 349398 495922 366970 495978
rect 367026 495922 367094 495978
rect 367150 495922 367218 495978
rect 367274 495922 367342 495978
rect 367398 495922 384970 495978
rect 385026 495922 385094 495978
rect 385150 495922 385218 495978
rect 385274 495922 385342 495978
rect 385398 495922 402970 495978
rect 403026 495922 403094 495978
rect 403150 495922 403218 495978
rect 403274 495922 403342 495978
rect 403398 495922 420970 495978
rect 421026 495922 421094 495978
rect 421150 495922 421218 495978
rect 421274 495922 421342 495978
rect 421398 495922 438970 495978
rect 439026 495922 439094 495978
rect 439150 495922 439218 495978
rect 439274 495922 439342 495978
rect 439398 495922 456970 495978
rect 457026 495922 457094 495978
rect 457150 495922 457218 495978
rect 457274 495922 457342 495978
rect 457398 495922 474970 495978
rect 475026 495922 475094 495978
rect 475150 495922 475218 495978
rect 475274 495922 475342 495978
rect 475398 495922 492970 495978
rect 493026 495922 493094 495978
rect 493150 495922 493218 495978
rect 493274 495922 493342 495978
rect 493398 495922 510970 495978
rect 511026 495922 511094 495978
rect 511150 495922 511218 495978
rect 511274 495922 511342 495978
rect 511398 495922 528970 495978
rect 529026 495922 529094 495978
rect 529150 495922 529218 495978
rect 529274 495922 529342 495978
rect 529398 495922 546970 495978
rect 547026 495922 547094 495978
rect 547150 495922 547218 495978
rect 547274 495922 547342 495978
rect 547398 495922 564970 495978
rect 565026 495922 565094 495978
rect 565150 495922 565218 495978
rect 565274 495922 565342 495978
rect 565398 495922 582970 495978
rect 583026 495922 583094 495978
rect 583150 495922 583218 495978
rect 583274 495922 583342 495978
rect 583398 495922 597456 495978
rect 597512 495922 597580 495978
rect 597636 495922 597704 495978
rect 597760 495922 597828 495978
rect 597884 495922 597980 495978
rect -1916 495826 597980 495922
rect -1916 490350 597980 490446
rect -1916 490294 -860 490350
rect -804 490294 -736 490350
rect -680 490294 -612 490350
rect -556 490294 -488 490350
rect -432 490294 3250 490350
rect 3306 490294 3374 490350
rect 3430 490294 3498 490350
rect 3554 490294 3622 490350
rect 3678 490294 21250 490350
rect 21306 490294 21374 490350
rect 21430 490294 21498 490350
rect 21554 490294 21622 490350
rect 21678 490294 39250 490350
rect 39306 490294 39374 490350
rect 39430 490294 39498 490350
rect 39554 490294 39622 490350
rect 39678 490294 57250 490350
rect 57306 490294 57374 490350
rect 57430 490294 57498 490350
rect 57554 490294 57622 490350
rect 57678 490294 75250 490350
rect 75306 490294 75374 490350
rect 75430 490294 75498 490350
rect 75554 490294 75622 490350
rect 75678 490294 93250 490350
rect 93306 490294 93374 490350
rect 93430 490294 93498 490350
rect 93554 490294 93622 490350
rect 93678 490294 111250 490350
rect 111306 490294 111374 490350
rect 111430 490294 111498 490350
rect 111554 490294 111622 490350
rect 111678 490294 129250 490350
rect 129306 490294 129374 490350
rect 129430 490294 129498 490350
rect 129554 490294 129622 490350
rect 129678 490294 147250 490350
rect 147306 490294 147374 490350
rect 147430 490294 147498 490350
rect 147554 490294 147622 490350
rect 147678 490294 165250 490350
rect 165306 490294 165374 490350
rect 165430 490294 165498 490350
rect 165554 490294 165622 490350
rect 165678 490294 183250 490350
rect 183306 490294 183374 490350
rect 183430 490294 183498 490350
rect 183554 490294 183622 490350
rect 183678 490294 201250 490350
rect 201306 490294 201374 490350
rect 201430 490294 201498 490350
rect 201554 490294 201622 490350
rect 201678 490294 219250 490350
rect 219306 490294 219374 490350
rect 219430 490294 219498 490350
rect 219554 490294 219622 490350
rect 219678 490294 237250 490350
rect 237306 490294 237374 490350
rect 237430 490294 237498 490350
rect 237554 490294 237622 490350
rect 237678 490294 255250 490350
rect 255306 490294 255374 490350
rect 255430 490294 255498 490350
rect 255554 490294 255622 490350
rect 255678 490294 273250 490350
rect 273306 490294 273374 490350
rect 273430 490294 273498 490350
rect 273554 490294 273622 490350
rect 273678 490294 291250 490350
rect 291306 490294 291374 490350
rect 291430 490294 291498 490350
rect 291554 490294 291622 490350
rect 291678 490294 309250 490350
rect 309306 490294 309374 490350
rect 309430 490294 309498 490350
rect 309554 490294 309622 490350
rect 309678 490294 327250 490350
rect 327306 490294 327374 490350
rect 327430 490294 327498 490350
rect 327554 490294 327622 490350
rect 327678 490294 345250 490350
rect 345306 490294 345374 490350
rect 345430 490294 345498 490350
rect 345554 490294 345622 490350
rect 345678 490294 363250 490350
rect 363306 490294 363374 490350
rect 363430 490294 363498 490350
rect 363554 490294 363622 490350
rect 363678 490294 381250 490350
rect 381306 490294 381374 490350
rect 381430 490294 381498 490350
rect 381554 490294 381622 490350
rect 381678 490294 399250 490350
rect 399306 490294 399374 490350
rect 399430 490294 399498 490350
rect 399554 490294 399622 490350
rect 399678 490294 417250 490350
rect 417306 490294 417374 490350
rect 417430 490294 417498 490350
rect 417554 490294 417622 490350
rect 417678 490294 435250 490350
rect 435306 490294 435374 490350
rect 435430 490294 435498 490350
rect 435554 490294 435622 490350
rect 435678 490294 453250 490350
rect 453306 490294 453374 490350
rect 453430 490294 453498 490350
rect 453554 490294 453622 490350
rect 453678 490294 471250 490350
rect 471306 490294 471374 490350
rect 471430 490294 471498 490350
rect 471554 490294 471622 490350
rect 471678 490294 489250 490350
rect 489306 490294 489374 490350
rect 489430 490294 489498 490350
rect 489554 490294 489622 490350
rect 489678 490294 507250 490350
rect 507306 490294 507374 490350
rect 507430 490294 507498 490350
rect 507554 490294 507622 490350
rect 507678 490294 525250 490350
rect 525306 490294 525374 490350
rect 525430 490294 525498 490350
rect 525554 490294 525622 490350
rect 525678 490294 543250 490350
rect 543306 490294 543374 490350
rect 543430 490294 543498 490350
rect 543554 490294 543622 490350
rect 543678 490294 561250 490350
rect 561306 490294 561374 490350
rect 561430 490294 561498 490350
rect 561554 490294 561622 490350
rect 561678 490294 579250 490350
rect 579306 490294 579374 490350
rect 579430 490294 579498 490350
rect 579554 490294 579622 490350
rect 579678 490294 596496 490350
rect 596552 490294 596620 490350
rect 596676 490294 596744 490350
rect 596800 490294 596868 490350
rect 596924 490294 597980 490350
rect -1916 490226 597980 490294
rect -1916 490170 -860 490226
rect -804 490170 -736 490226
rect -680 490170 -612 490226
rect -556 490170 -488 490226
rect -432 490170 3250 490226
rect 3306 490170 3374 490226
rect 3430 490170 3498 490226
rect 3554 490170 3622 490226
rect 3678 490170 21250 490226
rect 21306 490170 21374 490226
rect 21430 490170 21498 490226
rect 21554 490170 21622 490226
rect 21678 490170 39250 490226
rect 39306 490170 39374 490226
rect 39430 490170 39498 490226
rect 39554 490170 39622 490226
rect 39678 490170 57250 490226
rect 57306 490170 57374 490226
rect 57430 490170 57498 490226
rect 57554 490170 57622 490226
rect 57678 490170 75250 490226
rect 75306 490170 75374 490226
rect 75430 490170 75498 490226
rect 75554 490170 75622 490226
rect 75678 490170 93250 490226
rect 93306 490170 93374 490226
rect 93430 490170 93498 490226
rect 93554 490170 93622 490226
rect 93678 490170 111250 490226
rect 111306 490170 111374 490226
rect 111430 490170 111498 490226
rect 111554 490170 111622 490226
rect 111678 490170 129250 490226
rect 129306 490170 129374 490226
rect 129430 490170 129498 490226
rect 129554 490170 129622 490226
rect 129678 490170 147250 490226
rect 147306 490170 147374 490226
rect 147430 490170 147498 490226
rect 147554 490170 147622 490226
rect 147678 490170 165250 490226
rect 165306 490170 165374 490226
rect 165430 490170 165498 490226
rect 165554 490170 165622 490226
rect 165678 490170 183250 490226
rect 183306 490170 183374 490226
rect 183430 490170 183498 490226
rect 183554 490170 183622 490226
rect 183678 490170 201250 490226
rect 201306 490170 201374 490226
rect 201430 490170 201498 490226
rect 201554 490170 201622 490226
rect 201678 490170 219250 490226
rect 219306 490170 219374 490226
rect 219430 490170 219498 490226
rect 219554 490170 219622 490226
rect 219678 490170 237250 490226
rect 237306 490170 237374 490226
rect 237430 490170 237498 490226
rect 237554 490170 237622 490226
rect 237678 490170 255250 490226
rect 255306 490170 255374 490226
rect 255430 490170 255498 490226
rect 255554 490170 255622 490226
rect 255678 490170 273250 490226
rect 273306 490170 273374 490226
rect 273430 490170 273498 490226
rect 273554 490170 273622 490226
rect 273678 490170 291250 490226
rect 291306 490170 291374 490226
rect 291430 490170 291498 490226
rect 291554 490170 291622 490226
rect 291678 490170 309250 490226
rect 309306 490170 309374 490226
rect 309430 490170 309498 490226
rect 309554 490170 309622 490226
rect 309678 490170 327250 490226
rect 327306 490170 327374 490226
rect 327430 490170 327498 490226
rect 327554 490170 327622 490226
rect 327678 490170 345250 490226
rect 345306 490170 345374 490226
rect 345430 490170 345498 490226
rect 345554 490170 345622 490226
rect 345678 490170 363250 490226
rect 363306 490170 363374 490226
rect 363430 490170 363498 490226
rect 363554 490170 363622 490226
rect 363678 490170 381250 490226
rect 381306 490170 381374 490226
rect 381430 490170 381498 490226
rect 381554 490170 381622 490226
rect 381678 490170 399250 490226
rect 399306 490170 399374 490226
rect 399430 490170 399498 490226
rect 399554 490170 399622 490226
rect 399678 490170 417250 490226
rect 417306 490170 417374 490226
rect 417430 490170 417498 490226
rect 417554 490170 417622 490226
rect 417678 490170 435250 490226
rect 435306 490170 435374 490226
rect 435430 490170 435498 490226
rect 435554 490170 435622 490226
rect 435678 490170 453250 490226
rect 453306 490170 453374 490226
rect 453430 490170 453498 490226
rect 453554 490170 453622 490226
rect 453678 490170 471250 490226
rect 471306 490170 471374 490226
rect 471430 490170 471498 490226
rect 471554 490170 471622 490226
rect 471678 490170 489250 490226
rect 489306 490170 489374 490226
rect 489430 490170 489498 490226
rect 489554 490170 489622 490226
rect 489678 490170 507250 490226
rect 507306 490170 507374 490226
rect 507430 490170 507498 490226
rect 507554 490170 507622 490226
rect 507678 490170 525250 490226
rect 525306 490170 525374 490226
rect 525430 490170 525498 490226
rect 525554 490170 525622 490226
rect 525678 490170 543250 490226
rect 543306 490170 543374 490226
rect 543430 490170 543498 490226
rect 543554 490170 543622 490226
rect 543678 490170 561250 490226
rect 561306 490170 561374 490226
rect 561430 490170 561498 490226
rect 561554 490170 561622 490226
rect 561678 490170 579250 490226
rect 579306 490170 579374 490226
rect 579430 490170 579498 490226
rect 579554 490170 579622 490226
rect 579678 490170 596496 490226
rect 596552 490170 596620 490226
rect 596676 490170 596744 490226
rect 596800 490170 596868 490226
rect 596924 490170 597980 490226
rect -1916 490102 597980 490170
rect -1916 490046 -860 490102
rect -804 490046 -736 490102
rect -680 490046 -612 490102
rect -556 490046 -488 490102
rect -432 490046 3250 490102
rect 3306 490046 3374 490102
rect 3430 490046 3498 490102
rect 3554 490046 3622 490102
rect 3678 490046 21250 490102
rect 21306 490046 21374 490102
rect 21430 490046 21498 490102
rect 21554 490046 21622 490102
rect 21678 490046 39250 490102
rect 39306 490046 39374 490102
rect 39430 490046 39498 490102
rect 39554 490046 39622 490102
rect 39678 490046 57250 490102
rect 57306 490046 57374 490102
rect 57430 490046 57498 490102
rect 57554 490046 57622 490102
rect 57678 490046 75250 490102
rect 75306 490046 75374 490102
rect 75430 490046 75498 490102
rect 75554 490046 75622 490102
rect 75678 490046 93250 490102
rect 93306 490046 93374 490102
rect 93430 490046 93498 490102
rect 93554 490046 93622 490102
rect 93678 490046 111250 490102
rect 111306 490046 111374 490102
rect 111430 490046 111498 490102
rect 111554 490046 111622 490102
rect 111678 490046 129250 490102
rect 129306 490046 129374 490102
rect 129430 490046 129498 490102
rect 129554 490046 129622 490102
rect 129678 490046 147250 490102
rect 147306 490046 147374 490102
rect 147430 490046 147498 490102
rect 147554 490046 147622 490102
rect 147678 490046 165250 490102
rect 165306 490046 165374 490102
rect 165430 490046 165498 490102
rect 165554 490046 165622 490102
rect 165678 490046 183250 490102
rect 183306 490046 183374 490102
rect 183430 490046 183498 490102
rect 183554 490046 183622 490102
rect 183678 490046 201250 490102
rect 201306 490046 201374 490102
rect 201430 490046 201498 490102
rect 201554 490046 201622 490102
rect 201678 490046 219250 490102
rect 219306 490046 219374 490102
rect 219430 490046 219498 490102
rect 219554 490046 219622 490102
rect 219678 490046 237250 490102
rect 237306 490046 237374 490102
rect 237430 490046 237498 490102
rect 237554 490046 237622 490102
rect 237678 490046 255250 490102
rect 255306 490046 255374 490102
rect 255430 490046 255498 490102
rect 255554 490046 255622 490102
rect 255678 490046 273250 490102
rect 273306 490046 273374 490102
rect 273430 490046 273498 490102
rect 273554 490046 273622 490102
rect 273678 490046 291250 490102
rect 291306 490046 291374 490102
rect 291430 490046 291498 490102
rect 291554 490046 291622 490102
rect 291678 490046 309250 490102
rect 309306 490046 309374 490102
rect 309430 490046 309498 490102
rect 309554 490046 309622 490102
rect 309678 490046 327250 490102
rect 327306 490046 327374 490102
rect 327430 490046 327498 490102
rect 327554 490046 327622 490102
rect 327678 490046 345250 490102
rect 345306 490046 345374 490102
rect 345430 490046 345498 490102
rect 345554 490046 345622 490102
rect 345678 490046 363250 490102
rect 363306 490046 363374 490102
rect 363430 490046 363498 490102
rect 363554 490046 363622 490102
rect 363678 490046 381250 490102
rect 381306 490046 381374 490102
rect 381430 490046 381498 490102
rect 381554 490046 381622 490102
rect 381678 490046 399250 490102
rect 399306 490046 399374 490102
rect 399430 490046 399498 490102
rect 399554 490046 399622 490102
rect 399678 490046 417250 490102
rect 417306 490046 417374 490102
rect 417430 490046 417498 490102
rect 417554 490046 417622 490102
rect 417678 490046 435250 490102
rect 435306 490046 435374 490102
rect 435430 490046 435498 490102
rect 435554 490046 435622 490102
rect 435678 490046 453250 490102
rect 453306 490046 453374 490102
rect 453430 490046 453498 490102
rect 453554 490046 453622 490102
rect 453678 490046 471250 490102
rect 471306 490046 471374 490102
rect 471430 490046 471498 490102
rect 471554 490046 471622 490102
rect 471678 490046 489250 490102
rect 489306 490046 489374 490102
rect 489430 490046 489498 490102
rect 489554 490046 489622 490102
rect 489678 490046 507250 490102
rect 507306 490046 507374 490102
rect 507430 490046 507498 490102
rect 507554 490046 507622 490102
rect 507678 490046 525250 490102
rect 525306 490046 525374 490102
rect 525430 490046 525498 490102
rect 525554 490046 525622 490102
rect 525678 490046 543250 490102
rect 543306 490046 543374 490102
rect 543430 490046 543498 490102
rect 543554 490046 543622 490102
rect 543678 490046 561250 490102
rect 561306 490046 561374 490102
rect 561430 490046 561498 490102
rect 561554 490046 561622 490102
rect 561678 490046 579250 490102
rect 579306 490046 579374 490102
rect 579430 490046 579498 490102
rect 579554 490046 579622 490102
rect 579678 490046 596496 490102
rect 596552 490046 596620 490102
rect 596676 490046 596744 490102
rect 596800 490046 596868 490102
rect 596924 490046 597980 490102
rect -1916 489978 597980 490046
rect -1916 489922 -860 489978
rect -804 489922 -736 489978
rect -680 489922 -612 489978
rect -556 489922 -488 489978
rect -432 489922 3250 489978
rect 3306 489922 3374 489978
rect 3430 489922 3498 489978
rect 3554 489922 3622 489978
rect 3678 489922 21250 489978
rect 21306 489922 21374 489978
rect 21430 489922 21498 489978
rect 21554 489922 21622 489978
rect 21678 489922 39250 489978
rect 39306 489922 39374 489978
rect 39430 489922 39498 489978
rect 39554 489922 39622 489978
rect 39678 489922 57250 489978
rect 57306 489922 57374 489978
rect 57430 489922 57498 489978
rect 57554 489922 57622 489978
rect 57678 489922 75250 489978
rect 75306 489922 75374 489978
rect 75430 489922 75498 489978
rect 75554 489922 75622 489978
rect 75678 489922 93250 489978
rect 93306 489922 93374 489978
rect 93430 489922 93498 489978
rect 93554 489922 93622 489978
rect 93678 489922 111250 489978
rect 111306 489922 111374 489978
rect 111430 489922 111498 489978
rect 111554 489922 111622 489978
rect 111678 489922 129250 489978
rect 129306 489922 129374 489978
rect 129430 489922 129498 489978
rect 129554 489922 129622 489978
rect 129678 489922 147250 489978
rect 147306 489922 147374 489978
rect 147430 489922 147498 489978
rect 147554 489922 147622 489978
rect 147678 489922 165250 489978
rect 165306 489922 165374 489978
rect 165430 489922 165498 489978
rect 165554 489922 165622 489978
rect 165678 489922 183250 489978
rect 183306 489922 183374 489978
rect 183430 489922 183498 489978
rect 183554 489922 183622 489978
rect 183678 489922 201250 489978
rect 201306 489922 201374 489978
rect 201430 489922 201498 489978
rect 201554 489922 201622 489978
rect 201678 489922 219250 489978
rect 219306 489922 219374 489978
rect 219430 489922 219498 489978
rect 219554 489922 219622 489978
rect 219678 489922 237250 489978
rect 237306 489922 237374 489978
rect 237430 489922 237498 489978
rect 237554 489922 237622 489978
rect 237678 489922 255250 489978
rect 255306 489922 255374 489978
rect 255430 489922 255498 489978
rect 255554 489922 255622 489978
rect 255678 489922 273250 489978
rect 273306 489922 273374 489978
rect 273430 489922 273498 489978
rect 273554 489922 273622 489978
rect 273678 489922 291250 489978
rect 291306 489922 291374 489978
rect 291430 489922 291498 489978
rect 291554 489922 291622 489978
rect 291678 489922 309250 489978
rect 309306 489922 309374 489978
rect 309430 489922 309498 489978
rect 309554 489922 309622 489978
rect 309678 489922 327250 489978
rect 327306 489922 327374 489978
rect 327430 489922 327498 489978
rect 327554 489922 327622 489978
rect 327678 489922 345250 489978
rect 345306 489922 345374 489978
rect 345430 489922 345498 489978
rect 345554 489922 345622 489978
rect 345678 489922 363250 489978
rect 363306 489922 363374 489978
rect 363430 489922 363498 489978
rect 363554 489922 363622 489978
rect 363678 489922 381250 489978
rect 381306 489922 381374 489978
rect 381430 489922 381498 489978
rect 381554 489922 381622 489978
rect 381678 489922 399250 489978
rect 399306 489922 399374 489978
rect 399430 489922 399498 489978
rect 399554 489922 399622 489978
rect 399678 489922 417250 489978
rect 417306 489922 417374 489978
rect 417430 489922 417498 489978
rect 417554 489922 417622 489978
rect 417678 489922 435250 489978
rect 435306 489922 435374 489978
rect 435430 489922 435498 489978
rect 435554 489922 435622 489978
rect 435678 489922 453250 489978
rect 453306 489922 453374 489978
rect 453430 489922 453498 489978
rect 453554 489922 453622 489978
rect 453678 489922 471250 489978
rect 471306 489922 471374 489978
rect 471430 489922 471498 489978
rect 471554 489922 471622 489978
rect 471678 489922 489250 489978
rect 489306 489922 489374 489978
rect 489430 489922 489498 489978
rect 489554 489922 489622 489978
rect 489678 489922 507250 489978
rect 507306 489922 507374 489978
rect 507430 489922 507498 489978
rect 507554 489922 507622 489978
rect 507678 489922 525250 489978
rect 525306 489922 525374 489978
rect 525430 489922 525498 489978
rect 525554 489922 525622 489978
rect 525678 489922 543250 489978
rect 543306 489922 543374 489978
rect 543430 489922 543498 489978
rect 543554 489922 543622 489978
rect 543678 489922 561250 489978
rect 561306 489922 561374 489978
rect 561430 489922 561498 489978
rect 561554 489922 561622 489978
rect 561678 489922 579250 489978
rect 579306 489922 579374 489978
rect 579430 489922 579498 489978
rect 579554 489922 579622 489978
rect 579678 489922 596496 489978
rect 596552 489922 596620 489978
rect 596676 489922 596744 489978
rect 596800 489922 596868 489978
rect 596924 489922 597980 489978
rect -1916 489826 597980 489922
rect -1916 478350 597980 478446
rect -1916 478294 -1820 478350
rect -1764 478294 -1696 478350
rect -1640 478294 -1572 478350
rect -1516 478294 -1448 478350
rect -1392 478294 6970 478350
rect 7026 478294 7094 478350
rect 7150 478294 7218 478350
rect 7274 478294 7342 478350
rect 7398 478294 24970 478350
rect 25026 478294 25094 478350
rect 25150 478294 25218 478350
rect 25274 478294 25342 478350
rect 25398 478294 42970 478350
rect 43026 478294 43094 478350
rect 43150 478294 43218 478350
rect 43274 478294 43342 478350
rect 43398 478294 60970 478350
rect 61026 478294 61094 478350
rect 61150 478294 61218 478350
rect 61274 478294 61342 478350
rect 61398 478294 78970 478350
rect 79026 478294 79094 478350
rect 79150 478294 79218 478350
rect 79274 478294 79342 478350
rect 79398 478294 96970 478350
rect 97026 478294 97094 478350
rect 97150 478294 97218 478350
rect 97274 478294 97342 478350
rect 97398 478294 114970 478350
rect 115026 478294 115094 478350
rect 115150 478294 115218 478350
rect 115274 478294 115342 478350
rect 115398 478294 132970 478350
rect 133026 478294 133094 478350
rect 133150 478294 133218 478350
rect 133274 478294 133342 478350
rect 133398 478294 150970 478350
rect 151026 478294 151094 478350
rect 151150 478294 151218 478350
rect 151274 478294 151342 478350
rect 151398 478294 168970 478350
rect 169026 478294 169094 478350
rect 169150 478294 169218 478350
rect 169274 478294 169342 478350
rect 169398 478294 186970 478350
rect 187026 478294 187094 478350
rect 187150 478294 187218 478350
rect 187274 478294 187342 478350
rect 187398 478294 204970 478350
rect 205026 478294 205094 478350
rect 205150 478294 205218 478350
rect 205274 478294 205342 478350
rect 205398 478294 222970 478350
rect 223026 478294 223094 478350
rect 223150 478294 223218 478350
rect 223274 478294 223342 478350
rect 223398 478294 240970 478350
rect 241026 478294 241094 478350
rect 241150 478294 241218 478350
rect 241274 478294 241342 478350
rect 241398 478294 258970 478350
rect 259026 478294 259094 478350
rect 259150 478294 259218 478350
rect 259274 478294 259342 478350
rect 259398 478294 276970 478350
rect 277026 478294 277094 478350
rect 277150 478294 277218 478350
rect 277274 478294 277342 478350
rect 277398 478294 294970 478350
rect 295026 478294 295094 478350
rect 295150 478294 295218 478350
rect 295274 478294 295342 478350
rect 295398 478294 312970 478350
rect 313026 478294 313094 478350
rect 313150 478294 313218 478350
rect 313274 478294 313342 478350
rect 313398 478294 330970 478350
rect 331026 478294 331094 478350
rect 331150 478294 331218 478350
rect 331274 478294 331342 478350
rect 331398 478294 348970 478350
rect 349026 478294 349094 478350
rect 349150 478294 349218 478350
rect 349274 478294 349342 478350
rect 349398 478294 366970 478350
rect 367026 478294 367094 478350
rect 367150 478294 367218 478350
rect 367274 478294 367342 478350
rect 367398 478294 384970 478350
rect 385026 478294 385094 478350
rect 385150 478294 385218 478350
rect 385274 478294 385342 478350
rect 385398 478294 402970 478350
rect 403026 478294 403094 478350
rect 403150 478294 403218 478350
rect 403274 478294 403342 478350
rect 403398 478294 420970 478350
rect 421026 478294 421094 478350
rect 421150 478294 421218 478350
rect 421274 478294 421342 478350
rect 421398 478294 438970 478350
rect 439026 478294 439094 478350
rect 439150 478294 439218 478350
rect 439274 478294 439342 478350
rect 439398 478294 456970 478350
rect 457026 478294 457094 478350
rect 457150 478294 457218 478350
rect 457274 478294 457342 478350
rect 457398 478294 474970 478350
rect 475026 478294 475094 478350
rect 475150 478294 475218 478350
rect 475274 478294 475342 478350
rect 475398 478294 492970 478350
rect 493026 478294 493094 478350
rect 493150 478294 493218 478350
rect 493274 478294 493342 478350
rect 493398 478294 510970 478350
rect 511026 478294 511094 478350
rect 511150 478294 511218 478350
rect 511274 478294 511342 478350
rect 511398 478294 528970 478350
rect 529026 478294 529094 478350
rect 529150 478294 529218 478350
rect 529274 478294 529342 478350
rect 529398 478294 546970 478350
rect 547026 478294 547094 478350
rect 547150 478294 547218 478350
rect 547274 478294 547342 478350
rect 547398 478294 564970 478350
rect 565026 478294 565094 478350
rect 565150 478294 565218 478350
rect 565274 478294 565342 478350
rect 565398 478294 582970 478350
rect 583026 478294 583094 478350
rect 583150 478294 583218 478350
rect 583274 478294 583342 478350
rect 583398 478294 597456 478350
rect 597512 478294 597580 478350
rect 597636 478294 597704 478350
rect 597760 478294 597828 478350
rect 597884 478294 597980 478350
rect -1916 478226 597980 478294
rect -1916 478170 -1820 478226
rect -1764 478170 -1696 478226
rect -1640 478170 -1572 478226
rect -1516 478170 -1448 478226
rect -1392 478170 6970 478226
rect 7026 478170 7094 478226
rect 7150 478170 7218 478226
rect 7274 478170 7342 478226
rect 7398 478170 24970 478226
rect 25026 478170 25094 478226
rect 25150 478170 25218 478226
rect 25274 478170 25342 478226
rect 25398 478170 42970 478226
rect 43026 478170 43094 478226
rect 43150 478170 43218 478226
rect 43274 478170 43342 478226
rect 43398 478170 60970 478226
rect 61026 478170 61094 478226
rect 61150 478170 61218 478226
rect 61274 478170 61342 478226
rect 61398 478170 78970 478226
rect 79026 478170 79094 478226
rect 79150 478170 79218 478226
rect 79274 478170 79342 478226
rect 79398 478170 96970 478226
rect 97026 478170 97094 478226
rect 97150 478170 97218 478226
rect 97274 478170 97342 478226
rect 97398 478170 114970 478226
rect 115026 478170 115094 478226
rect 115150 478170 115218 478226
rect 115274 478170 115342 478226
rect 115398 478170 132970 478226
rect 133026 478170 133094 478226
rect 133150 478170 133218 478226
rect 133274 478170 133342 478226
rect 133398 478170 150970 478226
rect 151026 478170 151094 478226
rect 151150 478170 151218 478226
rect 151274 478170 151342 478226
rect 151398 478170 168970 478226
rect 169026 478170 169094 478226
rect 169150 478170 169218 478226
rect 169274 478170 169342 478226
rect 169398 478170 186970 478226
rect 187026 478170 187094 478226
rect 187150 478170 187218 478226
rect 187274 478170 187342 478226
rect 187398 478170 204970 478226
rect 205026 478170 205094 478226
rect 205150 478170 205218 478226
rect 205274 478170 205342 478226
rect 205398 478170 222970 478226
rect 223026 478170 223094 478226
rect 223150 478170 223218 478226
rect 223274 478170 223342 478226
rect 223398 478170 240970 478226
rect 241026 478170 241094 478226
rect 241150 478170 241218 478226
rect 241274 478170 241342 478226
rect 241398 478170 258970 478226
rect 259026 478170 259094 478226
rect 259150 478170 259218 478226
rect 259274 478170 259342 478226
rect 259398 478170 276970 478226
rect 277026 478170 277094 478226
rect 277150 478170 277218 478226
rect 277274 478170 277342 478226
rect 277398 478170 294970 478226
rect 295026 478170 295094 478226
rect 295150 478170 295218 478226
rect 295274 478170 295342 478226
rect 295398 478170 312970 478226
rect 313026 478170 313094 478226
rect 313150 478170 313218 478226
rect 313274 478170 313342 478226
rect 313398 478170 330970 478226
rect 331026 478170 331094 478226
rect 331150 478170 331218 478226
rect 331274 478170 331342 478226
rect 331398 478170 348970 478226
rect 349026 478170 349094 478226
rect 349150 478170 349218 478226
rect 349274 478170 349342 478226
rect 349398 478170 366970 478226
rect 367026 478170 367094 478226
rect 367150 478170 367218 478226
rect 367274 478170 367342 478226
rect 367398 478170 384970 478226
rect 385026 478170 385094 478226
rect 385150 478170 385218 478226
rect 385274 478170 385342 478226
rect 385398 478170 402970 478226
rect 403026 478170 403094 478226
rect 403150 478170 403218 478226
rect 403274 478170 403342 478226
rect 403398 478170 420970 478226
rect 421026 478170 421094 478226
rect 421150 478170 421218 478226
rect 421274 478170 421342 478226
rect 421398 478170 438970 478226
rect 439026 478170 439094 478226
rect 439150 478170 439218 478226
rect 439274 478170 439342 478226
rect 439398 478170 456970 478226
rect 457026 478170 457094 478226
rect 457150 478170 457218 478226
rect 457274 478170 457342 478226
rect 457398 478170 474970 478226
rect 475026 478170 475094 478226
rect 475150 478170 475218 478226
rect 475274 478170 475342 478226
rect 475398 478170 492970 478226
rect 493026 478170 493094 478226
rect 493150 478170 493218 478226
rect 493274 478170 493342 478226
rect 493398 478170 510970 478226
rect 511026 478170 511094 478226
rect 511150 478170 511218 478226
rect 511274 478170 511342 478226
rect 511398 478170 528970 478226
rect 529026 478170 529094 478226
rect 529150 478170 529218 478226
rect 529274 478170 529342 478226
rect 529398 478170 546970 478226
rect 547026 478170 547094 478226
rect 547150 478170 547218 478226
rect 547274 478170 547342 478226
rect 547398 478170 564970 478226
rect 565026 478170 565094 478226
rect 565150 478170 565218 478226
rect 565274 478170 565342 478226
rect 565398 478170 582970 478226
rect 583026 478170 583094 478226
rect 583150 478170 583218 478226
rect 583274 478170 583342 478226
rect 583398 478170 597456 478226
rect 597512 478170 597580 478226
rect 597636 478170 597704 478226
rect 597760 478170 597828 478226
rect 597884 478170 597980 478226
rect -1916 478102 597980 478170
rect -1916 478046 -1820 478102
rect -1764 478046 -1696 478102
rect -1640 478046 -1572 478102
rect -1516 478046 -1448 478102
rect -1392 478046 6970 478102
rect 7026 478046 7094 478102
rect 7150 478046 7218 478102
rect 7274 478046 7342 478102
rect 7398 478046 24970 478102
rect 25026 478046 25094 478102
rect 25150 478046 25218 478102
rect 25274 478046 25342 478102
rect 25398 478046 42970 478102
rect 43026 478046 43094 478102
rect 43150 478046 43218 478102
rect 43274 478046 43342 478102
rect 43398 478046 60970 478102
rect 61026 478046 61094 478102
rect 61150 478046 61218 478102
rect 61274 478046 61342 478102
rect 61398 478046 78970 478102
rect 79026 478046 79094 478102
rect 79150 478046 79218 478102
rect 79274 478046 79342 478102
rect 79398 478046 96970 478102
rect 97026 478046 97094 478102
rect 97150 478046 97218 478102
rect 97274 478046 97342 478102
rect 97398 478046 114970 478102
rect 115026 478046 115094 478102
rect 115150 478046 115218 478102
rect 115274 478046 115342 478102
rect 115398 478046 132970 478102
rect 133026 478046 133094 478102
rect 133150 478046 133218 478102
rect 133274 478046 133342 478102
rect 133398 478046 150970 478102
rect 151026 478046 151094 478102
rect 151150 478046 151218 478102
rect 151274 478046 151342 478102
rect 151398 478046 168970 478102
rect 169026 478046 169094 478102
rect 169150 478046 169218 478102
rect 169274 478046 169342 478102
rect 169398 478046 186970 478102
rect 187026 478046 187094 478102
rect 187150 478046 187218 478102
rect 187274 478046 187342 478102
rect 187398 478046 204970 478102
rect 205026 478046 205094 478102
rect 205150 478046 205218 478102
rect 205274 478046 205342 478102
rect 205398 478046 222970 478102
rect 223026 478046 223094 478102
rect 223150 478046 223218 478102
rect 223274 478046 223342 478102
rect 223398 478046 240970 478102
rect 241026 478046 241094 478102
rect 241150 478046 241218 478102
rect 241274 478046 241342 478102
rect 241398 478046 258970 478102
rect 259026 478046 259094 478102
rect 259150 478046 259218 478102
rect 259274 478046 259342 478102
rect 259398 478046 276970 478102
rect 277026 478046 277094 478102
rect 277150 478046 277218 478102
rect 277274 478046 277342 478102
rect 277398 478046 294970 478102
rect 295026 478046 295094 478102
rect 295150 478046 295218 478102
rect 295274 478046 295342 478102
rect 295398 478046 312970 478102
rect 313026 478046 313094 478102
rect 313150 478046 313218 478102
rect 313274 478046 313342 478102
rect 313398 478046 330970 478102
rect 331026 478046 331094 478102
rect 331150 478046 331218 478102
rect 331274 478046 331342 478102
rect 331398 478046 348970 478102
rect 349026 478046 349094 478102
rect 349150 478046 349218 478102
rect 349274 478046 349342 478102
rect 349398 478046 366970 478102
rect 367026 478046 367094 478102
rect 367150 478046 367218 478102
rect 367274 478046 367342 478102
rect 367398 478046 384970 478102
rect 385026 478046 385094 478102
rect 385150 478046 385218 478102
rect 385274 478046 385342 478102
rect 385398 478046 402970 478102
rect 403026 478046 403094 478102
rect 403150 478046 403218 478102
rect 403274 478046 403342 478102
rect 403398 478046 420970 478102
rect 421026 478046 421094 478102
rect 421150 478046 421218 478102
rect 421274 478046 421342 478102
rect 421398 478046 438970 478102
rect 439026 478046 439094 478102
rect 439150 478046 439218 478102
rect 439274 478046 439342 478102
rect 439398 478046 456970 478102
rect 457026 478046 457094 478102
rect 457150 478046 457218 478102
rect 457274 478046 457342 478102
rect 457398 478046 474970 478102
rect 475026 478046 475094 478102
rect 475150 478046 475218 478102
rect 475274 478046 475342 478102
rect 475398 478046 492970 478102
rect 493026 478046 493094 478102
rect 493150 478046 493218 478102
rect 493274 478046 493342 478102
rect 493398 478046 510970 478102
rect 511026 478046 511094 478102
rect 511150 478046 511218 478102
rect 511274 478046 511342 478102
rect 511398 478046 528970 478102
rect 529026 478046 529094 478102
rect 529150 478046 529218 478102
rect 529274 478046 529342 478102
rect 529398 478046 546970 478102
rect 547026 478046 547094 478102
rect 547150 478046 547218 478102
rect 547274 478046 547342 478102
rect 547398 478046 564970 478102
rect 565026 478046 565094 478102
rect 565150 478046 565218 478102
rect 565274 478046 565342 478102
rect 565398 478046 582970 478102
rect 583026 478046 583094 478102
rect 583150 478046 583218 478102
rect 583274 478046 583342 478102
rect 583398 478046 597456 478102
rect 597512 478046 597580 478102
rect 597636 478046 597704 478102
rect 597760 478046 597828 478102
rect 597884 478046 597980 478102
rect -1916 477978 597980 478046
rect -1916 477922 -1820 477978
rect -1764 477922 -1696 477978
rect -1640 477922 -1572 477978
rect -1516 477922 -1448 477978
rect -1392 477922 6970 477978
rect 7026 477922 7094 477978
rect 7150 477922 7218 477978
rect 7274 477922 7342 477978
rect 7398 477922 24970 477978
rect 25026 477922 25094 477978
rect 25150 477922 25218 477978
rect 25274 477922 25342 477978
rect 25398 477922 42970 477978
rect 43026 477922 43094 477978
rect 43150 477922 43218 477978
rect 43274 477922 43342 477978
rect 43398 477922 60970 477978
rect 61026 477922 61094 477978
rect 61150 477922 61218 477978
rect 61274 477922 61342 477978
rect 61398 477922 78970 477978
rect 79026 477922 79094 477978
rect 79150 477922 79218 477978
rect 79274 477922 79342 477978
rect 79398 477922 96970 477978
rect 97026 477922 97094 477978
rect 97150 477922 97218 477978
rect 97274 477922 97342 477978
rect 97398 477922 114970 477978
rect 115026 477922 115094 477978
rect 115150 477922 115218 477978
rect 115274 477922 115342 477978
rect 115398 477922 132970 477978
rect 133026 477922 133094 477978
rect 133150 477922 133218 477978
rect 133274 477922 133342 477978
rect 133398 477922 150970 477978
rect 151026 477922 151094 477978
rect 151150 477922 151218 477978
rect 151274 477922 151342 477978
rect 151398 477922 168970 477978
rect 169026 477922 169094 477978
rect 169150 477922 169218 477978
rect 169274 477922 169342 477978
rect 169398 477922 186970 477978
rect 187026 477922 187094 477978
rect 187150 477922 187218 477978
rect 187274 477922 187342 477978
rect 187398 477922 204970 477978
rect 205026 477922 205094 477978
rect 205150 477922 205218 477978
rect 205274 477922 205342 477978
rect 205398 477922 222970 477978
rect 223026 477922 223094 477978
rect 223150 477922 223218 477978
rect 223274 477922 223342 477978
rect 223398 477922 240970 477978
rect 241026 477922 241094 477978
rect 241150 477922 241218 477978
rect 241274 477922 241342 477978
rect 241398 477922 258970 477978
rect 259026 477922 259094 477978
rect 259150 477922 259218 477978
rect 259274 477922 259342 477978
rect 259398 477922 276970 477978
rect 277026 477922 277094 477978
rect 277150 477922 277218 477978
rect 277274 477922 277342 477978
rect 277398 477922 294970 477978
rect 295026 477922 295094 477978
rect 295150 477922 295218 477978
rect 295274 477922 295342 477978
rect 295398 477922 312970 477978
rect 313026 477922 313094 477978
rect 313150 477922 313218 477978
rect 313274 477922 313342 477978
rect 313398 477922 330970 477978
rect 331026 477922 331094 477978
rect 331150 477922 331218 477978
rect 331274 477922 331342 477978
rect 331398 477922 348970 477978
rect 349026 477922 349094 477978
rect 349150 477922 349218 477978
rect 349274 477922 349342 477978
rect 349398 477922 366970 477978
rect 367026 477922 367094 477978
rect 367150 477922 367218 477978
rect 367274 477922 367342 477978
rect 367398 477922 384970 477978
rect 385026 477922 385094 477978
rect 385150 477922 385218 477978
rect 385274 477922 385342 477978
rect 385398 477922 402970 477978
rect 403026 477922 403094 477978
rect 403150 477922 403218 477978
rect 403274 477922 403342 477978
rect 403398 477922 420970 477978
rect 421026 477922 421094 477978
rect 421150 477922 421218 477978
rect 421274 477922 421342 477978
rect 421398 477922 438970 477978
rect 439026 477922 439094 477978
rect 439150 477922 439218 477978
rect 439274 477922 439342 477978
rect 439398 477922 456970 477978
rect 457026 477922 457094 477978
rect 457150 477922 457218 477978
rect 457274 477922 457342 477978
rect 457398 477922 474970 477978
rect 475026 477922 475094 477978
rect 475150 477922 475218 477978
rect 475274 477922 475342 477978
rect 475398 477922 492970 477978
rect 493026 477922 493094 477978
rect 493150 477922 493218 477978
rect 493274 477922 493342 477978
rect 493398 477922 510970 477978
rect 511026 477922 511094 477978
rect 511150 477922 511218 477978
rect 511274 477922 511342 477978
rect 511398 477922 528970 477978
rect 529026 477922 529094 477978
rect 529150 477922 529218 477978
rect 529274 477922 529342 477978
rect 529398 477922 546970 477978
rect 547026 477922 547094 477978
rect 547150 477922 547218 477978
rect 547274 477922 547342 477978
rect 547398 477922 564970 477978
rect 565026 477922 565094 477978
rect 565150 477922 565218 477978
rect 565274 477922 565342 477978
rect 565398 477922 582970 477978
rect 583026 477922 583094 477978
rect 583150 477922 583218 477978
rect 583274 477922 583342 477978
rect 583398 477922 597456 477978
rect 597512 477922 597580 477978
rect 597636 477922 597704 477978
rect 597760 477922 597828 477978
rect 597884 477922 597980 477978
rect -1916 477826 597980 477922
rect -1916 472350 597980 472446
rect -1916 472294 -860 472350
rect -804 472294 -736 472350
rect -680 472294 -612 472350
rect -556 472294 -488 472350
rect -432 472294 3250 472350
rect 3306 472294 3374 472350
rect 3430 472294 3498 472350
rect 3554 472294 3622 472350
rect 3678 472294 21250 472350
rect 21306 472294 21374 472350
rect 21430 472294 21498 472350
rect 21554 472294 21622 472350
rect 21678 472294 39250 472350
rect 39306 472294 39374 472350
rect 39430 472294 39498 472350
rect 39554 472294 39622 472350
rect 39678 472294 57250 472350
rect 57306 472294 57374 472350
rect 57430 472294 57498 472350
rect 57554 472294 57622 472350
rect 57678 472294 75250 472350
rect 75306 472294 75374 472350
rect 75430 472294 75498 472350
rect 75554 472294 75622 472350
rect 75678 472294 93250 472350
rect 93306 472294 93374 472350
rect 93430 472294 93498 472350
rect 93554 472294 93622 472350
rect 93678 472294 111250 472350
rect 111306 472294 111374 472350
rect 111430 472294 111498 472350
rect 111554 472294 111622 472350
rect 111678 472294 129250 472350
rect 129306 472294 129374 472350
rect 129430 472294 129498 472350
rect 129554 472294 129622 472350
rect 129678 472294 147250 472350
rect 147306 472294 147374 472350
rect 147430 472294 147498 472350
rect 147554 472294 147622 472350
rect 147678 472294 165250 472350
rect 165306 472294 165374 472350
rect 165430 472294 165498 472350
rect 165554 472294 165622 472350
rect 165678 472294 183250 472350
rect 183306 472294 183374 472350
rect 183430 472294 183498 472350
rect 183554 472294 183622 472350
rect 183678 472294 201250 472350
rect 201306 472294 201374 472350
rect 201430 472294 201498 472350
rect 201554 472294 201622 472350
rect 201678 472294 219250 472350
rect 219306 472294 219374 472350
rect 219430 472294 219498 472350
rect 219554 472294 219622 472350
rect 219678 472294 237250 472350
rect 237306 472294 237374 472350
rect 237430 472294 237498 472350
rect 237554 472294 237622 472350
rect 237678 472294 255250 472350
rect 255306 472294 255374 472350
rect 255430 472294 255498 472350
rect 255554 472294 255622 472350
rect 255678 472294 273250 472350
rect 273306 472294 273374 472350
rect 273430 472294 273498 472350
rect 273554 472294 273622 472350
rect 273678 472294 291250 472350
rect 291306 472294 291374 472350
rect 291430 472294 291498 472350
rect 291554 472294 291622 472350
rect 291678 472294 309250 472350
rect 309306 472294 309374 472350
rect 309430 472294 309498 472350
rect 309554 472294 309622 472350
rect 309678 472294 327250 472350
rect 327306 472294 327374 472350
rect 327430 472294 327498 472350
rect 327554 472294 327622 472350
rect 327678 472294 345250 472350
rect 345306 472294 345374 472350
rect 345430 472294 345498 472350
rect 345554 472294 345622 472350
rect 345678 472294 363250 472350
rect 363306 472294 363374 472350
rect 363430 472294 363498 472350
rect 363554 472294 363622 472350
rect 363678 472294 381250 472350
rect 381306 472294 381374 472350
rect 381430 472294 381498 472350
rect 381554 472294 381622 472350
rect 381678 472294 399250 472350
rect 399306 472294 399374 472350
rect 399430 472294 399498 472350
rect 399554 472294 399622 472350
rect 399678 472294 417250 472350
rect 417306 472294 417374 472350
rect 417430 472294 417498 472350
rect 417554 472294 417622 472350
rect 417678 472294 435250 472350
rect 435306 472294 435374 472350
rect 435430 472294 435498 472350
rect 435554 472294 435622 472350
rect 435678 472294 453250 472350
rect 453306 472294 453374 472350
rect 453430 472294 453498 472350
rect 453554 472294 453622 472350
rect 453678 472294 471250 472350
rect 471306 472294 471374 472350
rect 471430 472294 471498 472350
rect 471554 472294 471622 472350
rect 471678 472294 489250 472350
rect 489306 472294 489374 472350
rect 489430 472294 489498 472350
rect 489554 472294 489622 472350
rect 489678 472294 507250 472350
rect 507306 472294 507374 472350
rect 507430 472294 507498 472350
rect 507554 472294 507622 472350
rect 507678 472294 525250 472350
rect 525306 472294 525374 472350
rect 525430 472294 525498 472350
rect 525554 472294 525622 472350
rect 525678 472294 543250 472350
rect 543306 472294 543374 472350
rect 543430 472294 543498 472350
rect 543554 472294 543622 472350
rect 543678 472294 561250 472350
rect 561306 472294 561374 472350
rect 561430 472294 561498 472350
rect 561554 472294 561622 472350
rect 561678 472294 579250 472350
rect 579306 472294 579374 472350
rect 579430 472294 579498 472350
rect 579554 472294 579622 472350
rect 579678 472294 596496 472350
rect 596552 472294 596620 472350
rect 596676 472294 596744 472350
rect 596800 472294 596868 472350
rect 596924 472294 597980 472350
rect -1916 472226 597980 472294
rect -1916 472170 -860 472226
rect -804 472170 -736 472226
rect -680 472170 -612 472226
rect -556 472170 -488 472226
rect -432 472170 3250 472226
rect 3306 472170 3374 472226
rect 3430 472170 3498 472226
rect 3554 472170 3622 472226
rect 3678 472170 21250 472226
rect 21306 472170 21374 472226
rect 21430 472170 21498 472226
rect 21554 472170 21622 472226
rect 21678 472170 39250 472226
rect 39306 472170 39374 472226
rect 39430 472170 39498 472226
rect 39554 472170 39622 472226
rect 39678 472170 57250 472226
rect 57306 472170 57374 472226
rect 57430 472170 57498 472226
rect 57554 472170 57622 472226
rect 57678 472170 75250 472226
rect 75306 472170 75374 472226
rect 75430 472170 75498 472226
rect 75554 472170 75622 472226
rect 75678 472170 93250 472226
rect 93306 472170 93374 472226
rect 93430 472170 93498 472226
rect 93554 472170 93622 472226
rect 93678 472170 111250 472226
rect 111306 472170 111374 472226
rect 111430 472170 111498 472226
rect 111554 472170 111622 472226
rect 111678 472170 129250 472226
rect 129306 472170 129374 472226
rect 129430 472170 129498 472226
rect 129554 472170 129622 472226
rect 129678 472170 147250 472226
rect 147306 472170 147374 472226
rect 147430 472170 147498 472226
rect 147554 472170 147622 472226
rect 147678 472170 165250 472226
rect 165306 472170 165374 472226
rect 165430 472170 165498 472226
rect 165554 472170 165622 472226
rect 165678 472170 183250 472226
rect 183306 472170 183374 472226
rect 183430 472170 183498 472226
rect 183554 472170 183622 472226
rect 183678 472170 201250 472226
rect 201306 472170 201374 472226
rect 201430 472170 201498 472226
rect 201554 472170 201622 472226
rect 201678 472170 219250 472226
rect 219306 472170 219374 472226
rect 219430 472170 219498 472226
rect 219554 472170 219622 472226
rect 219678 472170 237250 472226
rect 237306 472170 237374 472226
rect 237430 472170 237498 472226
rect 237554 472170 237622 472226
rect 237678 472170 255250 472226
rect 255306 472170 255374 472226
rect 255430 472170 255498 472226
rect 255554 472170 255622 472226
rect 255678 472170 273250 472226
rect 273306 472170 273374 472226
rect 273430 472170 273498 472226
rect 273554 472170 273622 472226
rect 273678 472170 291250 472226
rect 291306 472170 291374 472226
rect 291430 472170 291498 472226
rect 291554 472170 291622 472226
rect 291678 472170 309250 472226
rect 309306 472170 309374 472226
rect 309430 472170 309498 472226
rect 309554 472170 309622 472226
rect 309678 472170 327250 472226
rect 327306 472170 327374 472226
rect 327430 472170 327498 472226
rect 327554 472170 327622 472226
rect 327678 472170 345250 472226
rect 345306 472170 345374 472226
rect 345430 472170 345498 472226
rect 345554 472170 345622 472226
rect 345678 472170 363250 472226
rect 363306 472170 363374 472226
rect 363430 472170 363498 472226
rect 363554 472170 363622 472226
rect 363678 472170 381250 472226
rect 381306 472170 381374 472226
rect 381430 472170 381498 472226
rect 381554 472170 381622 472226
rect 381678 472170 399250 472226
rect 399306 472170 399374 472226
rect 399430 472170 399498 472226
rect 399554 472170 399622 472226
rect 399678 472170 417250 472226
rect 417306 472170 417374 472226
rect 417430 472170 417498 472226
rect 417554 472170 417622 472226
rect 417678 472170 435250 472226
rect 435306 472170 435374 472226
rect 435430 472170 435498 472226
rect 435554 472170 435622 472226
rect 435678 472170 453250 472226
rect 453306 472170 453374 472226
rect 453430 472170 453498 472226
rect 453554 472170 453622 472226
rect 453678 472170 471250 472226
rect 471306 472170 471374 472226
rect 471430 472170 471498 472226
rect 471554 472170 471622 472226
rect 471678 472170 489250 472226
rect 489306 472170 489374 472226
rect 489430 472170 489498 472226
rect 489554 472170 489622 472226
rect 489678 472170 507250 472226
rect 507306 472170 507374 472226
rect 507430 472170 507498 472226
rect 507554 472170 507622 472226
rect 507678 472170 525250 472226
rect 525306 472170 525374 472226
rect 525430 472170 525498 472226
rect 525554 472170 525622 472226
rect 525678 472170 543250 472226
rect 543306 472170 543374 472226
rect 543430 472170 543498 472226
rect 543554 472170 543622 472226
rect 543678 472170 561250 472226
rect 561306 472170 561374 472226
rect 561430 472170 561498 472226
rect 561554 472170 561622 472226
rect 561678 472170 579250 472226
rect 579306 472170 579374 472226
rect 579430 472170 579498 472226
rect 579554 472170 579622 472226
rect 579678 472170 596496 472226
rect 596552 472170 596620 472226
rect 596676 472170 596744 472226
rect 596800 472170 596868 472226
rect 596924 472170 597980 472226
rect -1916 472102 597980 472170
rect -1916 472046 -860 472102
rect -804 472046 -736 472102
rect -680 472046 -612 472102
rect -556 472046 -488 472102
rect -432 472046 3250 472102
rect 3306 472046 3374 472102
rect 3430 472046 3498 472102
rect 3554 472046 3622 472102
rect 3678 472046 21250 472102
rect 21306 472046 21374 472102
rect 21430 472046 21498 472102
rect 21554 472046 21622 472102
rect 21678 472046 39250 472102
rect 39306 472046 39374 472102
rect 39430 472046 39498 472102
rect 39554 472046 39622 472102
rect 39678 472046 57250 472102
rect 57306 472046 57374 472102
rect 57430 472046 57498 472102
rect 57554 472046 57622 472102
rect 57678 472046 75250 472102
rect 75306 472046 75374 472102
rect 75430 472046 75498 472102
rect 75554 472046 75622 472102
rect 75678 472046 93250 472102
rect 93306 472046 93374 472102
rect 93430 472046 93498 472102
rect 93554 472046 93622 472102
rect 93678 472046 111250 472102
rect 111306 472046 111374 472102
rect 111430 472046 111498 472102
rect 111554 472046 111622 472102
rect 111678 472046 129250 472102
rect 129306 472046 129374 472102
rect 129430 472046 129498 472102
rect 129554 472046 129622 472102
rect 129678 472046 147250 472102
rect 147306 472046 147374 472102
rect 147430 472046 147498 472102
rect 147554 472046 147622 472102
rect 147678 472046 165250 472102
rect 165306 472046 165374 472102
rect 165430 472046 165498 472102
rect 165554 472046 165622 472102
rect 165678 472046 183250 472102
rect 183306 472046 183374 472102
rect 183430 472046 183498 472102
rect 183554 472046 183622 472102
rect 183678 472046 201250 472102
rect 201306 472046 201374 472102
rect 201430 472046 201498 472102
rect 201554 472046 201622 472102
rect 201678 472046 219250 472102
rect 219306 472046 219374 472102
rect 219430 472046 219498 472102
rect 219554 472046 219622 472102
rect 219678 472046 237250 472102
rect 237306 472046 237374 472102
rect 237430 472046 237498 472102
rect 237554 472046 237622 472102
rect 237678 472046 255250 472102
rect 255306 472046 255374 472102
rect 255430 472046 255498 472102
rect 255554 472046 255622 472102
rect 255678 472046 273250 472102
rect 273306 472046 273374 472102
rect 273430 472046 273498 472102
rect 273554 472046 273622 472102
rect 273678 472046 291250 472102
rect 291306 472046 291374 472102
rect 291430 472046 291498 472102
rect 291554 472046 291622 472102
rect 291678 472046 309250 472102
rect 309306 472046 309374 472102
rect 309430 472046 309498 472102
rect 309554 472046 309622 472102
rect 309678 472046 327250 472102
rect 327306 472046 327374 472102
rect 327430 472046 327498 472102
rect 327554 472046 327622 472102
rect 327678 472046 345250 472102
rect 345306 472046 345374 472102
rect 345430 472046 345498 472102
rect 345554 472046 345622 472102
rect 345678 472046 363250 472102
rect 363306 472046 363374 472102
rect 363430 472046 363498 472102
rect 363554 472046 363622 472102
rect 363678 472046 381250 472102
rect 381306 472046 381374 472102
rect 381430 472046 381498 472102
rect 381554 472046 381622 472102
rect 381678 472046 399250 472102
rect 399306 472046 399374 472102
rect 399430 472046 399498 472102
rect 399554 472046 399622 472102
rect 399678 472046 417250 472102
rect 417306 472046 417374 472102
rect 417430 472046 417498 472102
rect 417554 472046 417622 472102
rect 417678 472046 435250 472102
rect 435306 472046 435374 472102
rect 435430 472046 435498 472102
rect 435554 472046 435622 472102
rect 435678 472046 453250 472102
rect 453306 472046 453374 472102
rect 453430 472046 453498 472102
rect 453554 472046 453622 472102
rect 453678 472046 471250 472102
rect 471306 472046 471374 472102
rect 471430 472046 471498 472102
rect 471554 472046 471622 472102
rect 471678 472046 489250 472102
rect 489306 472046 489374 472102
rect 489430 472046 489498 472102
rect 489554 472046 489622 472102
rect 489678 472046 507250 472102
rect 507306 472046 507374 472102
rect 507430 472046 507498 472102
rect 507554 472046 507622 472102
rect 507678 472046 525250 472102
rect 525306 472046 525374 472102
rect 525430 472046 525498 472102
rect 525554 472046 525622 472102
rect 525678 472046 543250 472102
rect 543306 472046 543374 472102
rect 543430 472046 543498 472102
rect 543554 472046 543622 472102
rect 543678 472046 561250 472102
rect 561306 472046 561374 472102
rect 561430 472046 561498 472102
rect 561554 472046 561622 472102
rect 561678 472046 579250 472102
rect 579306 472046 579374 472102
rect 579430 472046 579498 472102
rect 579554 472046 579622 472102
rect 579678 472046 596496 472102
rect 596552 472046 596620 472102
rect 596676 472046 596744 472102
rect 596800 472046 596868 472102
rect 596924 472046 597980 472102
rect -1916 471978 597980 472046
rect -1916 471922 -860 471978
rect -804 471922 -736 471978
rect -680 471922 -612 471978
rect -556 471922 -488 471978
rect -432 471922 3250 471978
rect 3306 471922 3374 471978
rect 3430 471922 3498 471978
rect 3554 471922 3622 471978
rect 3678 471922 21250 471978
rect 21306 471922 21374 471978
rect 21430 471922 21498 471978
rect 21554 471922 21622 471978
rect 21678 471922 39250 471978
rect 39306 471922 39374 471978
rect 39430 471922 39498 471978
rect 39554 471922 39622 471978
rect 39678 471922 57250 471978
rect 57306 471922 57374 471978
rect 57430 471922 57498 471978
rect 57554 471922 57622 471978
rect 57678 471922 75250 471978
rect 75306 471922 75374 471978
rect 75430 471922 75498 471978
rect 75554 471922 75622 471978
rect 75678 471922 93250 471978
rect 93306 471922 93374 471978
rect 93430 471922 93498 471978
rect 93554 471922 93622 471978
rect 93678 471922 111250 471978
rect 111306 471922 111374 471978
rect 111430 471922 111498 471978
rect 111554 471922 111622 471978
rect 111678 471922 129250 471978
rect 129306 471922 129374 471978
rect 129430 471922 129498 471978
rect 129554 471922 129622 471978
rect 129678 471922 147250 471978
rect 147306 471922 147374 471978
rect 147430 471922 147498 471978
rect 147554 471922 147622 471978
rect 147678 471922 165250 471978
rect 165306 471922 165374 471978
rect 165430 471922 165498 471978
rect 165554 471922 165622 471978
rect 165678 471922 183250 471978
rect 183306 471922 183374 471978
rect 183430 471922 183498 471978
rect 183554 471922 183622 471978
rect 183678 471922 201250 471978
rect 201306 471922 201374 471978
rect 201430 471922 201498 471978
rect 201554 471922 201622 471978
rect 201678 471922 219250 471978
rect 219306 471922 219374 471978
rect 219430 471922 219498 471978
rect 219554 471922 219622 471978
rect 219678 471922 237250 471978
rect 237306 471922 237374 471978
rect 237430 471922 237498 471978
rect 237554 471922 237622 471978
rect 237678 471922 255250 471978
rect 255306 471922 255374 471978
rect 255430 471922 255498 471978
rect 255554 471922 255622 471978
rect 255678 471922 273250 471978
rect 273306 471922 273374 471978
rect 273430 471922 273498 471978
rect 273554 471922 273622 471978
rect 273678 471922 291250 471978
rect 291306 471922 291374 471978
rect 291430 471922 291498 471978
rect 291554 471922 291622 471978
rect 291678 471922 309250 471978
rect 309306 471922 309374 471978
rect 309430 471922 309498 471978
rect 309554 471922 309622 471978
rect 309678 471922 327250 471978
rect 327306 471922 327374 471978
rect 327430 471922 327498 471978
rect 327554 471922 327622 471978
rect 327678 471922 345250 471978
rect 345306 471922 345374 471978
rect 345430 471922 345498 471978
rect 345554 471922 345622 471978
rect 345678 471922 363250 471978
rect 363306 471922 363374 471978
rect 363430 471922 363498 471978
rect 363554 471922 363622 471978
rect 363678 471922 381250 471978
rect 381306 471922 381374 471978
rect 381430 471922 381498 471978
rect 381554 471922 381622 471978
rect 381678 471922 399250 471978
rect 399306 471922 399374 471978
rect 399430 471922 399498 471978
rect 399554 471922 399622 471978
rect 399678 471922 417250 471978
rect 417306 471922 417374 471978
rect 417430 471922 417498 471978
rect 417554 471922 417622 471978
rect 417678 471922 435250 471978
rect 435306 471922 435374 471978
rect 435430 471922 435498 471978
rect 435554 471922 435622 471978
rect 435678 471922 453250 471978
rect 453306 471922 453374 471978
rect 453430 471922 453498 471978
rect 453554 471922 453622 471978
rect 453678 471922 471250 471978
rect 471306 471922 471374 471978
rect 471430 471922 471498 471978
rect 471554 471922 471622 471978
rect 471678 471922 489250 471978
rect 489306 471922 489374 471978
rect 489430 471922 489498 471978
rect 489554 471922 489622 471978
rect 489678 471922 507250 471978
rect 507306 471922 507374 471978
rect 507430 471922 507498 471978
rect 507554 471922 507622 471978
rect 507678 471922 525250 471978
rect 525306 471922 525374 471978
rect 525430 471922 525498 471978
rect 525554 471922 525622 471978
rect 525678 471922 543250 471978
rect 543306 471922 543374 471978
rect 543430 471922 543498 471978
rect 543554 471922 543622 471978
rect 543678 471922 561250 471978
rect 561306 471922 561374 471978
rect 561430 471922 561498 471978
rect 561554 471922 561622 471978
rect 561678 471922 579250 471978
rect 579306 471922 579374 471978
rect 579430 471922 579498 471978
rect 579554 471922 579622 471978
rect 579678 471922 596496 471978
rect 596552 471922 596620 471978
rect 596676 471922 596744 471978
rect 596800 471922 596868 471978
rect 596924 471922 597980 471978
rect -1916 471826 597980 471922
rect -1916 460350 597980 460446
rect -1916 460294 -1820 460350
rect -1764 460294 -1696 460350
rect -1640 460294 -1572 460350
rect -1516 460294 -1448 460350
rect -1392 460294 6970 460350
rect 7026 460294 7094 460350
rect 7150 460294 7218 460350
rect 7274 460294 7342 460350
rect 7398 460294 24970 460350
rect 25026 460294 25094 460350
rect 25150 460294 25218 460350
rect 25274 460294 25342 460350
rect 25398 460294 42970 460350
rect 43026 460294 43094 460350
rect 43150 460294 43218 460350
rect 43274 460294 43342 460350
rect 43398 460294 60970 460350
rect 61026 460294 61094 460350
rect 61150 460294 61218 460350
rect 61274 460294 61342 460350
rect 61398 460294 78970 460350
rect 79026 460294 79094 460350
rect 79150 460294 79218 460350
rect 79274 460294 79342 460350
rect 79398 460294 96970 460350
rect 97026 460294 97094 460350
rect 97150 460294 97218 460350
rect 97274 460294 97342 460350
rect 97398 460294 114970 460350
rect 115026 460294 115094 460350
rect 115150 460294 115218 460350
rect 115274 460294 115342 460350
rect 115398 460294 132970 460350
rect 133026 460294 133094 460350
rect 133150 460294 133218 460350
rect 133274 460294 133342 460350
rect 133398 460294 150970 460350
rect 151026 460294 151094 460350
rect 151150 460294 151218 460350
rect 151274 460294 151342 460350
rect 151398 460294 168970 460350
rect 169026 460294 169094 460350
rect 169150 460294 169218 460350
rect 169274 460294 169342 460350
rect 169398 460294 186970 460350
rect 187026 460294 187094 460350
rect 187150 460294 187218 460350
rect 187274 460294 187342 460350
rect 187398 460294 204970 460350
rect 205026 460294 205094 460350
rect 205150 460294 205218 460350
rect 205274 460294 205342 460350
rect 205398 460294 222970 460350
rect 223026 460294 223094 460350
rect 223150 460294 223218 460350
rect 223274 460294 223342 460350
rect 223398 460294 240970 460350
rect 241026 460294 241094 460350
rect 241150 460294 241218 460350
rect 241274 460294 241342 460350
rect 241398 460294 258970 460350
rect 259026 460294 259094 460350
rect 259150 460294 259218 460350
rect 259274 460294 259342 460350
rect 259398 460294 276970 460350
rect 277026 460294 277094 460350
rect 277150 460294 277218 460350
rect 277274 460294 277342 460350
rect 277398 460294 294970 460350
rect 295026 460294 295094 460350
rect 295150 460294 295218 460350
rect 295274 460294 295342 460350
rect 295398 460294 312970 460350
rect 313026 460294 313094 460350
rect 313150 460294 313218 460350
rect 313274 460294 313342 460350
rect 313398 460294 330970 460350
rect 331026 460294 331094 460350
rect 331150 460294 331218 460350
rect 331274 460294 331342 460350
rect 331398 460294 348970 460350
rect 349026 460294 349094 460350
rect 349150 460294 349218 460350
rect 349274 460294 349342 460350
rect 349398 460294 366970 460350
rect 367026 460294 367094 460350
rect 367150 460294 367218 460350
rect 367274 460294 367342 460350
rect 367398 460294 384970 460350
rect 385026 460294 385094 460350
rect 385150 460294 385218 460350
rect 385274 460294 385342 460350
rect 385398 460294 402970 460350
rect 403026 460294 403094 460350
rect 403150 460294 403218 460350
rect 403274 460294 403342 460350
rect 403398 460294 420970 460350
rect 421026 460294 421094 460350
rect 421150 460294 421218 460350
rect 421274 460294 421342 460350
rect 421398 460294 438970 460350
rect 439026 460294 439094 460350
rect 439150 460294 439218 460350
rect 439274 460294 439342 460350
rect 439398 460294 456970 460350
rect 457026 460294 457094 460350
rect 457150 460294 457218 460350
rect 457274 460294 457342 460350
rect 457398 460294 474970 460350
rect 475026 460294 475094 460350
rect 475150 460294 475218 460350
rect 475274 460294 475342 460350
rect 475398 460294 492970 460350
rect 493026 460294 493094 460350
rect 493150 460294 493218 460350
rect 493274 460294 493342 460350
rect 493398 460294 510970 460350
rect 511026 460294 511094 460350
rect 511150 460294 511218 460350
rect 511274 460294 511342 460350
rect 511398 460294 528970 460350
rect 529026 460294 529094 460350
rect 529150 460294 529218 460350
rect 529274 460294 529342 460350
rect 529398 460294 546970 460350
rect 547026 460294 547094 460350
rect 547150 460294 547218 460350
rect 547274 460294 547342 460350
rect 547398 460294 564970 460350
rect 565026 460294 565094 460350
rect 565150 460294 565218 460350
rect 565274 460294 565342 460350
rect 565398 460294 582970 460350
rect 583026 460294 583094 460350
rect 583150 460294 583218 460350
rect 583274 460294 583342 460350
rect 583398 460294 597456 460350
rect 597512 460294 597580 460350
rect 597636 460294 597704 460350
rect 597760 460294 597828 460350
rect 597884 460294 597980 460350
rect -1916 460226 597980 460294
rect -1916 460170 -1820 460226
rect -1764 460170 -1696 460226
rect -1640 460170 -1572 460226
rect -1516 460170 -1448 460226
rect -1392 460170 6970 460226
rect 7026 460170 7094 460226
rect 7150 460170 7218 460226
rect 7274 460170 7342 460226
rect 7398 460170 24970 460226
rect 25026 460170 25094 460226
rect 25150 460170 25218 460226
rect 25274 460170 25342 460226
rect 25398 460170 42970 460226
rect 43026 460170 43094 460226
rect 43150 460170 43218 460226
rect 43274 460170 43342 460226
rect 43398 460170 60970 460226
rect 61026 460170 61094 460226
rect 61150 460170 61218 460226
rect 61274 460170 61342 460226
rect 61398 460170 78970 460226
rect 79026 460170 79094 460226
rect 79150 460170 79218 460226
rect 79274 460170 79342 460226
rect 79398 460170 96970 460226
rect 97026 460170 97094 460226
rect 97150 460170 97218 460226
rect 97274 460170 97342 460226
rect 97398 460170 114970 460226
rect 115026 460170 115094 460226
rect 115150 460170 115218 460226
rect 115274 460170 115342 460226
rect 115398 460170 132970 460226
rect 133026 460170 133094 460226
rect 133150 460170 133218 460226
rect 133274 460170 133342 460226
rect 133398 460170 150970 460226
rect 151026 460170 151094 460226
rect 151150 460170 151218 460226
rect 151274 460170 151342 460226
rect 151398 460170 168970 460226
rect 169026 460170 169094 460226
rect 169150 460170 169218 460226
rect 169274 460170 169342 460226
rect 169398 460170 186970 460226
rect 187026 460170 187094 460226
rect 187150 460170 187218 460226
rect 187274 460170 187342 460226
rect 187398 460170 204970 460226
rect 205026 460170 205094 460226
rect 205150 460170 205218 460226
rect 205274 460170 205342 460226
rect 205398 460170 222970 460226
rect 223026 460170 223094 460226
rect 223150 460170 223218 460226
rect 223274 460170 223342 460226
rect 223398 460170 240970 460226
rect 241026 460170 241094 460226
rect 241150 460170 241218 460226
rect 241274 460170 241342 460226
rect 241398 460170 258970 460226
rect 259026 460170 259094 460226
rect 259150 460170 259218 460226
rect 259274 460170 259342 460226
rect 259398 460170 276970 460226
rect 277026 460170 277094 460226
rect 277150 460170 277218 460226
rect 277274 460170 277342 460226
rect 277398 460170 294970 460226
rect 295026 460170 295094 460226
rect 295150 460170 295218 460226
rect 295274 460170 295342 460226
rect 295398 460170 312970 460226
rect 313026 460170 313094 460226
rect 313150 460170 313218 460226
rect 313274 460170 313342 460226
rect 313398 460170 330970 460226
rect 331026 460170 331094 460226
rect 331150 460170 331218 460226
rect 331274 460170 331342 460226
rect 331398 460170 348970 460226
rect 349026 460170 349094 460226
rect 349150 460170 349218 460226
rect 349274 460170 349342 460226
rect 349398 460170 366970 460226
rect 367026 460170 367094 460226
rect 367150 460170 367218 460226
rect 367274 460170 367342 460226
rect 367398 460170 384970 460226
rect 385026 460170 385094 460226
rect 385150 460170 385218 460226
rect 385274 460170 385342 460226
rect 385398 460170 402970 460226
rect 403026 460170 403094 460226
rect 403150 460170 403218 460226
rect 403274 460170 403342 460226
rect 403398 460170 420970 460226
rect 421026 460170 421094 460226
rect 421150 460170 421218 460226
rect 421274 460170 421342 460226
rect 421398 460170 438970 460226
rect 439026 460170 439094 460226
rect 439150 460170 439218 460226
rect 439274 460170 439342 460226
rect 439398 460170 456970 460226
rect 457026 460170 457094 460226
rect 457150 460170 457218 460226
rect 457274 460170 457342 460226
rect 457398 460170 474970 460226
rect 475026 460170 475094 460226
rect 475150 460170 475218 460226
rect 475274 460170 475342 460226
rect 475398 460170 492970 460226
rect 493026 460170 493094 460226
rect 493150 460170 493218 460226
rect 493274 460170 493342 460226
rect 493398 460170 510970 460226
rect 511026 460170 511094 460226
rect 511150 460170 511218 460226
rect 511274 460170 511342 460226
rect 511398 460170 528970 460226
rect 529026 460170 529094 460226
rect 529150 460170 529218 460226
rect 529274 460170 529342 460226
rect 529398 460170 546970 460226
rect 547026 460170 547094 460226
rect 547150 460170 547218 460226
rect 547274 460170 547342 460226
rect 547398 460170 564970 460226
rect 565026 460170 565094 460226
rect 565150 460170 565218 460226
rect 565274 460170 565342 460226
rect 565398 460170 582970 460226
rect 583026 460170 583094 460226
rect 583150 460170 583218 460226
rect 583274 460170 583342 460226
rect 583398 460170 597456 460226
rect 597512 460170 597580 460226
rect 597636 460170 597704 460226
rect 597760 460170 597828 460226
rect 597884 460170 597980 460226
rect -1916 460102 597980 460170
rect -1916 460046 -1820 460102
rect -1764 460046 -1696 460102
rect -1640 460046 -1572 460102
rect -1516 460046 -1448 460102
rect -1392 460046 6970 460102
rect 7026 460046 7094 460102
rect 7150 460046 7218 460102
rect 7274 460046 7342 460102
rect 7398 460046 24970 460102
rect 25026 460046 25094 460102
rect 25150 460046 25218 460102
rect 25274 460046 25342 460102
rect 25398 460046 42970 460102
rect 43026 460046 43094 460102
rect 43150 460046 43218 460102
rect 43274 460046 43342 460102
rect 43398 460046 60970 460102
rect 61026 460046 61094 460102
rect 61150 460046 61218 460102
rect 61274 460046 61342 460102
rect 61398 460046 78970 460102
rect 79026 460046 79094 460102
rect 79150 460046 79218 460102
rect 79274 460046 79342 460102
rect 79398 460046 96970 460102
rect 97026 460046 97094 460102
rect 97150 460046 97218 460102
rect 97274 460046 97342 460102
rect 97398 460046 114970 460102
rect 115026 460046 115094 460102
rect 115150 460046 115218 460102
rect 115274 460046 115342 460102
rect 115398 460046 132970 460102
rect 133026 460046 133094 460102
rect 133150 460046 133218 460102
rect 133274 460046 133342 460102
rect 133398 460046 150970 460102
rect 151026 460046 151094 460102
rect 151150 460046 151218 460102
rect 151274 460046 151342 460102
rect 151398 460046 168970 460102
rect 169026 460046 169094 460102
rect 169150 460046 169218 460102
rect 169274 460046 169342 460102
rect 169398 460046 186970 460102
rect 187026 460046 187094 460102
rect 187150 460046 187218 460102
rect 187274 460046 187342 460102
rect 187398 460046 204970 460102
rect 205026 460046 205094 460102
rect 205150 460046 205218 460102
rect 205274 460046 205342 460102
rect 205398 460046 222970 460102
rect 223026 460046 223094 460102
rect 223150 460046 223218 460102
rect 223274 460046 223342 460102
rect 223398 460046 240970 460102
rect 241026 460046 241094 460102
rect 241150 460046 241218 460102
rect 241274 460046 241342 460102
rect 241398 460046 258970 460102
rect 259026 460046 259094 460102
rect 259150 460046 259218 460102
rect 259274 460046 259342 460102
rect 259398 460046 276970 460102
rect 277026 460046 277094 460102
rect 277150 460046 277218 460102
rect 277274 460046 277342 460102
rect 277398 460046 294970 460102
rect 295026 460046 295094 460102
rect 295150 460046 295218 460102
rect 295274 460046 295342 460102
rect 295398 460046 312970 460102
rect 313026 460046 313094 460102
rect 313150 460046 313218 460102
rect 313274 460046 313342 460102
rect 313398 460046 330970 460102
rect 331026 460046 331094 460102
rect 331150 460046 331218 460102
rect 331274 460046 331342 460102
rect 331398 460046 348970 460102
rect 349026 460046 349094 460102
rect 349150 460046 349218 460102
rect 349274 460046 349342 460102
rect 349398 460046 366970 460102
rect 367026 460046 367094 460102
rect 367150 460046 367218 460102
rect 367274 460046 367342 460102
rect 367398 460046 384970 460102
rect 385026 460046 385094 460102
rect 385150 460046 385218 460102
rect 385274 460046 385342 460102
rect 385398 460046 402970 460102
rect 403026 460046 403094 460102
rect 403150 460046 403218 460102
rect 403274 460046 403342 460102
rect 403398 460046 420970 460102
rect 421026 460046 421094 460102
rect 421150 460046 421218 460102
rect 421274 460046 421342 460102
rect 421398 460046 438970 460102
rect 439026 460046 439094 460102
rect 439150 460046 439218 460102
rect 439274 460046 439342 460102
rect 439398 460046 456970 460102
rect 457026 460046 457094 460102
rect 457150 460046 457218 460102
rect 457274 460046 457342 460102
rect 457398 460046 474970 460102
rect 475026 460046 475094 460102
rect 475150 460046 475218 460102
rect 475274 460046 475342 460102
rect 475398 460046 492970 460102
rect 493026 460046 493094 460102
rect 493150 460046 493218 460102
rect 493274 460046 493342 460102
rect 493398 460046 510970 460102
rect 511026 460046 511094 460102
rect 511150 460046 511218 460102
rect 511274 460046 511342 460102
rect 511398 460046 528970 460102
rect 529026 460046 529094 460102
rect 529150 460046 529218 460102
rect 529274 460046 529342 460102
rect 529398 460046 546970 460102
rect 547026 460046 547094 460102
rect 547150 460046 547218 460102
rect 547274 460046 547342 460102
rect 547398 460046 564970 460102
rect 565026 460046 565094 460102
rect 565150 460046 565218 460102
rect 565274 460046 565342 460102
rect 565398 460046 582970 460102
rect 583026 460046 583094 460102
rect 583150 460046 583218 460102
rect 583274 460046 583342 460102
rect 583398 460046 597456 460102
rect 597512 460046 597580 460102
rect 597636 460046 597704 460102
rect 597760 460046 597828 460102
rect 597884 460046 597980 460102
rect -1916 459978 597980 460046
rect -1916 459922 -1820 459978
rect -1764 459922 -1696 459978
rect -1640 459922 -1572 459978
rect -1516 459922 -1448 459978
rect -1392 459922 6970 459978
rect 7026 459922 7094 459978
rect 7150 459922 7218 459978
rect 7274 459922 7342 459978
rect 7398 459922 24970 459978
rect 25026 459922 25094 459978
rect 25150 459922 25218 459978
rect 25274 459922 25342 459978
rect 25398 459922 42970 459978
rect 43026 459922 43094 459978
rect 43150 459922 43218 459978
rect 43274 459922 43342 459978
rect 43398 459922 60970 459978
rect 61026 459922 61094 459978
rect 61150 459922 61218 459978
rect 61274 459922 61342 459978
rect 61398 459922 78970 459978
rect 79026 459922 79094 459978
rect 79150 459922 79218 459978
rect 79274 459922 79342 459978
rect 79398 459922 96970 459978
rect 97026 459922 97094 459978
rect 97150 459922 97218 459978
rect 97274 459922 97342 459978
rect 97398 459922 114970 459978
rect 115026 459922 115094 459978
rect 115150 459922 115218 459978
rect 115274 459922 115342 459978
rect 115398 459922 132970 459978
rect 133026 459922 133094 459978
rect 133150 459922 133218 459978
rect 133274 459922 133342 459978
rect 133398 459922 150970 459978
rect 151026 459922 151094 459978
rect 151150 459922 151218 459978
rect 151274 459922 151342 459978
rect 151398 459922 168970 459978
rect 169026 459922 169094 459978
rect 169150 459922 169218 459978
rect 169274 459922 169342 459978
rect 169398 459922 186970 459978
rect 187026 459922 187094 459978
rect 187150 459922 187218 459978
rect 187274 459922 187342 459978
rect 187398 459922 204970 459978
rect 205026 459922 205094 459978
rect 205150 459922 205218 459978
rect 205274 459922 205342 459978
rect 205398 459922 222970 459978
rect 223026 459922 223094 459978
rect 223150 459922 223218 459978
rect 223274 459922 223342 459978
rect 223398 459922 240970 459978
rect 241026 459922 241094 459978
rect 241150 459922 241218 459978
rect 241274 459922 241342 459978
rect 241398 459922 258970 459978
rect 259026 459922 259094 459978
rect 259150 459922 259218 459978
rect 259274 459922 259342 459978
rect 259398 459922 276970 459978
rect 277026 459922 277094 459978
rect 277150 459922 277218 459978
rect 277274 459922 277342 459978
rect 277398 459922 294970 459978
rect 295026 459922 295094 459978
rect 295150 459922 295218 459978
rect 295274 459922 295342 459978
rect 295398 459922 312970 459978
rect 313026 459922 313094 459978
rect 313150 459922 313218 459978
rect 313274 459922 313342 459978
rect 313398 459922 330970 459978
rect 331026 459922 331094 459978
rect 331150 459922 331218 459978
rect 331274 459922 331342 459978
rect 331398 459922 348970 459978
rect 349026 459922 349094 459978
rect 349150 459922 349218 459978
rect 349274 459922 349342 459978
rect 349398 459922 366970 459978
rect 367026 459922 367094 459978
rect 367150 459922 367218 459978
rect 367274 459922 367342 459978
rect 367398 459922 384970 459978
rect 385026 459922 385094 459978
rect 385150 459922 385218 459978
rect 385274 459922 385342 459978
rect 385398 459922 402970 459978
rect 403026 459922 403094 459978
rect 403150 459922 403218 459978
rect 403274 459922 403342 459978
rect 403398 459922 420970 459978
rect 421026 459922 421094 459978
rect 421150 459922 421218 459978
rect 421274 459922 421342 459978
rect 421398 459922 438970 459978
rect 439026 459922 439094 459978
rect 439150 459922 439218 459978
rect 439274 459922 439342 459978
rect 439398 459922 456970 459978
rect 457026 459922 457094 459978
rect 457150 459922 457218 459978
rect 457274 459922 457342 459978
rect 457398 459922 474970 459978
rect 475026 459922 475094 459978
rect 475150 459922 475218 459978
rect 475274 459922 475342 459978
rect 475398 459922 492970 459978
rect 493026 459922 493094 459978
rect 493150 459922 493218 459978
rect 493274 459922 493342 459978
rect 493398 459922 510970 459978
rect 511026 459922 511094 459978
rect 511150 459922 511218 459978
rect 511274 459922 511342 459978
rect 511398 459922 528970 459978
rect 529026 459922 529094 459978
rect 529150 459922 529218 459978
rect 529274 459922 529342 459978
rect 529398 459922 546970 459978
rect 547026 459922 547094 459978
rect 547150 459922 547218 459978
rect 547274 459922 547342 459978
rect 547398 459922 564970 459978
rect 565026 459922 565094 459978
rect 565150 459922 565218 459978
rect 565274 459922 565342 459978
rect 565398 459922 582970 459978
rect 583026 459922 583094 459978
rect 583150 459922 583218 459978
rect 583274 459922 583342 459978
rect 583398 459922 597456 459978
rect 597512 459922 597580 459978
rect 597636 459922 597704 459978
rect 597760 459922 597828 459978
rect 597884 459922 597980 459978
rect -1916 459826 597980 459922
rect -1916 454350 597980 454446
rect -1916 454294 -860 454350
rect -804 454294 -736 454350
rect -680 454294 -612 454350
rect -556 454294 -488 454350
rect -432 454294 3250 454350
rect 3306 454294 3374 454350
rect 3430 454294 3498 454350
rect 3554 454294 3622 454350
rect 3678 454294 201250 454350
rect 201306 454294 201374 454350
rect 201430 454294 201498 454350
rect 201554 454294 201622 454350
rect 201678 454294 381250 454350
rect 381306 454294 381374 454350
rect 381430 454294 381498 454350
rect 381554 454294 381622 454350
rect 381678 454294 399250 454350
rect 399306 454294 399374 454350
rect 399430 454294 399498 454350
rect 399554 454294 399622 454350
rect 399678 454294 579250 454350
rect 579306 454294 579374 454350
rect 579430 454294 579498 454350
rect 579554 454294 579622 454350
rect 579678 454294 596496 454350
rect 596552 454294 596620 454350
rect 596676 454294 596744 454350
rect 596800 454294 596868 454350
rect 596924 454294 597980 454350
rect -1916 454226 597980 454294
rect -1916 454170 -860 454226
rect -804 454170 -736 454226
rect -680 454170 -612 454226
rect -556 454170 -488 454226
rect -432 454170 3250 454226
rect 3306 454170 3374 454226
rect 3430 454170 3498 454226
rect 3554 454170 3622 454226
rect 3678 454170 201250 454226
rect 201306 454170 201374 454226
rect 201430 454170 201498 454226
rect 201554 454170 201622 454226
rect 201678 454170 381250 454226
rect 381306 454170 381374 454226
rect 381430 454170 381498 454226
rect 381554 454170 381622 454226
rect 381678 454170 399250 454226
rect 399306 454170 399374 454226
rect 399430 454170 399498 454226
rect 399554 454170 399622 454226
rect 399678 454170 579250 454226
rect 579306 454170 579374 454226
rect 579430 454170 579498 454226
rect 579554 454170 579622 454226
rect 579678 454170 596496 454226
rect 596552 454170 596620 454226
rect 596676 454170 596744 454226
rect 596800 454170 596868 454226
rect 596924 454170 597980 454226
rect -1916 454102 597980 454170
rect -1916 454046 -860 454102
rect -804 454046 -736 454102
rect -680 454046 -612 454102
rect -556 454046 -488 454102
rect -432 454046 3250 454102
rect 3306 454046 3374 454102
rect 3430 454046 3498 454102
rect 3554 454046 3622 454102
rect 3678 454046 201250 454102
rect 201306 454046 201374 454102
rect 201430 454046 201498 454102
rect 201554 454046 201622 454102
rect 201678 454046 381250 454102
rect 381306 454046 381374 454102
rect 381430 454046 381498 454102
rect 381554 454046 381622 454102
rect 381678 454046 399250 454102
rect 399306 454046 399374 454102
rect 399430 454046 399498 454102
rect 399554 454046 399622 454102
rect 399678 454046 579250 454102
rect 579306 454046 579374 454102
rect 579430 454046 579498 454102
rect 579554 454046 579622 454102
rect 579678 454046 596496 454102
rect 596552 454046 596620 454102
rect 596676 454046 596744 454102
rect 596800 454046 596868 454102
rect 596924 454046 597980 454102
rect -1916 453978 597980 454046
rect -1916 453922 -860 453978
rect -804 453922 -736 453978
rect -680 453922 -612 453978
rect -556 453922 -488 453978
rect -432 453922 3250 453978
rect 3306 453922 3374 453978
rect 3430 453922 3498 453978
rect 3554 453922 3622 453978
rect 3678 453922 201250 453978
rect 201306 453922 201374 453978
rect 201430 453922 201498 453978
rect 201554 453922 201622 453978
rect 201678 453922 381250 453978
rect 381306 453922 381374 453978
rect 381430 453922 381498 453978
rect 381554 453922 381622 453978
rect 381678 453922 399250 453978
rect 399306 453922 399374 453978
rect 399430 453922 399498 453978
rect 399554 453922 399622 453978
rect 399678 453922 579250 453978
rect 579306 453922 579374 453978
rect 579430 453922 579498 453978
rect 579554 453922 579622 453978
rect 579678 453922 596496 453978
rect 596552 453922 596620 453978
rect 596676 453922 596744 453978
rect 596800 453922 596868 453978
rect 596924 453922 597980 453978
rect -1916 453826 597980 453922
rect -1916 442350 597980 442446
rect -1916 442294 -1820 442350
rect -1764 442294 -1696 442350
rect -1640 442294 -1572 442350
rect -1516 442294 -1448 442350
rect -1392 442294 6970 442350
rect 7026 442294 7094 442350
rect 7150 442294 7218 442350
rect 7274 442294 7342 442350
rect 7398 442294 204970 442350
rect 205026 442294 205094 442350
rect 205150 442294 205218 442350
rect 205274 442294 205342 442350
rect 205398 442294 384970 442350
rect 385026 442294 385094 442350
rect 385150 442294 385218 442350
rect 385274 442294 385342 442350
rect 385398 442294 402970 442350
rect 403026 442294 403094 442350
rect 403150 442294 403218 442350
rect 403274 442294 403342 442350
rect 403398 442294 582970 442350
rect 583026 442294 583094 442350
rect 583150 442294 583218 442350
rect 583274 442294 583342 442350
rect 583398 442294 597456 442350
rect 597512 442294 597580 442350
rect 597636 442294 597704 442350
rect 597760 442294 597828 442350
rect 597884 442294 597980 442350
rect -1916 442226 597980 442294
rect -1916 442170 -1820 442226
rect -1764 442170 -1696 442226
rect -1640 442170 -1572 442226
rect -1516 442170 -1448 442226
rect -1392 442170 6970 442226
rect 7026 442170 7094 442226
rect 7150 442170 7218 442226
rect 7274 442170 7342 442226
rect 7398 442170 204970 442226
rect 205026 442170 205094 442226
rect 205150 442170 205218 442226
rect 205274 442170 205342 442226
rect 205398 442170 384970 442226
rect 385026 442170 385094 442226
rect 385150 442170 385218 442226
rect 385274 442170 385342 442226
rect 385398 442170 402970 442226
rect 403026 442170 403094 442226
rect 403150 442170 403218 442226
rect 403274 442170 403342 442226
rect 403398 442170 582970 442226
rect 583026 442170 583094 442226
rect 583150 442170 583218 442226
rect 583274 442170 583342 442226
rect 583398 442170 597456 442226
rect 597512 442170 597580 442226
rect 597636 442170 597704 442226
rect 597760 442170 597828 442226
rect 597884 442170 597980 442226
rect -1916 442102 597980 442170
rect -1916 442046 -1820 442102
rect -1764 442046 -1696 442102
rect -1640 442046 -1572 442102
rect -1516 442046 -1448 442102
rect -1392 442046 6970 442102
rect 7026 442046 7094 442102
rect 7150 442046 7218 442102
rect 7274 442046 7342 442102
rect 7398 442046 204970 442102
rect 205026 442046 205094 442102
rect 205150 442046 205218 442102
rect 205274 442046 205342 442102
rect 205398 442046 384970 442102
rect 385026 442046 385094 442102
rect 385150 442046 385218 442102
rect 385274 442046 385342 442102
rect 385398 442046 402970 442102
rect 403026 442046 403094 442102
rect 403150 442046 403218 442102
rect 403274 442046 403342 442102
rect 403398 442046 582970 442102
rect 583026 442046 583094 442102
rect 583150 442046 583218 442102
rect 583274 442046 583342 442102
rect 583398 442046 597456 442102
rect 597512 442046 597580 442102
rect 597636 442046 597704 442102
rect 597760 442046 597828 442102
rect 597884 442046 597980 442102
rect -1916 441978 597980 442046
rect -1916 441922 -1820 441978
rect -1764 441922 -1696 441978
rect -1640 441922 -1572 441978
rect -1516 441922 -1448 441978
rect -1392 441922 6970 441978
rect 7026 441922 7094 441978
rect 7150 441922 7218 441978
rect 7274 441922 7342 441978
rect 7398 441922 204970 441978
rect 205026 441922 205094 441978
rect 205150 441922 205218 441978
rect 205274 441922 205342 441978
rect 205398 441922 384970 441978
rect 385026 441922 385094 441978
rect 385150 441922 385218 441978
rect 385274 441922 385342 441978
rect 385398 441922 402970 441978
rect 403026 441922 403094 441978
rect 403150 441922 403218 441978
rect 403274 441922 403342 441978
rect 403398 441922 582970 441978
rect 583026 441922 583094 441978
rect 583150 441922 583218 441978
rect 583274 441922 583342 441978
rect 583398 441922 597456 441978
rect 597512 441922 597580 441978
rect 597636 441922 597704 441978
rect 597760 441922 597828 441978
rect 597884 441922 597980 441978
rect -1916 441826 597980 441922
rect -1916 436350 597980 436446
rect -1916 436294 -860 436350
rect -804 436294 -736 436350
rect -680 436294 -612 436350
rect -556 436294 -488 436350
rect -432 436294 3250 436350
rect 3306 436294 3374 436350
rect 3430 436294 3498 436350
rect 3554 436294 3622 436350
rect 3678 436294 201250 436350
rect 201306 436294 201374 436350
rect 201430 436294 201498 436350
rect 201554 436294 201622 436350
rect 201678 436294 381250 436350
rect 381306 436294 381374 436350
rect 381430 436294 381498 436350
rect 381554 436294 381622 436350
rect 381678 436294 399250 436350
rect 399306 436294 399374 436350
rect 399430 436294 399498 436350
rect 399554 436294 399622 436350
rect 399678 436294 579250 436350
rect 579306 436294 579374 436350
rect 579430 436294 579498 436350
rect 579554 436294 579622 436350
rect 579678 436294 596496 436350
rect 596552 436294 596620 436350
rect 596676 436294 596744 436350
rect 596800 436294 596868 436350
rect 596924 436294 597980 436350
rect -1916 436226 597980 436294
rect -1916 436170 -860 436226
rect -804 436170 -736 436226
rect -680 436170 -612 436226
rect -556 436170 -488 436226
rect -432 436170 3250 436226
rect 3306 436170 3374 436226
rect 3430 436170 3498 436226
rect 3554 436170 3622 436226
rect 3678 436170 201250 436226
rect 201306 436170 201374 436226
rect 201430 436170 201498 436226
rect 201554 436170 201622 436226
rect 201678 436170 381250 436226
rect 381306 436170 381374 436226
rect 381430 436170 381498 436226
rect 381554 436170 381622 436226
rect 381678 436170 399250 436226
rect 399306 436170 399374 436226
rect 399430 436170 399498 436226
rect 399554 436170 399622 436226
rect 399678 436170 579250 436226
rect 579306 436170 579374 436226
rect 579430 436170 579498 436226
rect 579554 436170 579622 436226
rect 579678 436170 596496 436226
rect 596552 436170 596620 436226
rect 596676 436170 596744 436226
rect 596800 436170 596868 436226
rect 596924 436170 597980 436226
rect -1916 436102 597980 436170
rect -1916 436046 -860 436102
rect -804 436046 -736 436102
rect -680 436046 -612 436102
rect -556 436046 -488 436102
rect -432 436046 3250 436102
rect 3306 436046 3374 436102
rect 3430 436046 3498 436102
rect 3554 436046 3622 436102
rect 3678 436046 201250 436102
rect 201306 436046 201374 436102
rect 201430 436046 201498 436102
rect 201554 436046 201622 436102
rect 201678 436046 381250 436102
rect 381306 436046 381374 436102
rect 381430 436046 381498 436102
rect 381554 436046 381622 436102
rect 381678 436046 399250 436102
rect 399306 436046 399374 436102
rect 399430 436046 399498 436102
rect 399554 436046 399622 436102
rect 399678 436046 579250 436102
rect 579306 436046 579374 436102
rect 579430 436046 579498 436102
rect 579554 436046 579622 436102
rect 579678 436046 596496 436102
rect 596552 436046 596620 436102
rect 596676 436046 596744 436102
rect 596800 436046 596868 436102
rect 596924 436046 597980 436102
rect -1916 435978 597980 436046
rect -1916 435922 -860 435978
rect -804 435922 -736 435978
rect -680 435922 -612 435978
rect -556 435922 -488 435978
rect -432 435922 3250 435978
rect 3306 435922 3374 435978
rect 3430 435922 3498 435978
rect 3554 435922 3622 435978
rect 3678 435922 201250 435978
rect 201306 435922 201374 435978
rect 201430 435922 201498 435978
rect 201554 435922 201622 435978
rect 201678 435922 381250 435978
rect 381306 435922 381374 435978
rect 381430 435922 381498 435978
rect 381554 435922 381622 435978
rect 381678 435922 399250 435978
rect 399306 435922 399374 435978
rect 399430 435922 399498 435978
rect 399554 435922 399622 435978
rect 399678 435922 579250 435978
rect 579306 435922 579374 435978
rect 579430 435922 579498 435978
rect 579554 435922 579622 435978
rect 579678 435922 596496 435978
rect 596552 435922 596620 435978
rect 596676 435922 596744 435978
rect 596800 435922 596868 435978
rect 596924 435922 597980 435978
rect -1916 435826 597980 435922
rect -1916 424350 597980 424446
rect -1916 424294 -1820 424350
rect -1764 424294 -1696 424350
rect -1640 424294 -1572 424350
rect -1516 424294 -1448 424350
rect -1392 424294 6970 424350
rect 7026 424294 7094 424350
rect 7150 424294 7218 424350
rect 7274 424294 7342 424350
rect 7398 424294 204970 424350
rect 205026 424294 205094 424350
rect 205150 424294 205218 424350
rect 205274 424294 205342 424350
rect 205398 424294 384970 424350
rect 385026 424294 385094 424350
rect 385150 424294 385218 424350
rect 385274 424294 385342 424350
rect 385398 424294 402970 424350
rect 403026 424294 403094 424350
rect 403150 424294 403218 424350
rect 403274 424294 403342 424350
rect 403398 424294 582970 424350
rect 583026 424294 583094 424350
rect 583150 424294 583218 424350
rect 583274 424294 583342 424350
rect 583398 424294 597456 424350
rect 597512 424294 597580 424350
rect 597636 424294 597704 424350
rect 597760 424294 597828 424350
rect 597884 424294 597980 424350
rect -1916 424226 597980 424294
rect -1916 424170 -1820 424226
rect -1764 424170 -1696 424226
rect -1640 424170 -1572 424226
rect -1516 424170 -1448 424226
rect -1392 424170 6970 424226
rect 7026 424170 7094 424226
rect 7150 424170 7218 424226
rect 7274 424170 7342 424226
rect 7398 424170 204970 424226
rect 205026 424170 205094 424226
rect 205150 424170 205218 424226
rect 205274 424170 205342 424226
rect 205398 424170 384970 424226
rect 385026 424170 385094 424226
rect 385150 424170 385218 424226
rect 385274 424170 385342 424226
rect 385398 424170 402970 424226
rect 403026 424170 403094 424226
rect 403150 424170 403218 424226
rect 403274 424170 403342 424226
rect 403398 424170 582970 424226
rect 583026 424170 583094 424226
rect 583150 424170 583218 424226
rect 583274 424170 583342 424226
rect 583398 424170 597456 424226
rect 597512 424170 597580 424226
rect 597636 424170 597704 424226
rect 597760 424170 597828 424226
rect 597884 424170 597980 424226
rect -1916 424102 597980 424170
rect -1916 424046 -1820 424102
rect -1764 424046 -1696 424102
rect -1640 424046 -1572 424102
rect -1516 424046 -1448 424102
rect -1392 424046 6970 424102
rect 7026 424046 7094 424102
rect 7150 424046 7218 424102
rect 7274 424046 7342 424102
rect 7398 424046 204970 424102
rect 205026 424046 205094 424102
rect 205150 424046 205218 424102
rect 205274 424046 205342 424102
rect 205398 424046 384970 424102
rect 385026 424046 385094 424102
rect 385150 424046 385218 424102
rect 385274 424046 385342 424102
rect 385398 424046 402970 424102
rect 403026 424046 403094 424102
rect 403150 424046 403218 424102
rect 403274 424046 403342 424102
rect 403398 424046 582970 424102
rect 583026 424046 583094 424102
rect 583150 424046 583218 424102
rect 583274 424046 583342 424102
rect 583398 424046 597456 424102
rect 597512 424046 597580 424102
rect 597636 424046 597704 424102
rect 597760 424046 597828 424102
rect 597884 424046 597980 424102
rect -1916 423978 597980 424046
rect -1916 423922 -1820 423978
rect -1764 423922 -1696 423978
rect -1640 423922 -1572 423978
rect -1516 423922 -1448 423978
rect -1392 423922 6970 423978
rect 7026 423922 7094 423978
rect 7150 423922 7218 423978
rect 7274 423922 7342 423978
rect 7398 423922 204970 423978
rect 205026 423922 205094 423978
rect 205150 423922 205218 423978
rect 205274 423922 205342 423978
rect 205398 423922 384970 423978
rect 385026 423922 385094 423978
rect 385150 423922 385218 423978
rect 385274 423922 385342 423978
rect 385398 423922 402970 423978
rect 403026 423922 403094 423978
rect 403150 423922 403218 423978
rect 403274 423922 403342 423978
rect 403398 423922 582970 423978
rect 583026 423922 583094 423978
rect 583150 423922 583218 423978
rect 583274 423922 583342 423978
rect 583398 423922 597456 423978
rect 597512 423922 597580 423978
rect 597636 423922 597704 423978
rect 597760 423922 597828 423978
rect 597884 423922 597980 423978
rect -1916 423826 597980 423922
rect -1916 418350 597980 418446
rect -1916 418294 -860 418350
rect -804 418294 -736 418350
rect -680 418294 -612 418350
rect -556 418294 -488 418350
rect -432 418294 3250 418350
rect 3306 418294 3374 418350
rect 3430 418294 3498 418350
rect 3554 418294 3622 418350
rect 3678 418294 201250 418350
rect 201306 418294 201374 418350
rect 201430 418294 201498 418350
rect 201554 418294 201622 418350
rect 201678 418294 381250 418350
rect 381306 418294 381374 418350
rect 381430 418294 381498 418350
rect 381554 418294 381622 418350
rect 381678 418294 399250 418350
rect 399306 418294 399374 418350
rect 399430 418294 399498 418350
rect 399554 418294 399622 418350
rect 399678 418294 579250 418350
rect 579306 418294 579374 418350
rect 579430 418294 579498 418350
rect 579554 418294 579622 418350
rect 579678 418294 596496 418350
rect 596552 418294 596620 418350
rect 596676 418294 596744 418350
rect 596800 418294 596868 418350
rect 596924 418294 597980 418350
rect -1916 418226 597980 418294
rect -1916 418170 -860 418226
rect -804 418170 -736 418226
rect -680 418170 -612 418226
rect -556 418170 -488 418226
rect -432 418170 3250 418226
rect 3306 418170 3374 418226
rect 3430 418170 3498 418226
rect 3554 418170 3622 418226
rect 3678 418170 201250 418226
rect 201306 418170 201374 418226
rect 201430 418170 201498 418226
rect 201554 418170 201622 418226
rect 201678 418170 381250 418226
rect 381306 418170 381374 418226
rect 381430 418170 381498 418226
rect 381554 418170 381622 418226
rect 381678 418170 399250 418226
rect 399306 418170 399374 418226
rect 399430 418170 399498 418226
rect 399554 418170 399622 418226
rect 399678 418170 579250 418226
rect 579306 418170 579374 418226
rect 579430 418170 579498 418226
rect 579554 418170 579622 418226
rect 579678 418170 596496 418226
rect 596552 418170 596620 418226
rect 596676 418170 596744 418226
rect 596800 418170 596868 418226
rect 596924 418170 597980 418226
rect -1916 418102 597980 418170
rect -1916 418046 -860 418102
rect -804 418046 -736 418102
rect -680 418046 -612 418102
rect -556 418046 -488 418102
rect -432 418046 3250 418102
rect 3306 418046 3374 418102
rect 3430 418046 3498 418102
rect 3554 418046 3622 418102
rect 3678 418046 201250 418102
rect 201306 418046 201374 418102
rect 201430 418046 201498 418102
rect 201554 418046 201622 418102
rect 201678 418046 381250 418102
rect 381306 418046 381374 418102
rect 381430 418046 381498 418102
rect 381554 418046 381622 418102
rect 381678 418046 399250 418102
rect 399306 418046 399374 418102
rect 399430 418046 399498 418102
rect 399554 418046 399622 418102
rect 399678 418046 579250 418102
rect 579306 418046 579374 418102
rect 579430 418046 579498 418102
rect 579554 418046 579622 418102
rect 579678 418046 596496 418102
rect 596552 418046 596620 418102
rect 596676 418046 596744 418102
rect 596800 418046 596868 418102
rect 596924 418046 597980 418102
rect -1916 417978 597980 418046
rect -1916 417922 -860 417978
rect -804 417922 -736 417978
rect -680 417922 -612 417978
rect -556 417922 -488 417978
rect -432 417922 3250 417978
rect 3306 417922 3374 417978
rect 3430 417922 3498 417978
rect 3554 417922 3622 417978
rect 3678 417922 201250 417978
rect 201306 417922 201374 417978
rect 201430 417922 201498 417978
rect 201554 417922 201622 417978
rect 201678 417922 381250 417978
rect 381306 417922 381374 417978
rect 381430 417922 381498 417978
rect 381554 417922 381622 417978
rect 381678 417922 399250 417978
rect 399306 417922 399374 417978
rect 399430 417922 399498 417978
rect 399554 417922 399622 417978
rect 399678 417922 579250 417978
rect 579306 417922 579374 417978
rect 579430 417922 579498 417978
rect 579554 417922 579622 417978
rect 579678 417922 596496 417978
rect 596552 417922 596620 417978
rect 596676 417922 596744 417978
rect 596800 417922 596868 417978
rect 596924 417922 597980 417978
rect -1916 417826 597980 417922
rect -1916 406350 597980 406446
rect -1916 406294 -1820 406350
rect -1764 406294 -1696 406350
rect -1640 406294 -1572 406350
rect -1516 406294 -1448 406350
rect -1392 406294 6970 406350
rect 7026 406294 7094 406350
rect 7150 406294 7218 406350
rect 7274 406294 7342 406350
rect 7398 406294 204970 406350
rect 205026 406294 205094 406350
rect 205150 406294 205218 406350
rect 205274 406294 205342 406350
rect 205398 406294 384970 406350
rect 385026 406294 385094 406350
rect 385150 406294 385218 406350
rect 385274 406294 385342 406350
rect 385398 406294 402970 406350
rect 403026 406294 403094 406350
rect 403150 406294 403218 406350
rect 403274 406294 403342 406350
rect 403398 406294 582970 406350
rect 583026 406294 583094 406350
rect 583150 406294 583218 406350
rect 583274 406294 583342 406350
rect 583398 406294 597456 406350
rect 597512 406294 597580 406350
rect 597636 406294 597704 406350
rect 597760 406294 597828 406350
rect 597884 406294 597980 406350
rect -1916 406226 597980 406294
rect -1916 406170 -1820 406226
rect -1764 406170 -1696 406226
rect -1640 406170 -1572 406226
rect -1516 406170 -1448 406226
rect -1392 406170 6970 406226
rect 7026 406170 7094 406226
rect 7150 406170 7218 406226
rect 7274 406170 7342 406226
rect 7398 406170 204970 406226
rect 205026 406170 205094 406226
rect 205150 406170 205218 406226
rect 205274 406170 205342 406226
rect 205398 406170 384970 406226
rect 385026 406170 385094 406226
rect 385150 406170 385218 406226
rect 385274 406170 385342 406226
rect 385398 406170 402970 406226
rect 403026 406170 403094 406226
rect 403150 406170 403218 406226
rect 403274 406170 403342 406226
rect 403398 406170 582970 406226
rect 583026 406170 583094 406226
rect 583150 406170 583218 406226
rect 583274 406170 583342 406226
rect 583398 406170 597456 406226
rect 597512 406170 597580 406226
rect 597636 406170 597704 406226
rect 597760 406170 597828 406226
rect 597884 406170 597980 406226
rect -1916 406102 597980 406170
rect -1916 406046 -1820 406102
rect -1764 406046 -1696 406102
rect -1640 406046 -1572 406102
rect -1516 406046 -1448 406102
rect -1392 406046 6970 406102
rect 7026 406046 7094 406102
rect 7150 406046 7218 406102
rect 7274 406046 7342 406102
rect 7398 406046 204970 406102
rect 205026 406046 205094 406102
rect 205150 406046 205218 406102
rect 205274 406046 205342 406102
rect 205398 406046 384970 406102
rect 385026 406046 385094 406102
rect 385150 406046 385218 406102
rect 385274 406046 385342 406102
rect 385398 406046 402970 406102
rect 403026 406046 403094 406102
rect 403150 406046 403218 406102
rect 403274 406046 403342 406102
rect 403398 406046 582970 406102
rect 583026 406046 583094 406102
rect 583150 406046 583218 406102
rect 583274 406046 583342 406102
rect 583398 406046 597456 406102
rect 597512 406046 597580 406102
rect 597636 406046 597704 406102
rect 597760 406046 597828 406102
rect 597884 406046 597980 406102
rect -1916 405978 597980 406046
rect -1916 405922 -1820 405978
rect -1764 405922 -1696 405978
rect -1640 405922 -1572 405978
rect -1516 405922 -1448 405978
rect -1392 405922 6970 405978
rect 7026 405922 7094 405978
rect 7150 405922 7218 405978
rect 7274 405922 7342 405978
rect 7398 405922 204970 405978
rect 205026 405922 205094 405978
rect 205150 405922 205218 405978
rect 205274 405922 205342 405978
rect 205398 405922 384970 405978
rect 385026 405922 385094 405978
rect 385150 405922 385218 405978
rect 385274 405922 385342 405978
rect 385398 405922 402970 405978
rect 403026 405922 403094 405978
rect 403150 405922 403218 405978
rect 403274 405922 403342 405978
rect 403398 405922 582970 405978
rect 583026 405922 583094 405978
rect 583150 405922 583218 405978
rect 583274 405922 583342 405978
rect 583398 405922 597456 405978
rect 597512 405922 597580 405978
rect 597636 405922 597704 405978
rect 597760 405922 597828 405978
rect 597884 405922 597980 405978
rect -1916 405826 597980 405922
rect -1916 400350 597980 400446
rect -1916 400294 -860 400350
rect -804 400294 -736 400350
rect -680 400294 -612 400350
rect -556 400294 -488 400350
rect -432 400294 3250 400350
rect 3306 400294 3374 400350
rect 3430 400294 3498 400350
rect 3554 400294 3622 400350
rect 3678 400294 201250 400350
rect 201306 400294 201374 400350
rect 201430 400294 201498 400350
rect 201554 400294 201622 400350
rect 201678 400294 381250 400350
rect 381306 400294 381374 400350
rect 381430 400294 381498 400350
rect 381554 400294 381622 400350
rect 381678 400294 399250 400350
rect 399306 400294 399374 400350
rect 399430 400294 399498 400350
rect 399554 400294 399622 400350
rect 399678 400294 579250 400350
rect 579306 400294 579374 400350
rect 579430 400294 579498 400350
rect 579554 400294 579622 400350
rect 579678 400294 596496 400350
rect 596552 400294 596620 400350
rect 596676 400294 596744 400350
rect 596800 400294 596868 400350
rect 596924 400294 597980 400350
rect -1916 400226 597980 400294
rect -1916 400170 -860 400226
rect -804 400170 -736 400226
rect -680 400170 -612 400226
rect -556 400170 -488 400226
rect -432 400170 3250 400226
rect 3306 400170 3374 400226
rect 3430 400170 3498 400226
rect 3554 400170 3622 400226
rect 3678 400170 201250 400226
rect 201306 400170 201374 400226
rect 201430 400170 201498 400226
rect 201554 400170 201622 400226
rect 201678 400170 381250 400226
rect 381306 400170 381374 400226
rect 381430 400170 381498 400226
rect 381554 400170 381622 400226
rect 381678 400170 399250 400226
rect 399306 400170 399374 400226
rect 399430 400170 399498 400226
rect 399554 400170 399622 400226
rect 399678 400170 579250 400226
rect 579306 400170 579374 400226
rect 579430 400170 579498 400226
rect 579554 400170 579622 400226
rect 579678 400170 596496 400226
rect 596552 400170 596620 400226
rect 596676 400170 596744 400226
rect 596800 400170 596868 400226
rect 596924 400170 597980 400226
rect -1916 400102 597980 400170
rect -1916 400046 -860 400102
rect -804 400046 -736 400102
rect -680 400046 -612 400102
rect -556 400046 -488 400102
rect -432 400046 3250 400102
rect 3306 400046 3374 400102
rect 3430 400046 3498 400102
rect 3554 400046 3622 400102
rect 3678 400046 201250 400102
rect 201306 400046 201374 400102
rect 201430 400046 201498 400102
rect 201554 400046 201622 400102
rect 201678 400046 381250 400102
rect 381306 400046 381374 400102
rect 381430 400046 381498 400102
rect 381554 400046 381622 400102
rect 381678 400046 399250 400102
rect 399306 400046 399374 400102
rect 399430 400046 399498 400102
rect 399554 400046 399622 400102
rect 399678 400046 579250 400102
rect 579306 400046 579374 400102
rect 579430 400046 579498 400102
rect 579554 400046 579622 400102
rect 579678 400046 596496 400102
rect 596552 400046 596620 400102
rect 596676 400046 596744 400102
rect 596800 400046 596868 400102
rect 596924 400046 597980 400102
rect -1916 399978 597980 400046
rect -1916 399922 -860 399978
rect -804 399922 -736 399978
rect -680 399922 -612 399978
rect -556 399922 -488 399978
rect -432 399922 3250 399978
rect 3306 399922 3374 399978
rect 3430 399922 3498 399978
rect 3554 399922 3622 399978
rect 3678 399922 201250 399978
rect 201306 399922 201374 399978
rect 201430 399922 201498 399978
rect 201554 399922 201622 399978
rect 201678 399922 381250 399978
rect 381306 399922 381374 399978
rect 381430 399922 381498 399978
rect 381554 399922 381622 399978
rect 381678 399922 399250 399978
rect 399306 399922 399374 399978
rect 399430 399922 399498 399978
rect 399554 399922 399622 399978
rect 399678 399922 579250 399978
rect 579306 399922 579374 399978
rect 579430 399922 579498 399978
rect 579554 399922 579622 399978
rect 579678 399922 596496 399978
rect 596552 399922 596620 399978
rect 596676 399922 596744 399978
rect 596800 399922 596868 399978
rect 596924 399922 597980 399978
rect -1916 399826 597980 399922
rect -1916 388350 597980 388446
rect -1916 388294 -1820 388350
rect -1764 388294 -1696 388350
rect -1640 388294 -1572 388350
rect -1516 388294 -1448 388350
rect -1392 388294 6970 388350
rect 7026 388294 7094 388350
rect 7150 388294 7218 388350
rect 7274 388294 7342 388350
rect 7398 388294 204970 388350
rect 205026 388294 205094 388350
rect 205150 388294 205218 388350
rect 205274 388294 205342 388350
rect 205398 388294 384970 388350
rect 385026 388294 385094 388350
rect 385150 388294 385218 388350
rect 385274 388294 385342 388350
rect 385398 388294 402970 388350
rect 403026 388294 403094 388350
rect 403150 388294 403218 388350
rect 403274 388294 403342 388350
rect 403398 388294 582970 388350
rect 583026 388294 583094 388350
rect 583150 388294 583218 388350
rect 583274 388294 583342 388350
rect 583398 388294 597456 388350
rect 597512 388294 597580 388350
rect 597636 388294 597704 388350
rect 597760 388294 597828 388350
rect 597884 388294 597980 388350
rect -1916 388226 597980 388294
rect -1916 388170 -1820 388226
rect -1764 388170 -1696 388226
rect -1640 388170 -1572 388226
rect -1516 388170 -1448 388226
rect -1392 388170 6970 388226
rect 7026 388170 7094 388226
rect 7150 388170 7218 388226
rect 7274 388170 7342 388226
rect 7398 388170 204970 388226
rect 205026 388170 205094 388226
rect 205150 388170 205218 388226
rect 205274 388170 205342 388226
rect 205398 388170 384970 388226
rect 385026 388170 385094 388226
rect 385150 388170 385218 388226
rect 385274 388170 385342 388226
rect 385398 388170 402970 388226
rect 403026 388170 403094 388226
rect 403150 388170 403218 388226
rect 403274 388170 403342 388226
rect 403398 388170 582970 388226
rect 583026 388170 583094 388226
rect 583150 388170 583218 388226
rect 583274 388170 583342 388226
rect 583398 388170 597456 388226
rect 597512 388170 597580 388226
rect 597636 388170 597704 388226
rect 597760 388170 597828 388226
rect 597884 388170 597980 388226
rect -1916 388102 597980 388170
rect -1916 388046 -1820 388102
rect -1764 388046 -1696 388102
rect -1640 388046 -1572 388102
rect -1516 388046 -1448 388102
rect -1392 388046 6970 388102
rect 7026 388046 7094 388102
rect 7150 388046 7218 388102
rect 7274 388046 7342 388102
rect 7398 388046 204970 388102
rect 205026 388046 205094 388102
rect 205150 388046 205218 388102
rect 205274 388046 205342 388102
rect 205398 388046 384970 388102
rect 385026 388046 385094 388102
rect 385150 388046 385218 388102
rect 385274 388046 385342 388102
rect 385398 388046 402970 388102
rect 403026 388046 403094 388102
rect 403150 388046 403218 388102
rect 403274 388046 403342 388102
rect 403398 388046 582970 388102
rect 583026 388046 583094 388102
rect 583150 388046 583218 388102
rect 583274 388046 583342 388102
rect 583398 388046 597456 388102
rect 597512 388046 597580 388102
rect 597636 388046 597704 388102
rect 597760 388046 597828 388102
rect 597884 388046 597980 388102
rect -1916 387978 597980 388046
rect -1916 387922 -1820 387978
rect -1764 387922 -1696 387978
rect -1640 387922 -1572 387978
rect -1516 387922 -1448 387978
rect -1392 387922 6970 387978
rect 7026 387922 7094 387978
rect 7150 387922 7218 387978
rect 7274 387922 7342 387978
rect 7398 387922 204970 387978
rect 205026 387922 205094 387978
rect 205150 387922 205218 387978
rect 205274 387922 205342 387978
rect 205398 387922 384970 387978
rect 385026 387922 385094 387978
rect 385150 387922 385218 387978
rect 385274 387922 385342 387978
rect 385398 387922 402970 387978
rect 403026 387922 403094 387978
rect 403150 387922 403218 387978
rect 403274 387922 403342 387978
rect 403398 387922 582970 387978
rect 583026 387922 583094 387978
rect 583150 387922 583218 387978
rect 583274 387922 583342 387978
rect 583398 387922 597456 387978
rect 597512 387922 597580 387978
rect 597636 387922 597704 387978
rect 597760 387922 597828 387978
rect 597884 387922 597980 387978
rect -1916 387826 597980 387922
rect -1916 382350 597980 382446
rect -1916 382294 -860 382350
rect -804 382294 -736 382350
rect -680 382294 -612 382350
rect -556 382294 -488 382350
rect -432 382294 3250 382350
rect 3306 382294 3374 382350
rect 3430 382294 3498 382350
rect 3554 382294 3622 382350
rect 3678 382294 201250 382350
rect 201306 382294 201374 382350
rect 201430 382294 201498 382350
rect 201554 382294 201622 382350
rect 201678 382294 381250 382350
rect 381306 382294 381374 382350
rect 381430 382294 381498 382350
rect 381554 382294 381622 382350
rect 381678 382294 399250 382350
rect 399306 382294 399374 382350
rect 399430 382294 399498 382350
rect 399554 382294 399622 382350
rect 399678 382294 579250 382350
rect 579306 382294 579374 382350
rect 579430 382294 579498 382350
rect 579554 382294 579622 382350
rect 579678 382294 596496 382350
rect 596552 382294 596620 382350
rect 596676 382294 596744 382350
rect 596800 382294 596868 382350
rect 596924 382294 597980 382350
rect -1916 382226 597980 382294
rect -1916 382170 -860 382226
rect -804 382170 -736 382226
rect -680 382170 -612 382226
rect -556 382170 -488 382226
rect -432 382170 3250 382226
rect 3306 382170 3374 382226
rect 3430 382170 3498 382226
rect 3554 382170 3622 382226
rect 3678 382170 201250 382226
rect 201306 382170 201374 382226
rect 201430 382170 201498 382226
rect 201554 382170 201622 382226
rect 201678 382170 381250 382226
rect 381306 382170 381374 382226
rect 381430 382170 381498 382226
rect 381554 382170 381622 382226
rect 381678 382170 399250 382226
rect 399306 382170 399374 382226
rect 399430 382170 399498 382226
rect 399554 382170 399622 382226
rect 399678 382170 579250 382226
rect 579306 382170 579374 382226
rect 579430 382170 579498 382226
rect 579554 382170 579622 382226
rect 579678 382170 596496 382226
rect 596552 382170 596620 382226
rect 596676 382170 596744 382226
rect 596800 382170 596868 382226
rect 596924 382170 597980 382226
rect -1916 382102 597980 382170
rect -1916 382046 -860 382102
rect -804 382046 -736 382102
rect -680 382046 -612 382102
rect -556 382046 -488 382102
rect -432 382046 3250 382102
rect 3306 382046 3374 382102
rect 3430 382046 3498 382102
rect 3554 382046 3622 382102
rect 3678 382046 201250 382102
rect 201306 382046 201374 382102
rect 201430 382046 201498 382102
rect 201554 382046 201622 382102
rect 201678 382046 381250 382102
rect 381306 382046 381374 382102
rect 381430 382046 381498 382102
rect 381554 382046 381622 382102
rect 381678 382046 399250 382102
rect 399306 382046 399374 382102
rect 399430 382046 399498 382102
rect 399554 382046 399622 382102
rect 399678 382046 579250 382102
rect 579306 382046 579374 382102
rect 579430 382046 579498 382102
rect 579554 382046 579622 382102
rect 579678 382046 596496 382102
rect 596552 382046 596620 382102
rect 596676 382046 596744 382102
rect 596800 382046 596868 382102
rect 596924 382046 597980 382102
rect -1916 381978 597980 382046
rect -1916 381922 -860 381978
rect -804 381922 -736 381978
rect -680 381922 -612 381978
rect -556 381922 -488 381978
rect -432 381922 3250 381978
rect 3306 381922 3374 381978
rect 3430 381922 3498 381978
rect 3554 381922 3622 381978
rect 3678 381922 201250 381978
rect 201306 381922 201374 381978
rect 201430 381922 201498 381978
rect 201554 381922 201622 381978
rect 201678 381922 381250 381978
rect 381306 381922 381374 381978
rect 381430 381922 381498 381978
rect 381554 381922 381622 381978
rect 381678 381922 399250 381978
rect 399306 381922 399374 381978
rect 399430 381922 399498 381978
rect 399554 381922 399622 381978
rect 399678 381922 579250 381978
rect 579306 381922 579374 381978
rect 579430 381922 579498 381978
rect 579554 381922 579622 381978
rect 579678 381922 596496 381978
rect 596552 381922 596620 381978
rect 596676 381922 596744 381978
rect 596800 381922 596868 381978
rect 596924 381922 597980 381978
rect -1916 381826 597980 381922
rect -1916 370350 597980 370446
rect -1916 370294 -1820 370350
rect -1764 370294 -1696 370350
rect -1640 370294 -1572 370350
rect -1516 370294 -1448 370350
rect -1392 370294 6970 370350
rect 7026 370294 7094 370350
rect 7150 370294 7218 370350
rect 7274 370294 7342 370350
rect 7398 370294 204970 370350
rect 205026 370294 205094 370350
rect 205150 370294 205218 370350
rect 205274 370294 205342 370350
rect 205398 370294 384970 370350
rect 385026 370294 385094 370350
rect 385150 370294 385218 370350
rect 385274 370294 385342 370350
rect 385398 370294 402970 370350
rect 403026 370294 403094 370350
rect 403150 370294 403218 370350
rect 403274 370294 403342 370350
rect 403398 370294 582970 370350
rect 583026 370294 583094 370350
rect 583150 370294 583218 370350
rect 583274 370294 583342 370350
rect 583398 370294 597456 370350
rect 597512 370294 597580 370350
rect 597636 370294 597704 370350
rect 597760 370294 597828 370350
rect 597884 370294 597980 370350
rect -1916 370226 597980 370294
rect -1916 370170 -1820 370226
rect -1764 370170 -1696 370226
rect -1640 370170 -1572 370226
rect -1516 370170 -1448 370226
rect -1392 370170 6970 370226
rect 7026 370170 7094 370226
rect 7150 370170 7218 370226
rect 7274 370170 7342 370226
rect 7398 370170 204970 370226
rect 205026 370170 205094 370226
rect 205150 370170 205218 370226
rect 205274 370170 205342 370226
rect 205398 370170 384970 370226
rect 385026 370170 385094 370226
rect 385150 370170 385218 370226
rect 385274 370170 385342 370226
rect 385398 370170 402970 370226
rect 403026 370170 403094 370226
rect 403150 370170 403218 370226
rect 403274 370170 403342 370226
rect 403398 370170 582970 370226
rect 583026 370170 583094 370226
rect 583150 370170 583218 370226
rect 583274 370170 583342 370226
rect 583398 370170 597456 370226
rect 597512 370170 597580 370226
rect 597636 370170 597704 370226
rect 597760 370170 597828 370226
rect 597884 370170 597980 370226
rect -1916 370102 597980 370170
rect -1916 370046 -1820 370102
rect -1764 370046 -1696 370102
rect -1640 370046 -1572 370102
rect -1516 370046 -1448 370102
rect -1392 370046 6970 370102
rect 7026 370046 7094 370102
rect 7150 370046 7218 370102
rect 7274 370046 7342 370102
rect 7398 370046 204970 370102
rect 205026 370046 205094 370102
rect 205150 370046 205218 370102
rect 205274 370046 205342 370102
rect 205398 370046 384970 370102
rect 385026 370046 385094 370102
rect 385150 370046 385218 370102
rect 385274 370046 385342 370102
rect 385398 370046 402970 370102
rect 403026 370046 403094 370102
rect 403150 370046 403218 370102
rect 403274 370046 403342 370102
rect 403398 370046 582970 370102
rect 583026 370046 583094 370102
rect 583150 370046 583218 370102
rect 583274 370046 583342 370102
rect 583398 370046 597456 370102
rect 597512 370046 597580 370102
rect 597636 370046 597704 370102
rect 597760 370046 597828 370102
rect 597884 370046 597980 370102
rect -1916 369978 597980 370046
rect -1916 369922 -1820 369978
rect -1764 369922 -1696 369978
rect -1640 369922 -1572 369978
rect -1516 369922 -1448 369978
rect -1392 369922 6970 369978
rect 7026 369922 7094 369978
rect 7150 369922 7218 369978
rect 7274 369922 7342 369978
rect 7398 369922 204970 369978
rect 205026 369922 205094 369978
rect 205150 369922 205218 369978
rect 205274 369922 205342 369978
rect 205398 369922 384970 369978
rect 385026 369922 385094 369978
rect 385150 369922 385218 369978
rect 385274 369922 385342 369978
rect 385398 369922 402970 369978
rect 403026 369922 403094 369978
rect 403150 369922 403218 369978
rect 403274 369922 403342 369978
rect 403398 369922 582970 369978
rect 583026 369922 583094 369978
rect 583150 369922 583218 369978
rect 583274 369922 583342 369978
rect 583398 369922 597456 369978
rect 597512 369922 597580 369978
rect 597636 369922 597704 369978
rect 597760 369922 597828 369978
rect 597884 369922 597980 369978
rect -1916 369826 597980 369922
rect -1916 364350 597980 364446
rect -1916 364294 -860 364350
rect -804 364294 -736 364350
rect -680 364294 -612 364350
rect -556 364294 -488 364350
rect -432 364294 3250 364350
rect 3306 364294 3374 364350
rect 3430 364294 3498 364350
rect 3554 364294 3622 364350
rect 3678 364294 201250 364350
rect 201306 364294 201374 364350
rect 201430 364294 201498 364350
rect 201554 364294 201622 364350
rect 201678 364294 381250 364350
rect 381306 364294 381374 364350
rect 381430 364294 381498 364350
rect 381554 364294 381622 364350
rect 381678 364294 399250 364350
rect 399306 364294 399374 364350
rect 399430 364294 399498 364350
rect 399554 364294 399622 364350
rect 399678 364294 579250 364350
rect 579306 364294 579374 364350
rect 579430 364294 579498 364350
rect 579554 364294 579622 364350
rect 579678 364294 596496 364350
rect 596552 364294 596620 364350
rect 596676 364294 596744 364350
rect 596800 364294 596868 364350
rect 596924 364294 597980 364350
rect -1916 364226 597980 364294
rect -1916 364170 -860 364226
rect -804 364170 -736 364226
rect -680 364170 -612 364226
rect -556 364170 -488 364226
rect -432 364170 3250 364226
rect 3306 364170 3374 364226
rect 3430 364170 3498 364226
rect 3554 364170 3622 364226
rect 3678 364170 201250 364226
rect 201306 364170 201374 364226
rect 201430 364170 201498 364226
rect 201554 364170 201622 364226
rect 201678 364170 381250 364226
rect 381306 364170 381374 364226
rect 381430 364170 381498 364226
rect 381554 364170 381622 364226
rect 381678 364170 399250 364226
rect 399306 364170 399374 364226
rect 399430 364170 399498 364226
rect 399554 364170 399622 364226
rect 399678 364170 579250 364226
rect 579306 364170 579374 364226
rect 579430 364170 579498 364226
rect 579554 364170 579622 364226
rect 579678 364170 596496 364226
rect 596552 364170 596620 364226
rect 596676 364170 596744 364226
rect 596800 364170 596868 364226
rect 596924 364170 597980 364226
rect -1916 364102 597980 364170
rect -1916 364046 -860 364102
rect -804 364046 -736 364102
rect -680 364046 -612 364102
rect -556 364046 -488 364102
rect -432 364046 3250 364102
rect 3306 364046 3374 364102
rect 3430 364046 3498 364102
rect 3554 364046 3622 364102
rect 3678 364046 201250 364102
rect 201306 364046 201374 364102
rect 201430 364046 201498 364102
rect 201554 364046 201622 364102
rect 201678 364046 381250 364102
rect 381306 364046 381374 364102
rect 381430 364046 381498 364102
rect 381554 364046 381622 364102
rect 381678 364046 399250 364102
rect 399306 364046 399374 364102
rect 399430 364046 399498 364102
rect 399554 364046 399622 364102
rect 399678 364046 579250 364102
rect 579306 364046 579374 364102
rect 579430 364046 579498 364102
rect 579554 364046 579622 364102
rect 579678 364046 596496 364102
rect 596552 364046 596620 364102
rect 596676 364046 596744 364102
rect 596800 364046 596868 364102
rect 596924 364046 597980 364102
rect -1916 363978 597980 364046
rect -1916 363922 -860 363978
rect -804 363922 -736 363978
rect -680 363922 -612 363978
rect -556 363922 -488 363978
rect -432 363922 3250 363978
rect 3306 363922 3374 363978
rect 3430 363922 3498 363978
rect 3554 363922 3622 363978
rect 3678 363922 201250 363978
rect 201306 363922 201374 363978
rect 201430 363922 201498 363978
rect 201554 363922 201622 363978
rect 201678 363922 381250 363978
rect 381306 363922 381374 363978
rect 381430 363922 381498 363978
rect 381554 363922 381622 363978
rect 381678 363922 399250 363978
rect 399306 363922 399374 363978
rect 399430 363922 399498 363978
rect 399554 363922 399622 363978
rect 399678 363922 579250 363978
rect 579306 363922 579374 363978
rect 579430 363922 579498 363978
rect 579554 363922 579622 363978
rect 579678 363922 596496 363978
rect 596552 363922 596620 363978
rect 596676 363922 596744 363978
rect 596800 363922 596868 363978
rect 596924 363922 597980 363978
rect -1916 363826 597980 363922
rect -1916 352350 597980 352446
rect -1916 352294 -1820 352350
rect -1764 352294 -1696 352350
rect -1640 352294 -1572 352350
rect -1516 352294 -1448 352350
rect -1392 352294 6970 352350
rect 7026 352294 7094 352350
rect 7150 352294 7218 352350
rect 7274 352294 7342 352350
rect 7398 352294 204970 352350
rect 205026 352294 205094 352350
rect 205150 352294 205218 352350
rect 205274 352294 205342 352350
rect 205398 352294 384970 352350
rect 385026 352294 385094 352350
rect 385150 352294 385218 352350
rect 385274 352294 385342 352350
rect 385398 352294 402970 352350
rect 403026 352294 403094 352350
rect 403150 352294 403218 352350
rect 403274 352294 403342 352350
rect 403398 352294 582970 352350
rect 583026 352294 583094 352350
rect 583150 352294 583218 352350
rect 583274 352294 583342 352350
rect 583398 352294 597456 352350
rect 597512 352294 597580 352350
rect 597636 352294 597704 352350
rect 597760 352294 597828 352350
rect 597884 352294 597980 352350
rect -1916 352226 597980 352294
rect -1916 352170 -1820 352226
rect -1764 352170 -1696 352226
rect -1640 352170 -1572 352226
rect -1516 352170 -1448 352226
rect -1392 352170 6970 352226
rect 7026 352170 7094 352226
rect 7150 352170 7218 352226
rect 7274 352170 7342 352226
rect 7398 352170 204970 352226
rect 205026 352170 205094 352226
rect 205150 352170 205218 352226
rect 205274 352170 205342 352226
rect 205398 352170 384970 352226
rect 385026 352170 385094 352226
rect 385150 352170 385218 352226
rect 385274 352170 385342 352226
rect 385398 352170 402970 352226
rect 403026 352170 403094 352226
rect 403150 352170 403218 352226
rect 403274 352170 403342 352226
rect 403398 352170 582970 352226
rect 583026 352170 583094 352226
rect 583150 352170 583218 352226
rect 583274 352170 583342 352226
rect 583398 352170 597456 352226
rect 597512 352170 597580 352226
rect 597636 352170 597704 352226
rect 597760 352170 597828 352226
rect 597884 352170 597980 352226
rect -1916 352102 597980 352170
rect -1916 352046 -1820 352102
rect -1764 352046 -1696 352102
rect -1640 352046 -1572 352102
rect -1516 352046 -1448 352102
rect -1392 352046 6970 352102
rect 7026 352046 7094 352102
rect 7150 352046 7218 352102
rect 7274 352046 7342 352102
rect 7398 352046 204970 352102
rect 205026 352046 205094 352102
rect 205150 352046 205218 352102
rect 205274 352046 205342 352102
rect 205398 352046 384970 352102
rect 385026 352046 385094 352102
rect 385150 352046 385218 352102
rect 385274 352046 385342 352102
rect 385398 352046 402970 352102
rect 403026 352046 403094 352102
rect 403150 352046 403218 352102
rect 403274 352046 403342 352102
rect 403398 352046 582970 352102
rect 583026 352046 583094 352102
rect 583150 352046 583218 352102
rect 583274 352046 583342 352102
rect 583398 352046 597456 352102
rect 597512 352046 597580 352102
rect 597636 352046 597704 352102
rect 597760 352046 597828 352102
rect 597884 352046 597980 352102
rect -1916 351978 597980 352046
rect -1916 351922 -1820 351978
rect -1764 351922 -1696 351978
rect -1640 351922 -1572 351978
rect -1516 351922 -1448 351978
rect -1392 351922 6970 351978
rect 7026 351922 7094 351978
rect 7150 351922 7218 351978
rect 7274 351922 7342 351978
rect 7398 351922 204970 351978
rect 205026 351922 205094 351978
rect 205150 351922 205218 351978
rect 205274 351922 205342 351978
rect 205398 351922 384970 351978
rect 385026 351922 385094 351978
rect 385150 351922 385218 351978
rect 385274 351922 385342 351978
rect 385398 351922 402970 351978
rect 403026 351922 403094 351978
rect 403150 351922 403218 351978
rect 403274 351922 403342 351978
rect 403398 351922 582970 351978
rect 583026 351922 583094 351978
rect 583150 351922 583218 351978
rect 583274 351922 583342 351978
rect 583398 351922 597456 351978
rect 597512 351922 597580 351978
rect 597636 351922 597704 351978
rect 597760 351922 597828 351978
rect 597884 351922 597980 351978
rect -1916 351826 597980 351922
rect -1916 346350 597980 346446
rect -1916 346294 -860 346350
rect -804 346294 -736 346350
rect -680 346294 -612 346350
rect -556 346294 -488 346350
rect -432 346294 3250 346350
rect 3306 346294 3374 346350
rect 3430 346294 3498 346350
rect 3554 346294 3622 346350
rect 3678 346294 201250 346350
rect 201306 346294 201374 346350
rect 201430 346294 201498 346350
rect 201554 346294 201622 346350
rect 201678 346294 381250 346350
rect 381306 346294 381374 346350
rect 381430 346294 381498 346350
rect 381554 346294 381622 346350
rect 381678 346294 399250 346350
rect 399306 346294 399374 346350
rect 399430 346294 399498 346350
rect 399554 346294 399622 346350
rect 399678 346294 579250 346350
rect 579306 346294 579374 346350
rect 579430 346294 579498 346350
rect 579554 346294 579622 346350
rect 579678 346294 596496 346350
rect 596552 346294 596620 346350
rect 596676 346294 596744 346350
rect 596800 346294 596868 346350
rect 596924 346294 597980 346350
rect -1916 346226 597980 346294
rect -1916 346170 -860 346226
rect -804 346170 -736 346226
rect -680 346170 -612 346226
rect -556 346170 -488 346226
rect -432 346170 3250 346226
rect 3306 346170 3374 346226
rect 3430 346170 3498 346226
rect 3554 346170 3622 346226
rect 3678 346170 201250 346226
rect 201306 346170 201374 346226
rect 201430 346170 201498 346226
rect 201554 346170 201622 346226
rect 201678 346170 381250 346226
rect 381306 346170 381374 346226
rect 381430 346170 381498 346226
rect 381554 346170 381622 346226
rect 381678 346170 399250 346226
rect 399306 346170 399374 346226
rect 399430 346170 399498 346226
rect 399554 346170 399622 346226
rect 399678 346170 579250 346226
rect 579306 346170 579374 346226
rect 579430 346170 579498 346226
rect 579554 346170 579622 346226
rect 579678 346170 596496 346226
rect 596552 346170 596620 346226
rect 596676 346170 596744 346226
rect 596800 346170 596868 346226
rect 596924 346170 597980 346226
rect -1916 346102 597980 346170
rect -1916 346046 -860 346102
rect -804 346046 -736 346102
rect -680 346046 -612 346102
rect -556 346046 -488 346102
rect -432 346046 3250 346102
rect 3306 346046 3374 346102
rect 3430 346046 3498 346102
rect 3554 346046 3622 346102
rect 3678 346046 201250 346102
rect 201306 346046 201374 346102
rect 201430 346046 201498 346102
rect 201554 346046 201622 346102
rect 201678 346046 381250 346102
rect 381306 346046 381374 346102
rect 381430 346046 381498 346102
rect 381554 346046 381622 346102
rect 381678 346046 399250 346102
rect 399306 346046 399374 346102
rect 399430 346046 399498 346102
rect 399554 346046 399622 346102
rect 399678 346046 579250 346102
rect 579306 346046 579374 346102
rect 579430 346046 579498 346102
rect 579554 346046 579622 346102
rect 579678 346046 596496 346102
rect 596552 346046 596620 346102
rect 596676 346046 596744 346102
rect 596800 346046 596868 346102
rect 596924 346046 597980 346102
rect -1916 345978 597980 346046
rect -1916 345922 -860 345978
rect -804 345922 -736 345978
rect -680 345922 -612 345978
rect -556 345922 -488 345978
rect -432 345922 3250 345978
rect 3306 345922 3374 345978
rect 3430 345922 3498 345978
rect 3554 345922 3622 345978
rect 3678 345922 201250 345978
rect 201306 345922 201374 345978
rect 201430 345922 201498 345978
rect 201554 345922 201622 345978
rect 201678 345922 381250 345978
rect 381306 345922 381374 345978
rect 381430 345922 381498 345978
rect 381554 345922 381622 345978
rect 381678 345922 399250 345978
rect 399306 345922 399374 345978
rect 399430 345922 399498 345978
rect 399554 345922 399622 345978
rect 399678 345922 579250 345978
rect 579306 345922 579374 345978
rect 579430 345922 579498 345978
rect 579554 345922 579622 345978
rect 579678 345922 596496 345978
rect 596552 345922 596620 345978
rect 596676 345922 596744 345978
rect 596800 345922 596868 345978
rect 596924 345922 597980 345978
rect -1916 345826 597980 345922
rect -1916 334350 597980 334446
rect -1916 334294 -1820 334350
rect -1764 334294 -1696 334350
rect -1640 334294 -1572 334350
rect -1516 334294 -1448 334350
rect -1392 334294 6970 334350
rect 7026 334294 7094 334350
rect 7150 334294 7218 334350
rect 7274 334294 7342 334350
rect 7398 334294 204970 334350
rect 205026 334294 205094 334350
rect 205150 334294 205218 334350
rect 205274 334294 205342 334350
rect 205398 334294 384970 334350
rect 385026 334294 385094 334350
rect 385150 334294 385218 334350
rect 385274 334294 385342 334350
rect 385398 334294 402970 334350
rect 403026 334294 403094 334350
rect 403150 334294 403218 334350
rect 403274 334294 403342 334350
rect 403398 334294 582970 334350
rect 583026 334294 583094 334350
rect 583150 334294 583218 334350
rect 583274 334294 583342 334350
rect 583398 334294 597456 334350
rect 597512 334294 597580 334350
rect 597636 334294 597704 334350
rect 597760 334294 597828 334350
rect 597884 334294 597980 334350
rect -1916 334226 597980 334294
rect -1916 334170 -1820 334226
rect -1764 334170 -1696 334226
rect -1640 334170 -1572 334226
rect -1516 334170 -1448 334226
rect -1392 334170 6970 334226
rect 7026 334170 7094 334226
rect 7150 334170 7218 334226
rect 7274 334170 7342 334226
rect 7398 334170 204970 334226
rect 205026 334170 205094 334226
rect 205150 334170 205218 334226
rect 205274 334170 205342 334226
rect 205398 334170 384970 334226
rect 385026 334170 385094 334226
rect 385150 334170 385218 334226
rect 385274 334170 385342 334226
rect 385398 334170 402970 334226
rect 403026 334170 403094 334226
rect 403150 334170 403218 334226
rect 403274 334170 403342 334226
rect 403398 334170 582970 334226
rect 583026 334170 583094 334226
rect 583150 334170 583218 334226
rect 583274 334170 583342 334226
rect 583398 334170 597456 334226
rect 597512 334170 597580 334226
rect 597636 334170 597704 334226
rect 597760 334170 597828 334226
rect 597884 334170 597980 334226
rect -1916 334102 597980 334170
rect -1916 334046 -1820 334102
rect -1764 334046 -1696 334102
rect -1640 334046 -1572 334102
rect -1516 334046 -1448 334102
rect -1392 334046 6970 334102
rect 7026 334046 7094 334102
rect 7150 334046 7218 334102
rect 7274 334046 7342 334102
rect 7398 334046 204970 334102
rect 205026 334046 205094 334102
rect 205150 334046 205218 334102
rect 205274 334046 205342 334102
rect 205398 334046 384970 334102
rect 385026 334046 385094 334102
rect 385150 334046 385218 334102
rect 385274 334046 385342 334102
rect 385398 334046 402970 334102
rect 403026 334046 403094 334102
rect 403150 334046 403218 334102
rect 403274 334046 403342 334102
rect 403398 334046 582970 334102
rect 583026 334046 583094 334102
rect 583150 334046 583218 334102
rect 583274 334046 583342 334102
rect 583398 334046 597456 334102
rect 597512 334046 597580 334102
rect 597636 334046 597704 334102
rect 597760 334046 597828 334102
rect 597884 334046 597980 334102
rect -1916 333978 597980 334046
rect -1916 333922 -1820 333978
rect -1764 333922 -1696 333978
rect -1640 333922 -1572 333978
rect -1516 333922 -1448 333978
rect -1392 333922 6970 333978
rect 7026 333922 7094 333978
rect 7150 333922 7218 333978
rect 7274 333922 7342 333978
rect 7398 333922 204970 333978
rect 205026 333922 205094 333978
rect 205150 333922 205218 333978
rect 205274 333922 205342 333978
rect 205398 333922 384970 333978
rect 385026 333922 385094 333978
rect 385150 333922 385218 333978
rect 385274 333922 385342 333978
rect 385398 333922 402970 333978
rect 403026 333922 403094 333978
rect 403150 333922 403218 333978
rect 403274 333922 403342 333978
rect 403398 333922 582970 333978
rect 583026 333922 583094 333978
rect 583150 333922 583218 333978
rect 583274 333922 583342 333978
rect 583398 333922 597456 333978
rect 597512 333922 597580 333978
rect 597636 333922 597704 333978
rect 597760 333922 597828 333978
rect 597884 333922 597980 333978
rect -1916 333826 597980 333922
rect -1916 328350 597980 328446
rect -1916 328294 -860 328350
rect -804 328294 -736 328350
rect -680 328294 -612 328350
rect -556 328294 -488 328350
rect -432 328294 3250 328350
rect 3306 328294 3374 328350
rect 3430 328294 3498 328350
rect 3554 328294 3622 328350
rect 3678 328294 201250 328350
rect 201306 328294 201374 328350
rect 201430 328294 201498 328350
rect 201554 328294 201622 328350
rect 201678 328294 381250 328350
rect 381306 328294 381374 328350
rect 381430 328294 381498 328350
rect 381554 328294 381622 328350
rect 381678 328294 399250 328350
rect 399306 328294 399374 328350
rect 399430 328294 399498 328350
rect 399554 328294 399622 328350
rect 399678 328294 579250 328350
rect 579306 328294 579374 328350
rect 579430 328294 579498 328350
rect 579554 328294 579622 328350
rect 579678 328294 596496 328350
rect 596552 328294 596620 328350
rect 596676 328294 596744 328350
rect 596800 328294 596868 328350
rect 596924 328294 597980 328350
rect -1916 328226 597980 328294
rect -1916 328170 -860 328226
rect -804 328170 -736 328226
rect -680 328170 -612 328226
rect -556 328170 -488 328226
rect -432 328170 3250 328226
rect 3306 328170 3374 328226
rect 3430 328170 3498 328226
rect 3554 328170 3622 328226
rect 3678 328170 201250 328226
rect 201306 328170 201374 328226
rect 201430 328170 201498 328226
rect 201554 328170 201622 328226
rect 201678 328170 381250 328226
rect 381306 328170 381374 328226
rect 381430 328170 381498 328226
rect 381554 328170 381622 328226
rect 381678 328170 399250 328226
rect 399306 328170 399374 328226
rect 399430 328170 399498 328226
rect 399554 328170 399622 328226
rect 399678 328170 579250 328226
rect 579306 328170 579374 328226
rect 579430 328170 579498 328226
rect 579554 328170 579622 328226
rect 579678 328170 596496 328226
rect 596552 328170 596620 328226
rect 596676 328170 596744 328226
rect 596800 328170 596868 328226
rect 596924 328170 597980 328226
rect -1916 328102 597980 328170
rect -1916 328046 -860 328102
rect -804 328046 -736 328102
rect -680 328046 -612 328102
rect -556 328046 -488 328102
rect -432 328046 3250 328102
rect 3306 328046 3374 328102
rect 3430 328046 3498 328102
rect 3554 328046 3622 328102
rect 3678 328046 201250 328102
rect 201306 328046 201374 328102
rect 201430 328046 201498 328102
rect 201554 328046 201622 328102
rect 201678 328046 381250 328102
rect 381306 328046 381374 328102
rect 381430 328046 381498 328102
rect 381554 328046 381622 328102
rect 381678 328046 399250 328102
rect 399306 328046 399374 328102
rect 399430 328046 399498 328102
rect 399554 328046 399622 328102
rect 399678 328046 579250 328102
rect 579306 328046 579374 328102
rect 579430 328046 579498 328102
rect 579554 328046 579622 328102
rect 579678 328046 596496 328102
rect 596552 328046 596620 328102
rect 596676 328046 596744 328102
rect 596800 328046 596868 328102
rect 596924 328046 597980 328102
rect -1916 327978 597980 328046
rect -1916 327922 -860 327978
rect -804 327922 -736 327978
rect -680 327922 -612 327978
rect -556 327922 -488 327978
rect -432 327922 3250 327978
rect 3306 327922 3374 327978
rect 3430 327922 3498 327978
rect 3554 327922 3622 327978
rect 3678 327922 201250 327978
rect 201306 327922 201374 327978
rect 201430 327922 201498 327978
rect 201554 327922 201622 327978
rect 201678 327922 381250 327978
rect 381306 327922 381374 327978
rect 381430 327922 381498 327978
rect 381554 327922 381622 327978
rect 381678 327922 399250 327978
rect 399306 327922 399374 327978
rect 399430 327922 399498 327978
rect 399554 327922 399622 327978
rect 399678 327922 579250 327978
rect 579306 327922 579374 327978
rect 579430 327922 579498 327978
rect 579554 327922 579622 327978
rect 579678 327922 596496 327978
rect 596552 327922 596620 327978
rect 596676 327922 596744 327978
rect 596800 327922 596868 327978
rect 596924 327922 597980 327978
rect -1916 327826 597980 327922
rect -1916 316350 597980 316446
rect -1916 316294 -1820 316350
rect -1764 316294 -1696 316350
rect -1640 316294 -1572 316350
rect -1516 316294 -1448 316350
rect -1392 316294 6970 316350
rect 7026 316294 7094 316350
rect 7150 316294 7218 316350
rect 7274 316294 7342 316350
rect 7398 316294 24970 316350
rect 25026 316294 25094 316350
rect 25150 316294 25218 316350
rect 25274 316294 25342 316350
rect 25398 316294 42970 316350
rect 43026 316294 43094 316350
rect 43150 316294 43218 316350
rect 43274 316294 43342 316350
rect 43398 316294 60970 316350
rect 61026 316294 61094 316350
rect 61150 316294 61218 316350
rect 61274 316294 61342 316350
rect 61398 316294 78970 316350
rect 79026 316294 79094 316350
rect 79150 316294 79218 316350
rect 79274 316294 79342 316350
rect 79398 316294 96970 316350
rect 97026 316294 97094 316350
rect 97150 316294 97218 316350
rect 97274 316294 97342 316350
rect 97398 316294 114970 316350
rect 115026 316294 115094 316350
rect 115150 316294 115218 316350
rect 115274 316294 115342 316350
rect 115398 316294 132970 316350
rect 133026 316294 133094 316350
rect 133150 316294 133218 316350
rect 133274 316294 133342 316350
rect 133398 316294 150970 316350
rect 151026 316294 151094 316350
rect 151150 316294 151218 316350
rect 151274 316294 151342 316350
rect 151398 316294 168970 316350
rect 169026 316294 169094 316350
rect 169150 316294 169218 316350
rect 169274 316294 169342 316350
rect 169398 316294 186970 316350
rect 187026 316294 187094 316350
rect 187150 316294 187218 316350
rect 187274 316294 187342 316350
rect 187398 316294 204970 316350
rect 205026 316294 205094 316350
rect 205150 316294 205218 316350
rect 205274 316294 205342 316350
rect 205398 316294 222970 316350
rect 223026 316294 223094 316350
rect 223150 316294 223218 316350
rect 223274 316294 223342 316350
rect 223398 316294 240970 316350
rect 241026 316294 241094 316350
rect 241150 316294 241218 316350
rect 241274 316294 241342 316350
rect 241398 316294 258970 316350
rect 259026 316294 259094 316350
rect 259150 316294 259218 316350
rect 259274 316294 259342 316350
rect 259398 316294 276970 316350
rect 277026 316294 277094 316350
rect 277150 316294 277218 316350
rect 277274 316294 277342 316350
rect 277398 316294 294970 316350
rect 295026 316294 295094 316350
rect 295150 316294 295218 316350
rect 295274 316294 295342 316350
rect 295398 316294 312970 316350
rect 313026 316294 313094 316350
rect 313150 316294 313218 316350
rect 313274 316294 313342 316350
rect 313398 316294 330970 316350
rect 331026 316294 331094 316350
rect 331150 316294 331218 316350
rect 331274 316294 331342 316350
rect 331398 316294 348970 316350
rect 349026 316294 349094 316350
rect 349150 316294 349218 316350
rect 349274 316294 349342 316350
rect 349398 316294 366970 316350
rect 367026 316294 367094 316350
rect 367150 316294 367218 316350
rect 367274 316294 367342 316350
rect 367398 316294 384970 316350
rect 385026 316294 385094 316350
rect 385150 316294 385218 316350
rect 385274 316294 385342 316350
rect 385398 316294 402970 316350
rect 403026 316294 403094 316350
rect 403150 316294 403218 316350
rect 403274 316294 403342 316350
rect 403398 316294 420970 316350
rect 421026 316294 421094 316350
rect 421150 316294 421218 316350
rect 421274 316294 421342 316350
rect 421398 316294 438970 316350
rect 439026 316294 439094 316350
rect 439150 316294 439218 316350
rect 439274 316294 439342 316350
rect 439398 316294 456970 316350
rect 457026 316294 457094 316350
rect 457150 316294 457218 316350
rect 457274 316294 457342 316350
rect 457398 316294 474970 316350
rect 475026 316294 475094 316350
rect 475150 316294 475218 316350
rect 475274 316294 475342 316350
rect 475398 316294 492970 316350
rect 493026 316294 493094 316350
rect 493150 316294 493218 316350
rect 493274 316294 493342 316350
rect 493398 316294 510970 316350
rect 511026 316294 511094 316350
rect 511150 316294 511218 316350
rect 511274 316294 511342 316350
rect 511398 316294 528970 316350
rect 529026 316294 529094 316350
rect 529150 316294 529218 316350
rect 529274 316294 529342 316350
rect 529398 316294 546970 316350
rect 547026 316294 547094 316350
rect 547150 316294 547218 316350
rect 547274 316294 547342 316350
rect 547398 316294 564970 316350
rect 565026 316294 565094 316350
rect 565150 316294 565218 316350
rect 565274 316294 565342 316350
rect 565398 316294 582970 316350
rect 583026 316294 583094 316350
rect 583150 316294 583218 316350
rect 583274 316294 583342 316350
rect 583398 316294 597456 316350
rect 597512 316294 597580 316350
rect 597636 316294 597704 316350
rect 597760 316294 597828 316350
rect 597884 316294 597980 316350
rect -1916 316226 597980 316294
rect -1916 316170 -1820 316226
rect -1764 316170 -1696 316226
rect -1640 316170 -1572 316226
rect -1516 316170 -1448 316226
rect -1392 316170 6970 316226
rect 7026 316170 7094 316226
rect 7150 316170 7218 316226
rect 7274 316170 7342 316226
rect 7398 316170 24970 316226
rect 25026 316170 25094 316226
rect 25150 316170 25218 316226
rect 25274 316170 25342 316226
rect 25398 316170 42970 316226
rect 43026 316170 43094 316226
rect 43150 316170 43218 316226
rect 43274 316170 43342 316226
rect 43398 316170 60970 316226
rect 61026 316170 61094 316226
rect 61150 316170 61218 316226
rect 61274 316170 61342 316226
rect 61398 316170 78970 316226
rect 79026 316170 79094 316226
rect 79150 316170 79218 316226
rect 79274 316170 79342 316226
rect 79398 316170 96970 316226
rect 97026 316170 97094 316226
rect 97150 316170 97218 316226
rect 97274 316170 97342 316226
rect 97398 316170 114970 316226
rect 115026 316170 115094 316226
rect 115150 316170 115218 316226
rect 115274 316170 115342 316226
rect 115398 316170 132970 316226
rect 133026 316170 133094 316226
rect 133150 316170 133218 316226
rect 133274 316170 133342 316226
rect 133398 316170 150970 316226
rect 151026 316170 151094 316226
rect 151150 316170 151218 316226
rect 151274 316170 151342 316226
rect 151398 316170 168970 316226
rect 169026 316170 169094 316226
rect 169150 316170 169218 316226
rect 169274 316170 169342 316226
rect 169398 316170 186970 316226
rect 187026 316170 187094 316226
rect 187150 316170 187218 316226
rect 187274 316170 187342 316226
rect 187398 316170 204970 316226
rect 205026 316170 205094 316226
rect 205150 316170 205218 316226
rect 205274 316170 205342 316226
rect 205398 316170 222970 316226
rect 223026 316170 223094 316226
rect 223150 316170 223218 316226
rect 223274 316170 223342 316226
rect 223398 316170 240970 316226
rect 241026 316170 241094 316226
rect 241150 316170 241218 316226
rect 241274 316170 241342 316226
rect 241398 316170 258970 316226
rect 259026 316170 259094 316226
rect 259150 316170 259218 316226
rect 259274 316170 259342 316226
rect 259398 316170 276970 316226
rect 277026 316170 277094 316226
rect 277150 316170 277218 316226
rect 277274 316170 277342 316226
rect 277398 316170 294970 316226
rect 295026 316170 295094 316226
rect 295150 316170 295218 316226
rect 295274 316170 295342 316226
rect 295398 316170 312970 316226
rect 313026 316170 313094 316226
rect 313150 316170 313218 316226
rect 313274 316170 313342 316226
rect 313398 316170 330970 316226
rect 331026 316170 331094 316226
rect 331150 316170 331218 316226
rect 331274 316170 331342 316226
rect 331398 316170 348970 316226
rect 349026 316170 349094 316226
rect 349150 316170 349218 316226
rect 349274 316170 349342 316226
rect 349398 316170 366970 316226
rect 367026 316170 367094 316226
rect 367150 316170 367218 316226
rect 367274 316170 367342 316226
rect 367398 316170 384970 316226
rect 385026 316170 385094 316226
rect 385150 316170 385218 316226
rect 385274 316170 385342 316226
rect 385398 316170 402970 316226
rect 403026 316170 403094 316226
rect 403150 316170 403218 316226
rect 403274 316170 403342 316226
rect 403398 316170 420970 316226
rect 421026 316170 421094 316226
rect 421150 316170 421218 316226
rect 421274 316170 421342 316226
rect 421398 316170 438970 316226
rect 439026 316170 439094 316226
rect 439150 316170 439218 316226
rect 439274 316170 439342 316226
rect 439398 316170 456970 316226
rect 457026 316170 457094 316226
rect 457150 316170 457218 316226
rect 457274 316170 457342 316226
rect 457398 316170 474970 316226
rect 475026 316170 475094 316226
rect 475150 316170 475218 316226
rect 475274 316170 475342 316226
rect 475398 316170 492970 316226
rect 493026 316170 493094 316226
rect 493150 316170 493218 316226
rect 493274 316170 493342 316226
rect 493398 316170 510970 316226
rect 511026 316170 511094 316226
rect 511150 316170 511218 316226
rect 511274 316170 511342 316226
rect 511398 316170 528970 316226
rect 529026 316170 529094 316226
rect 529150 316170 529218 316226
rect 529274 316170 529342 316226
rect 529398 316170 546970 316226
rect 547026 316170 547094 316226
rect 547150 316170 547218 316226
rect 547274 316170 547342 316226
rect 547398 316170 564970 316226
rect 565026 316170 565094 316226
rect 565150 316170 565218 316226
rect 565274 316170 565342 316226
rect 565398 316170 582970 316226
rect 583026 316170 583094 316226
rect 583150 316170 583218 316226
rect 583274 316170 583342 316226
rect 583398 316170 597456 316226
rect 597512 316170 597580 316226
rect 597636 316170 597704 316226
rect 597760 316170 597828 316226
rect 597884 316170 597980 316226
rect -1916 316102 597980 316170
rect -1916 316046 -1820 316102
rect -1764 316046 -1696 316102
rect -1640 316046 -1572 316102
rect -1516 316046 -1448 316102
rect -1392 316046 6970 316102
rect 7026 316046 7094 316102
rect 7150 316046 7218 316102
rect 7274 316046 7342 316102
rect 7398 316046 24970 316102
rect 25026 316046 25094 316102
rect 25150 316046 25218 316102
rect 25274 316046 25342 316102
rect 25398 316046 42970 316102
rect 43026 316046 43094 316102
rect 43150 316046 43218 316102
rect 43274 316046 43342 316102
rect 43398 316046 60970 316102
rect 61026 316046 61094 316102
rect 61150 316046 61218 316102
rect 61274 316046 61342 316102
rect 61398 316046 78970 316102
rect 79026 316046 79094 316102
rect 79150 316046 79218 316102
rect 79274 316046 79342 316102
rect 79398 316046 96970 316102
rect 97026 316046 97094 316102
rect 97150 316046 97218 316102
rect 97274 316046 97342 316102
rect 97398 316046 114970 316102
rect 115026 316046 115094 316102
rect 115150 316046 115218 316102
rect 115274 316046 115342 316102
rect 115398 316046 132970 316102
rect 133026 316046 133094 316102
rect 133150 316046 133218 316102
rect 133274 316046 133342 316102
rect 133398 316046 150970 316102
rect 151026 316046 151094 316102
rect 151150 316046 151218 316102
rect 151274 316046 151342 316102
rect 151398 316046 168970 316102
rect 169026 316046 169094 316102
rect 169150 316046 169218 316102
rect 169274 316046 169342 316102
rect 169398 316046 186970 316102
rect 187026 316046 187094 316102
rect 187150 316046 187218 316102
rect 187274 316046 187342 316102
rect 187398 316046 204970 316102
rect 205026 316046 205094 316102
rect 205150 316046 205218 316102
rect 205274 316046 205342 316102
rect 205398 316046 222970 316102
rect 223026 316046 223094 316102
rect 223150 316046 223218 316102
rect 223274 316046 223342 316102
rect 223398 316046 240970 316102
rect 241026 316046 241094 316102
rect 241150 316046 241218 316102
rect 241274 316046 241342 316102
rect 241398 316046 258970 316102
rect 259026 316046 259094 316102
rect 259150 316046 259218 316102
rect 259274 316046 259342 316102
rect 259398 316046 276970 316102
rect 277026 316046 277094 316102
rect 277150 316046 277218 316102
rect 277274 316046 277342 316102
rect 277398 316046 294970 316102
rect 295026 316046 295094 316102
rect 295150 316046 295218 316102
rect 295274 316046 295342 316102
rect 295398 316046 312970 316102
rect 313026 316046 313094 316102
rect 313150 316046 313218 316102
rect 313274 316046 313342 316102
rect 313398 316046 330970 316102
rect 331026 316046 331094 316102
rect 331150 316046 331218 316102
rect 331274 316046 331342 316102
rect 331398 316046 348970 316102
rect 349026 316046 349094 316102
rect 349150 316046 349218 316102
rect 349274 316046 349342 316102
rect 349398 316046 366970 316102
rect 367026 316046 367094 316102
rect 367150 316046 367218 316102
rect 367274 316046 367342 316102
rect 367398 316046 384970 316102
rect 385026 316046 385094 316102
rect 385150 316046 385218 316102
rect 385274 316046 385342 316102
rect 385398 316046 402970 316102
rect 403026 316046 403094 316102
rect 403150 316046 403218 316102
rect 403274 316046 403342 316102
rect 403398 316046 420970 316102
rect 421026 316046 421094 316102
rect 421150 316046 421218 316102
rect 421274 316046 421342 316102
rect 421398 316046 438970 316102
rect 439026 316046 439094 316102
rect 439150 316046 439218 316102
rect 439274 316046 439342 316102
rect 439398 316046 456970 316102
rect 457026 316046 457094 316102
rect 457150 316046 457218 316102
rect 457274 316046 457342 316102
rect 457398 316046 474970 316102
rect 475026 316046 475094 316102
rect 475150 316046 475218 316102
rect 475274 316046 475342 316102
rect 475398 316046 492970 316102
rect 493026 316046 493094 316102
rect 493150 316046 493218 316102
rect 493274 316046 493342 316102
rect 493398 316046 510970 316102
rect 511026 316046 511094 316102
rect 511150 316046 511218 316102
rect 511274 316046 511342 316102
rect 511398 316046 528970 316102
rect 529026 316046 529094 316102
rect 529150 316046 529218 316102
rect 529274 316046 529342 316102
rect 529398 316046 546970 316102
rect 547026 316046 547094 316102
rect 547150 316046 547218 316102
rect 547274 316046 547342 316102
rect 547398 316046 564970 316102
rect 565026 316046 565094 316102
rect 565150 316046 565218 316102
rect 565274 316046 565342 316102
rect 565398 316046 582970 316102
rect 583026 316046 583094 316102
rect 583150 316046 583218 316102
rect 583274 316046 583342 316102
rect 583398 316046 597456 316102
rect 597512 316046 597580 316102
rect 597636 316046 597704 316102
rect 597760 316046 597828 316102
rect 597884 316046 597980 316102
rect -1916 315978 597980 316046
rect -1916 315922 -1820 315978
rect -1764 315922 -1696 315978
rect -1640 315922 -1572 315978
rect -1516 315922 -1448 315978
rect -1392 315922 6970 315978
rect 7026 315922 7094 315978
rect 7150 315922 7218 315978
rect 7274 315922 7342 315978
rect 7398 315922 24970 315978
rect 25026 315922 25094 315978
rect 25150 315922 25218 315978
rect 25274 315922 25342 315978
rect 25398 315922 42970 315978
rect 43026 315922 43094 315978
rect 43150 315922 43218 315978
rect 43274 315922 43342 315978
rect 43398 315922 60970 315978
rect 61026 315922 61094 315978
rect 61150 315922 61218 315978
rect 61274 315922 61342 315978
rect 61398 315922 78970 315978
rect 79026 315922 79094 315978
rect 79150 315922 79218 315978
rect 79274 315922 79342 315978
rect 79398 315922 96970 315978
rect 97026 315922 97094 315978
rect 97150 315922 97218 315978
rect 97274 315922 97342 315978
rect 97398 315922 114970 315978
rect 115026 315922 115094 315978
rect 115150 315922 115218 315978
rect 115274 315922 115342 315978
rect 115398 315922 132970 315978
rect 133026 315922 133094 315978
rect 133150 315922 133218 315978
rect 133274 315922 133342 315978
rect 133398 315922 150970 315978
rect 151026 315922 151094 315978
rect 151150 315922 151218 315978
rect 151274 315922 151342 315978
rect 151398 315922 168970 315978
rect 169026 315922 169094 315978
rect 169150 315922 169218 315978
rect 169274 315922 169342 315978
rect 169398 315922 186970 315978
rect 187026 315922 187094 315978
rect 187150 315922 187218 315978
rect 187274 315922 187342 315978
rect 187398 315922 204970 315978
rect 205026 315922 205094 315978
rect 205150 315922 205218 315978
rect 205274 315922 205342 315978
rect 205398 315922 222970 315978
rect 223026 315922 223094 315978
rect 223150 315922 223218 315978
rect 223274 315922 223342 315978
rect 223398 315922 240970 315978
rect 241026 315922 241094 315978
rect 241150 315922 241218 315978
rect 241274 315922 241342 315978
rect 241398 315922 258970 315978
rect 259026 315922 259094 315978
rect 259150 315922 259218 315978
rect 259274 315922 259342 315978
rect 259398 315922 276970 315978
rect 277026 315922 277094 315978
rect 277150 315922 277218 315978
rect 277274 315922 277342 315978
rect 277398 315922 294970 315978
rect 295026 315922 295094 315978
rect 295150 315922 295218 315978
rect 295274 315922 295342 315978
rect 295398 315922 312970 315978
rect 313026 315922 313094 315978
rect 313150 315922 313218 315978
rect 313274 315922 313342 315978
rect 313398 315922 330970 315978
rect 331026 315922 331094 315978
rect 331150 315922 331218 315978
rect 331274 315922 331342 315978
rect 331398 315922 348970 315978
rect 349026 315922 349094 315978
rect 349150 315922 349218 315978
rect 349274 315922 349342 315978
rect 349398 315922 366970 315978
rect 367026 315922 367094 315978
rect 367150 315922 367218 315978
rect 367274 315922 367342 315978
rect 367398 315922 384970 315978
rect 385026 315922 385094 315978
rect 385150 315922 385218 315978
rect 385274 315922 385342 315978
rect 385398 315922 402970 315978
rect 403026 315922 403094 315978
rect 403150 315922 403218 315978
rect 403274 315922 403342 315978
rect 403398 315922 420970 315978
rect 421026 315922 421094 315978
rect 421150 315922 421218 315978
rect 421274 315922 421342 315978
rect 421398 315922 438970 315978
rect 439026 315922 439094 315978
rect 439150 315922 439218 315978
rect 439274 315922 439342 315978
rect 439398 315922 456970 315978
rect 457026 315922 457094 315978
rect 457150 315922 457218 315978
rect 457274 315922 457342 315978
rect 457398 315922 474970 315978
rect 475026 315922 475094 315978
rect 475150 315922 475218 315978
rect 475274 315922 475342 315978
rect 475398 315922 492970 315978
rect 493026 315922 493094 315978
rect 493150 315922 493218 315978
rect 493274 315922 493342 315978
rect 493398 315922 510970 315978
rect 511026 315922 511094 315978
rect 511150 315922 511218 315978
rect 511274 315922 511342 315978
rect 511398 315922 528970 315978
rect 529026 315922 529094 315978
rect 529150 315922 529218 315978
rect 529274 315922 529342 315978
rect 529398 315922 546970 315978
rect 547026 315922 547094 315978
rect 547150 315922 547218 315978
rect 547274 315922 547342 315978
rect 547398 315922 564970 315978
rect 565026 315922 565094 315978
rect 565150 315922 565218 315978
rect 565274 315922 565342 315978
rect 565398 315922 582970 315978
rect 583026 315922 583094 315978
rect 583150 315922 583218 315978
rect 583274 315922 583342 315978
rect 583398 315922 597456 315978
rect 597512 315922 597580 315978
rect 597636 315922 597704 315978
rect 597760 315922 597828 315978
rect 597884 315922 597980 315978
rect -1916 315826 597980 315922
rect -1916 310350 597980 310446
rect -1916 310294 -860 310350
rect -804 310294 -736 310350
rect -680 310294 -612 310350
rect -556 310294 -488 310350
rect -432 310294 3250 310350
rect 3306 310294 3374 310350
rect 3430 310294 3498 310350
rect 3554 310294 3622 310350
rect 3678 310294 201250 310350
rect 201306 310294 201374 310350
rect 201430 310294 201498 310350
rect 201554 310294 201622 310350
rect 201678 310294 381250 310350
rect 381306 310294 381374 310350
rect 381430 310294 381498 310350
rect 381554 310294 381622 310350
rect 381678 310294 399250 310350
rect 399306 310294 399374 310350
rect 399430 310294 399498 310350
rect 399554 310294 399622 310350
rect 399678 310294 579250 310350
rect 579306 310294 579374 310350
rect 579430 310294 579498 310350
rect 579554 310294 579622 310350
rect 579678 310294 596496 310350
rect 596552 310294 596620 310350
rect 596676 310294 596744 310350
rect 596800 310294 596868 310350
rect 596924 310294 597980 310350
rect -1916 310226 597980 310294
rect -1916 310170 -860 310226
rect -804 310170 -736 310226
rect -680 310170 -612 310226
rect -556 310170 -488 310226
rect -432 310170 3250 310226
rect 3306 310170 3374 310226
rect 3430 310170 3498 310226
rect 3554 310170 3622 310226
rect 3678 310170 201250 310226
rect 201306 310170 201374 310226
rect 201430 310170 201498 310226
rect 201554 310170 201622 310226
rect 201678 310170 381250 310226
rect 381306 310170 381374 310226
rect 381430 310170 381498 310226
rect 381554 310170 381622 310226
rect 381678 310170 399250 310226
rect 399306 310170 399374 310226
rect 399430 310170 399498 310226
rect 399554 310170 399622 310226
rect 399678 310170 579250 310226
rect 579306 310170 579374 310226
rect 579430 310170 579498 310226
rect 579554 310170 579622 310226
rect 579678 310170 596496 310226
rect 596552 310170 596620 310226
rect 596676 310170 596744 310226
rect 596800 310170 596868 310226
rect 596924 310170 597980 310226
rect -1916 310102 597980 310170
rect -1916 310046 -860 310102
rect -804 310046 -736 310102
rect -680 310046 -612 310102
rect -556 310046 -488 310102
rect -432 310046 3250 310102
rect 3306 310046 3374 310102
rect 3430 310046 3498 310102
rect 3554 310046 3622 310102
rect 3678 310046 201250 310102
rect 201306 310046 201374 310102
rect 201430 310046 201498 310102
rect 201554 310046 201622 310102
rect 201678 310046 381250 310102
rect 381306 310046 381374 310102
rect 381430 310046 381498 310102
rect 381554 310046 381622 310102
rect 381678 310046 399250 310102
rect 399306 310046 399374 310102
rect 399430 310046 399498 310102
rect 399554 310046 399622 310102
rect 399678 310046 579250 310102
rect 579306 310046 579374 310102
rect 579430 310046 579498 310102
rect 579554 310046 579622 310102
rect 579678 310046 596496 310102
rect 596552 310046 596620 310102
rect 596676 310046 596744 310102
rect 596800 310046 596868 310102
rect 596924 310046 597980 310102
rect -1916 309978 597980 310046
rect -1916 309922 -860 309978
rect -804 309922 -736 309978
rect -680 309922 -612 309978
rect -556 309922 -488 309978
rect -432 309922 3250 309978
rect 3306 309922 3374 309978
rect 3430 309922 3498 309978
rect 3554 309922 3622 309978
rect 3678 309922 201250 309978
rect 201306 309922 201374 309978
rect 201430 309922 201498 309978
rect 201554 309922 201622 309978
rect 201678 309922 381250 309978
rect 381306 309922 381374 309978
rect 381430 309922 381498 309978
rect 381554 309922 381622 309978
rect 381678 309922 399250 309978
rect 399306 309922 399374 309978
rect 399430 309922 399498 309978
rect 399554 309922 399622 309978
rect 399678 309922 579250 309978
rect 579306 309922 579374 309978
rect 579430 309922 579498 309978
rect 579554 309922 579622 309978
rect 579678 309922 596496 309978
rect 596552 309922 596620 309978
rect 596676 309922 596744 309978
rect 596800 309922 596868 309978
rect 596924 309922 597980 309978
rect -1916 309826 597980 309922
rect -1916 298422 597980 298446
rect -1916 298366 24970 298422
rect 25026 298366 25094 298422
rect 25150 298366 25218 298422
rect 25274 298366 25342 298422
rect 25398 298366 42970 298422
rect 43026 298366 43094 298422
rect 43150 298366 43218 298422
rect 43274 298366 43342 298422
rect 43398 298366 60970 298422
rect 61026 298366 61094 298422
rect 61150 298366 61218 298422
rect 61274 298366 61342 298422
rect 61398 298366 78970 298422
rect 79026 298366 79094 298422
rect 79150 298366 79218 298422
rect 79274 298366 79342 298422
rect 79398 298366 96970 298422
rect 97026 298366 97094 298422
rect 97150 298366 97218 298422
rect 97274 298366 97342 298422
rect 97398 298366 114970 298422
rect 115026 298366 115094 298422
rect 115150 298366 115218 298422
rect 115274 298366 115342 298422
rect 115398 298366 132970 298422
rect 133026 298366 133094 298422
rect 133150 298366 133218 298422
rect 133274 298366 133342 298422
rect 133398 298366 150970 298422
rect 151026 298366 151094 298422
rect 151150 298366 151218 298422
rect 151274 298366 151342 298422
rect 151398 298366 168970 298422
rect 169026 298366 169094 298422
rect 169150 298366 169218 298422
rect 169274 298366 169342 298422
rect 169398 298366 186970 298422
rect 187026 298366 187094 298422
rect 187150 298366 187218 298422
rect 187274 298366 187342 298422
rect 187398 298366 222970 298422
rect 223026 298366 223094 298422
rect 223150 298366 223218 298422
rect 223274 298366 223342 298422
rect 223398 298366 240970 298422
rect 241026 298366 241094 298422
rect 241150 298366 241218 298422
rect 241274 298366 241342 298422
rect 241398 298366 258970 298422
rect 259026 298366 259094 298422
rect 259150 298366 259218 298422
rect 259274 298366 259342 298422
rect 259398 298366 276970 298422
rect 277026 298366 277094 298422
rect 277150 298366 277218 298422
rect 277274 298366 277342 298422
rect 277398 298366 294970 298422
rect 295026 298366 295094 298422
rect 295150 298366 295218 298422
rect 295274 298366 295342 298422
rect 295398 298366 312970 298422
rect 313026 298366 313094 298422
rect 313150 298366 313218 298422
rect 313274 298366 313342 298422
rect 313398 298366 330970 298422
rect 331026 298366 331094 298422
rect 331150 298366 331218 298422
rect 331274 298366 331342 298422
rect 331398 298366 348970 298422
rect 349026 298366 349094 298422
rect 349150 298366 349218 298422
rect 349274 298366 349342 298422
rect 349398 298366 366970 298422
rect 367026 298366 367094 298422
rect 367150 298366 367218 298422
rect 367274 298366 367342 298422
rect 367398 298366 420970 298422
rect 421026 298366 421094 298422
rect 421150 298366 421218 298422
rect 421274 298366 421342 298422
rect 421398 298366 438970 298422
rect 439026 298366 439094 298422
rect 439150 298366 439218 298422
rect 439274 298366 439342 298422
rect 439398 298366 456970 298422
rect 457026 298366 457094 298422
rect 457150 298366 457218 298422
rect 457274 298366 457342 298422
rect 457398 298366 474970 298422
rect 475026 298366 475094 298422
rect 475150 298366 475218 298422
rect 475274 298366 475342 298422
rect 475398 298366 492970 298422
rect 493026 298366 493094 298422
rect 493150 298366 493218 298422
rect 493274 298366 493342 298422
rect 493398 298366 510970 298422
rect 511026 298366 511094 298422
rect 511150 298366 511218 298422
rect 511274 298366 511342 298422
rect 511398 298366 528970 298422
rect 529026 298366 529094 298422
rect 529150 298366 529218 298422
rect 529274 298366 529342 298422
rect 529398 298366 546970 298422
rect 547026 298366 547094 298422
rect 547150 298366 547218 298422
rect 547274 298366 547342 298422
rect 547398 298366 564970 298422
rect 565026 298366 565094 298422
rect 565150 298366 565218 298422
rect 565274 298366 565342 298422
rect 565398 298366 597980 298422
rect -1916 298350 597980 298366
rect -1916 298294 -1820 298350
rect -1764 298294 -1696 298350
rect -1640 298294 -1572 298350
rect -1516 298294 -1448 298350
rect -1392 298294 6970 298350
rect 7026 298294 7094 298350
rect 7150 298294 7218 298350
rect 7274 298294 7342 298350
rect 7398 298294 204970 298350
rect 205026 298294 205094 298350
rect 205150 298294 205218 298350
rect 205274 298294 205342 298350
rect 205398 298294 384970 298350
rect 385026 298294 385094 298350
rect 385150 298294 385218 298350
rect 385274 298294 385342 298350
rect 385398 298294 402970 298350
rect 403026 298294 403094 298350
rect 403150 298294 403218 298350
rect 403274 298294 403342 298350
rect 403398 298294 582970 298350
rect 583026 298294 583094 298350
rect 583150 298294 583218 298350
rect 583274 298294 583342 298350
rect 583398 298294 597456 298350
rect 597512 298294 597580 298350
rect 597636 298294 597704 298350
rect 597760 298294 597828 298350
rect 597884 298294 597980 298350
rect -1916 298226 597980 298294
rect -1916 298170 -1820 298226
rect -1764 298170 -1696 298226
rect -1640 298170 -1572 298226
rect -1516 298170 -1448 298226
rect -1392 298170 6970 298226
rect 7026 298170 7094 298226
rect 7150 298170 7218 298226
rect 7274 298170 7342 298226
rect 7398 298170 204970 298226
rect 205026 298170 205094 298226
rect 205150 298170 205218 298226
rect 205274 298170 205342 298226
rect 205398 298170 384970 298226
rect 385026 298170 385094 298226
rect 385150 298170 385218 298226
rect 385274 298170 385342 298226
rect 385398 298170 402970 298226
rect 403026 298170 403094 298226
rect 403150 298170 403218 298226
rect 403274 298170 403342 298226
rect 403398 298170 582970 298226
rect 583026 298170 583094 298226
rect 583150 298170 583218 298226
rect 583274 298170 583342 298226
rect 583398 298170 597456 298226
rect 597512 298170 597580 298226
rect 597636 298170 597704 298226
rect 597760 298170 597828 298226
rect 597884 298170 597980 298226
rect -1916 298102 597980 298170
rect -1916 298046 -1820 298102
rect -1764 298046 -1696 298102
rect -1640 298046 -1572 298102
rect -1516 298046 -1448 298102
rect -1392 298046 6970 298102
rect 7026 298046 7094 298102
rect 7150 298046 7218 298102
rect 7274 298046 7342 298102
rect 7398 298046 204970 298102
rect 205026 298046 205094 298102
rect 205150 298046 205218 298102
rect 205274 298046 205342 298102
rect 205398 298046 384970 298102
rect 385026 298046 385094 298102
rect 385150 298046 385218 298102
rect 385274 298046 385342 298102
rect 385398 298046 402970 298102
rect 403026 298046 403094 298102
rect 403150 298046 403218 298102
rect 403274 298046 403342 298102
rect 403398 298046 582970 298102
rect 583026 298046 583094 298102
rect 583150 298046 583218 298102
rect 583274 298046 583342 298102
rect 583398 298046 597456 298102
rect 597512 298046 597580 298102
rect 597636 298046 597704 298102
rect 597760 298046 597828 298102
rect 597884 298046 597980 298102
rect -1916 297978 597980 298046
rect -1916 297922 -1820 297978
rect -1764 297922 -1696 297978
rect -1640 297922 -1572 297978
rect -1516 297922 -1448 297978
rect -1392 297922 6970 297978
rect 7026 297922 7094 297978
rect 7150 297922 7218 297978
rect 7274 297922 7342 297978
rect 7398 297922 204970 297978
rect 205026 297922 205094 297978
rect 205150 297922 205218 297978
rect 205274 297922 205342 297978
rect 205398 297922 384970 297978
rect 385026 297922 385094 297978
rect 385150 297922 385218 297978
rect 385274 297922 385342 297978
rect 385398 297922 402970 297978
rect 403026 297922 403094 297978
rect 403150 297922 403218 297978
rect 403274 297922 403342 297978
rect 403398 297922 582970 297978
rect 583026 297922 583094 297978
rect 583150 297922 583218 297978
rect 583274 297922 583342 297978
rect 583398 297922 597456 297978
rect 597512 297922 597580 297978
rect 597636 297922 597704 297978
rect 597760 297922 597828 297978
rect 597884 297922 597980 297978
rect -1916 297826 597980 297922
rect -1916 292350 597980 292446
rect -1916 292294 -860 292350
rect -804 292294 -736 292350
rect -680 292294 -612 292350
rect -556 292294 -488 292350
rect -432 292294 3250 292350
rect 3306 292294 3374 292350
rect 3430 292294 3498 292350
rect 3554 292294 3622 292350
rect 3678 292294 201250 292350
rect 201306 292294 201374 292350
rect 201430 292294 201498 292350
rect 201554 292294 201622 292350
rect 201678 292294 381250 292350
rect 381306 292294 381374 292350
rect 381430 292294 381498 292350
rect 381554 292294 381622 292350
rect 381678 292294 399250 292350
rect 399306 292294 399374 292350
rect 399430 292294 399498 292350
rect 399554 292294 399622 292350
rect 399678 292294 579250 292350
rect 579306 292294 579374 292350
rect 579430 292294 579498 292350
rect 579554 292294 579622 292350
rect 579678 292294 596496 292350
rect 596552 292294 596620 292350
rect 596676 292294 596744 292350
rect 596800 292294 596868 292350
rect 596924 292294 597980 292350
rect -1916 292226 597980 292294
rect -1916 292170 -860 292226
rect -804 292170 -736 292226
rect -680 292170 -612 292226
rect -556 292170 -488 292226
rect -432 292170 3250 292226
rect 3306 292170 3374 292226
rect 3430 292170 3498 292226
rect 3554 292170 3622 292226
rect 3678 292170 201250 292226
rect 201306 292170 201374 292226
rect 201430 292170 201498 292226
rect 201554 292170 201622 292226
rect 201678 292170 381250 292226
rect 381306 292170 381374 292226
rect 381430 292170 381498 292226
rect 381554 292170 381622 292226
rect 381678 292170 399250 292226
rect 399306 292170 399374 292226
rect 399430 292170 399498 292226
rect 399554 292170 399622 292226
rect 399678 292170 579250 292226
rect 579306 292170 579374 292226
rect 579430 292170 579498 292226
rect 579554 292170 579622 292226
rect 579678 292170 596496 292226
rect 596552 292170 596620 292226
rect 596676 292170 596744 292226
rect 596800 292170 596868 292226
rect 596924 292170 597980 292226
rect -1916 292102 597980 292170
rect -1916 292046 -860 292102
rect -804 292046 -736 292102
rect -680 292046 -612 292102
rect -556 292046 -488 292102
rect -432 292046 3250 292102
rect 3306 292046 3374 292102
rect 3430 292046 3498 292102
rect 3554 292046 3622 292102
rect 3678 292046 201250 292102
rect 201306 292046 201374 292102
rect 201430 292046 201498 292102
rect 201554 292046 201622 292102
rect 201678 292046 381250 292102
rect 381306 292046 381374 292102
rect 381430 292046 381498 292102
rect 381554 292046 381622 292102
rect 381678 292046 399250 292102
rect 399306 292046 399374 292102
rect 399430 292046 399498 292102
rect 399554 292046 399622 292102
rect 399678 292046 579250 292102
rect 579306 292046 579374 292102
rect 579430 292046 579498 292102
rect 579554 292046 579622 292102
rect 579678 292046 596496 292102
rect 596552 292046 596620 292102
rect 596676 292046 596744 292102
rect 596800 292046 596868 292102
rect 596924 292046 597980 292102
rect -1916 291978 597980 292046
rect -1916 291922 -860 291978
rect -804 291922 -736 291978
rect -680 291922 -612 291978
rect -556 291922 -488 291978
rect -432 291922 3250 291978
rect 3306 291922 3374 291978
rect 3430 291922 3498 291978
rect 3554 291922 3622 291978
rect 3678 291922 201250 291978
rect 201306 291922 201374 291978
rect 201430 291922 201498 291978
rect 201554 291922 201622 291978
rect 201678 291922 381250 291978
rect 381306 291922 381374 291978
rect 381430 291922 381498 291978
rect 381554 291922 381622 291978
rect 381678 291922 399250 291978
rect 399306 291922 399374 291978
rect 399430 291922 399498 291978
rect 399554 291922 399622 291978
rect 399678 291922 579250 291978
rect 579306 291922 579374 291978
rect 579430 291922 579498 291978
rect 579554 291922 579622 291978
rect 579678 291922 596496 291978
rect 596552 291922 596620 291978
rect 596676 291922 596744 291978
rect 596800 291922 596868 291978
rect 596924 291922 597980 291978
rect -1916 291826 597980 291922
rect -1916 280350 597980 280446
rect -1916 280294 -1820 280350
rect -1764 280294 -1696 280350
rect -1640 280294 -1572 280350
rect -1516 280294 -1448 280350
rect -1392 280294 6970 280350
rect 7026 280294 7094 280350
rect 7150 280294 7218 280350
rect 7274 280294 7342 280350
rect 7398 280294 204970 280350
rect 205026 280294 205094 280350
rect 205150 280294 205218 280350
rect 205274 280294 205342 280350
rect 205398 280294 384970 280350
rect 385026 280294 385094 280350
rect 385150 280294 385218 280350
rect 385274 280294 385342 280350
rect 385398 280294 402970 280350
rect 403026 280294 403094 280350
rect 403150 280294 403218 280350
rect 403274 280294 403342 280350
rect 403398 280294 582970 280350
rect 583026 280294 583094 280350
rect 583150 280294 583218 280350
rect 583274 280294 583342 280350
rect 583398 280294 597456 280350
rect 597512 280294 597580 280350
rect 597636 280294 597704 280350
rect 597760 280294 597828 280350
rect 597884 280294 597980 280350
rect -1916 280226 597980 280294
rect -1916 280170 -1820 280226
rect -1764 280170 -1696 280226
rect -1640 280170 -1572 280226
rect -1516 280170 -1448 280226
rect -1392 280170 6970 280226
rect 7026 280170 7094 280226
rect 7150 280170 7218 280226
rect 7274 280170 7342 280226
rect 7398 280170 204970 280226
rect 205026 280170 205094 280226
rect 205150 280170 205218 280226
rect 205274 280170 205342 280226
rect 205398 280170 384970 280226
rect 385026 280170 385094 280226
rect 385150 280170 385218 280226
rect 385274 280170 385342 280226
rect 385398 280170 402970 280226
rect 403026 280170 403094 280226
rect 403150 280170 403218 280226
rect 403274 280170 403342 280226
rect 403398 280170 582970 280226
rect 583026 280170 583094 280226
rect 583150 280170 583218 280226
rect 583274 280170 583342 280226
rect 583398 280170 597456 280226
rect 597512 280170 597580 280226
rect 597636 280170 597704 280226
rect 597760 280170 597828 280226
rect 597884 280170 597980 280226
rect -1916 280102 597980 280170
rect -1916 280046 -1820 280102
rect -1764 280046 -1696 280102
rect -1640 280046 -1572 280102
rect -1516 280046 -1448 280102
rect -1392 280046 6970 280102
rect 7026 280046 7094 280102
rect 7150 280046 7218 280102
rect 7274 280046 7342 280102
rect 7398 280046 204970 280102
rect 205026 280046 205094 280102
rect 205150 280046 205218 280102
rect 205274 280046 205342 280102
rect 205398 280046 384970 280102
rect 385026 280046 385094 280102
rect 385150 280046 385218 280102
rect 385274 280046 385342 280102
rect 385398 280046 402970 280102
rect 403026 280046 403094 280102
rect 403150 280046 403218 280102
rect 403274 280046 403342 280102
rect 403398 280046 582970 280102
rect 583026 280046 583094 280102
rect 583150 280046 583218 280102
rect 583274 280046 583342 280102
rect 583398 280046 597456 280102
rect 597512 280046 597580 280102
rect 597636 280046 597704 280102
rect 597760 280046 597828 280102
rect 597884 280046 597980 280102
rect -1916 279978 597980 280046
rect -1916 279922 -1820 279978
rect -1764 279922 -1696 279978
rect -1640 279922 -1572 279978
rect -1516 279922 -1448 279978
rect -1392 279922 6970 279978
rect 7026 279922 7094 279978
rect 7150 279922 7218 279978
rect 7274 279922 7342 279978
rect 7398 279922 204970 279978
rect 205026 279922 205094 279978
rect 205150 279922 205218 279978
rect 205274 279922 205342 279978
rect 205398 279922 384970 279978
rect 385026 279922 385094 279978
rect 385150 279922 385218 279978
rect 385274 279922 385342 279978
rect 385398 279922 402970 279978
rect 403026 279922 403094 279978
rect 403150 279922 403218 279978
rect 403274 279922 403342 279978
rect 403398 279922 582970 279978
rect 583026 279922 583094 279978
rect 583150 279922 583218 279978
rect 583274 279922 583342 279978
rect 583398 279922 597456 279978
rect 597512 279922 597580 279978
rect 597636 279922 597704 279978
rect 597760 279922 597828 279978
rect 597884 279922 597980 279978
rect -1916 279826 597980 279922
rect -1916 274350 597980 274446
rect -1916 274294 -860 274350
rect -804 274294 -736 274350
rect -680 274294 -612 274350
rect -556 274294 -488 274350
rect -432 274294 3250 274350
rect 3306 274294 3374 274350
rect 3430 274294 3498 274350
rect 3554 274294 3622 274350
rect 3678 274294 201250 274350
rect 201306 274294 201374 274350
rect 201430 274294 201498 274350
rect 201554 274294 201622 274350
rect 201678 274294 381250 274350
rect 381306 274294 381374 274350
rect 381430 274294 381498 274350
rect 381554 274294 381622 274350
rect 381678 274294 399250 274350
rect 399306 274294 399374 274350
rect 399430 274294 399498 274350
rect 399554 274294 399622 274350
rect 399678 274294 579250 274350
rect 579306 274294 579374 274350
rect 579430 274294 579498 274350
rect 579554 274294 579622 274350
rect 579678 274294 596496 274350
rect 596552 274294 596620 274350
rect 596676 274294 596744 274350
rect 596800 274294 596868 274350
rect 596924 274294 597980 274350
rect -1916 274226 597980 274294
rect -1916 274170 -860 274226
rect -804 274170 -736 274226
rect -680 274170 -612 274226
rect -556 274170 -488 274226
rect -432 274170 3250 274226
rect 3306 274170 3374 274226
rect 3430 274170 3498 274226
rect 3554 274170 3622 274226
rect 3678 274170 201250 274226
rect 201306 274170 201374 274226
rect 201430 274170 201498 274226
rect 201554 274170 201622 274226
rect 201678 274170 381250 274226
rect 381306 274170 381374 274226
rect 381430 274170 381498 274226
rect 381554 274170 381622 274226
rect 381678 274170 399250 274226
rect 399306 274170 399374 274226
rect 399430 274170 399498 274226
rect 399554 274170 399622 274226
rect 399678 274170 579250 274226
rect 579306 274170 579374 274226
rect 579430 274170 579498 274226
rect 579554 274170 579622 274226
rect 579678 274170 596496 274226
rect 596552 274170 596620 274226
rect 596676 274170 596744 274226
rect 596800 274170 596868 274226
rect 596924 274170 597980 274226
rect -1916 274102 597980 274170
rect -1916 274046 -860 274102
rect -804 274046 -736 274102
rect -680 274046 -612 274102
rect -556 274046 -488 274102
rect -432 274046 3250 274102
rect 3306 274046 3374 274102
rect 3430 274046 3498 274102
rect 3554 274046 3622 274102
rect 3678 274046 201250 274102
rect 201306 274046 201374 274102
rect 201430 274046 201498 274102
rect 201554 274046 201622 274102
rect 201678 274046 381250 274102
rect 381306 274046 381374 274102
rect 381430 274046 381498 274102
rect 381554 274046 381622 274102
rect 381678 274046 399250 274102
rect 399306 274046 399374 274102
rect 399430 274046 399498 274102
rect 399554 274046 399622 274102
rect 399678 274046 579250 274102
rect 579306 274046 579374 274102
rect 579430 274046 579498 274102
rect 579554 274046 579622 274102
rect 579678 274046 596496 274102
rect 596552 274046 596620 274102
rect 596676 274046 596744 274102
rect 596800 274046 596868 274102
rect 596924 274046 597980 274102
rect -1916 273978 597980 274046
rect -1916 273922 -860 273978
rect -804 273922 -736 273978
rect -680 273922 -612 273978
rect -556 273922 -488 273978
rect -432 273922 3250 273978
rect 3306 273922 3374 273978
rect 3430 273922 3498 273978
rect 3554 273922 3622 273978
rect 3678 273922 201250 273978
rect 201306 273922 201374 273978
rect 201430 273922 201498 273978
rect 201554 273922 201622 273978
rect 201678 273922 381250 273978
rect 381306 273922 381374 273978
rect 381430 273922 381498 273978
rect 381554 273922 381622 273978
rect 381678 273922 399250 273978
rect 399306 273922 399374 273978
rect 399430 273922 399498 273978
rect 399554 273922 399622 273978
rect 399678 273922 579250 273978
rect 579306 273922 579374 273978
rect 579430 273922 579498 273978
rect 579554 273922 579622 273978
rect 579678 273922 596496 273978
rect 596552 273922 596620 273978
rect 596676 273922 596744 273978
rect 596800 273922 596868 273978
rect 596924 273922 597980 273978
rect -1916 273826 597980 273922
rect -1916 262350 597980 262446
rect -1916 262294 -1820 262350
rect -1764 262294 -1696 262350
rect -1640 262294 -1572 262350
rect -1516 262294 -1448 262350
rect -1392 262294 6970 262350
rect 7026 262294 7094 262350
rect 7150 262294 7218 262350
rect 7274 262294 7342 262350
rect 7398 262294 204970 262350
rect 205026 262294 205094 262350
rect 205150 262294 205218 262350
rect 205274 262294 205342 262350
rect 205398 262294 384970 262350
rect 385026 262294 385094 262350
rect 385150 262294 385218 262350
rect 385274 262294 385342 262350
rect 385398 262294 402970 262350
rect 403026 262294 403094 262350
rect 403150 262294 403218 262350
rect 403274 262294 403342 262350
rect 403398 262294 582970 262350
rect 583026 262294 583094 262350
rect 583150 262294 583218 262350
rect 583274 262294 583342 262350
rect 583398 262294 597456 262350
rect 597512 262294 597580 262350
rect 597636 262294 597704 262350
rect 597760 262294 597828 262350
rect 597884 262294 597980 262350
rect -1916 262226 597980 262294
rect -1916 262170 -1820 262226
rect -1764 262170 -1696 262226
rect -1640 262170 -1572 262226
rect -1516 262170 -1448 262226
rect -1392 262170 6970 262226
rect 7026 262170 7094 262226
rect 7150 262170 7218 262226
rect 7274 262170 7342 262226
rect 7398 262170 204970 262226
rect 205026 262170 205094 262226
rect 205150 262170 205218 262226
rect 205274 262170 205342 262226
rect 205398 262170 384970 262226
rect 385026 262170 385094 262226
rect 385150 262170 385218 262226
rect 385274 262170 385342 262226
rect 385398 262170 402970 262226
rect 403026 262170 403094 262226
rect 403150 262170 403218 262226
rect 403274 262170 403342 262226
rect 403398 262170 582970 262226
rect 583026 262170 583094 262226
rect 583150 262170 583218 262226
rect 583274 262170 583342 262226
rect 583398 262170 597456 262226
rect 597512 262170 597580 262226
rect 597636 262170 597704 262226
rect 597760 262170 597828 262226
rect 597884 262170 597980 262226
rect -1916 262102 597980 262170
rect -1916 262046 -1820 262102
rect -1764 262046 -1696 262102
rect -1640 262046 -1572 262102
rect -1516 262046 -1448 262102
rect -1392 262046 6970 262102
rect 7026 262046 7094 262102
rect 7150 262046 7218 262102
rect 7274 262046 7342 262102
rect 7398 262046 204970 262102
rect 205026 262046 205094 262102
rect 205150 262046 205218 262102
rect 205274 262046 205342 262102
rect 205398 262046 384970 262102
rect 385026 262046 385094 262102
rect 385150 262046 385218 262102
rect 385274 262046 385342 262102
rect 385398 262046 402970 262102
rect 403026 262046 403094 262102
rect 403150 262046 403218 262102
rect 403274 262046 403342 262102
rect 403398 262046 582970 262102
rect 583026 262046 583094 262102
rect 583150 262046 583218 262102
rect 583274 262046 583342 262102
rect 583398 262046 597456 262102
rect 597512 262046 597580 262102
rect 597636 262046 597704 262102
rect 597760 262046 597828 262102
rect 597884 262046 597980 262102
rect -1916 261978 597980 262046
rect -1916 261922 -1820 261978
rect -1764 261922 -1696 261978
rect -1640 261922 -1572 261978
rect -1516 261922 -1448 261978
rect -1392 261922 6970 261978
rect 7026 261922 7094 261978
rect 7150 261922 7218 261978
rect 7274 261922 7342 261978
rect 7398 261922 204970 261978
rect 205026 261922 205094 261978
rect 205150 261922 205218 261978
rect 205274 261922 205342 261978
rect 205398 261922 384970 261978
rect 385026 261922 385094 261978
rect 385150 261922 385218 261978
rect 385274 261922 385342 261978
rect 385398 261922 402970 261978
rect 403026 261922 403094 261978
rect 403150 261922 403218 261978
rect 403274 261922 403342 261978
rect 403398 261922 582970 261978
rect 583026 261922 583094 261978
rect 583150 261922 583218 261978
rect 583274 261922 583342 261978
rect 583398 261922 597456 261978
rect 597512 261922 597580 261978
rect 597636 261922 597704 261978
rect 597760 261922 597828 261978
rect 597884 261922 597980 261978
rect -1916 261826 597980 261922
rect -1916 256350 597980 256446
rect -1916 256294 -860 256350
rect -804 256294 -736 256350
rect -680 256294 -612 256350
rect -556 256294 -488 256350
rect -432 256294 3250 256350
rect 3306 256294 3374 256350
rect 3430 256294 3498 256350
rect 3554 256294 3622 256350
rect 3678 256294 201250 256350
rect 201306 256294 201374 256350
rect 201430 256294 201498 256350
rect 201554 256294 201622 256350
rect 201678 256294 381250 256350
rect 381306 256294 381374 256350
rect 381430 256294 381498 256350
rect 381554 256294 381622 256350
rect 381678 256294 399250 256350
rect 399306 256294 399374 256350
rect 399430 256294 399498 256350
rect 399554 256294 399622 256350
rect 399678 256294 579250 256350
rect 579306 256294 579374 256350
rect 579430 256294 579498 256350
rect 579554 256294 579622 256350
rect 579678 256294 596496 256350
rect 596552 256294 596620 256350
rect 596676 256294 596744 256350
rect 596800 256294 596868 256350
rect 596924 256294 597980 256350
rect -1916 256226 597980 256294
rect -1916 256170 -860 256226
rect -804 256170 -736 256226
rect -680 256170 -612 256226
rect -556 256170 -488 256226
rect -432 256170 3250 256226
rect 3306 256170 3374 256226
rect 3430 256170 3498 256226
rect 3554 256170 3622 256226
rect 3678 256170 201250 256226
rect 201306 256170 201374 256226
rect 201430 256170 201498 256226
rect 201554 256170 201622 256226
rect 201678 256170 381250 256226
rect 381306 256170 381374 256226
rect 381430 256170 381498 256226
rect 381554 256170 381622 256226
rect 381678 256170 399250 256226
rect 399306 256170 399374 256226
rect 399430 256170 399498 256226
rect 399554 256170 399622 256226
rect 399678 256170 579250 256226
rect 579306 256170 579374 256226
rect 579430 256170 579498 256226
rect 579554 256170 579622 256226
rect 579678 256170 596496 256226
rect 596552 256170 596620 256226
rect 596676 256170 596744 256226
rect 596800 256170 596868 256226
rect 596924 256170 597980 256226
rect -1916 256102 597980 256170
rect -1916 256046 -860 256102
rect -804 256046 -736 256102
rect -680 256046 -612 256102
rect -556 256046 -488 256102
rect -432 256046 3250 256102
rect 3306 256046 3374 256102
rect 3430 256046 3498 256102
rect 3554 256046 3622 256102
rect 3678 256046 201250 256102
rect 201306 256046 201374 256102
rect 201430 256046 201498 256102
rect 201554 256046 201622 256102
rect 201678 256046 381250 256102
rect 381306 256046 381374 256102
rect 381430 256046 381498 256102
rect 381554 256046 381622 256102
rect 381678 256046 399250 256102
rect 399306 256046 399374 256102
rect 399430 256046 399498 256102
rect 399554 256046 399622 256102
rect 399678 256046 579250 256102
rect 579306 256046 579374 256102
rect 579430 256046 579498 256102
rect 579554 256046 579622 256102
rect 579678 256046 596496 256102
rect 596552 256046 596620 256102
rect 596676 256046 596744 256102
rect 596800 256046 596868 256102
rect 596924 256046 597980 256102
rect -1916 255978 597980 256046
rect -1916 255922 -860 255978
rect -804 255922 -736 255978
rect -680 255922 -612 255978
rect -556 255922 -488 255978
rect -432 255922 3250 255978
rect 3306 255922 3374 255978
rect 3430 255922 3498 255978
rect 3554 255922 3622 255978
rect 3678 255922 201250 255978
rect 201306 255922 201374 255978
rect 201430 255922 201498 255978
rect 201554 255922 201622 255978
rect 201678 255922 381250 255978
rect 381306 255922 381374 255978
rect 381430 255922 381498 255978
rect 381554 255922 381622 255978
rect 381678 255922 399250 255978
rect 399306 255922 399374 255978
rect 399430 255922 399498 255978
rect 399554 255922 399622 255978
rect 399678 255922 579250 255978
rect 579306 255922 579374 255978
rect 579430 255922 579498 255978
rect 579554 255922 579622 255978
rect 579678 255922 596496 255978
rect 596552 255922 596620 255978
rect 596676 255922 596744 255978
rect 596800 255922 596868 255978
rect 596924 255922 597980 255978
rect -1916 255826 597980 255922
rect -1916 244350 597980 244446
rect -1916 244294 -1820 244350
rect -1764 244294 -1696 244350
rect -1640 244294 -1572 244350
rect -1516 244294 -1448 244350
rect -1392 244294 6970 244350
rect 7026 244294 7094 244350
rect 7150 244294 7218 244350
rect 7274 244294 7342 244350
rect 7398 244294 204970 244350
rect 205026 244294 205094 244350
rect 205150 244294 205218 244350
rect 205274 244294 205342 244350
rect 205398 244294 384970 244350
rect 385026 244294 385094 244350
rect 385150 244294 385218 244350
rect 385274 244294 385342 244350
rect 385398 244294 402970 244350
rect 403026 244294 403094 244350
rect 403150 244294 403218 244350
rect 403274 244294 403342 244350
rect 403398 244294 582970 244350
rect 583026 244294 583094 244350
rect 583150 244294 583218 244350
rect 583274 244294 583342 244350
rect 583398 244294 597456 244350
rect 597512 244294 597580 244350
rect 597636 244294 597704 244350
rect 597760 244294 597828 244350
rect 597884 244294 597980 244350
rect -1916 244226 597980 244294
rect -1916 244170 -1820 244226
rect -1764 244170 -1696 244226
rect -1640 244170 -1572 244226
rect -1516 244170 -1448 244226
rect -1392 244170 6970 244226
rect 7026 244170 7094 244226
rect 7150 244170 7218 244226
rect 7274 244170 7342 244226
rect 7398 244170 204970 244226
rect 205026 244170 205094 244226
rect 205150 244170 205218 244226
rect 205274 244170 205342 244226
rect 205398 244170 384970 244226
rect 385026 244170 385094 244226
rect 385150 244170 385218 244226
rect 385274 244170 385342 244226
rect 385398 244170 402970 244226
rect 403026 244170 403094 244226
rect 403150 244170 403218 244226
rect 403274 244170 403342 244226
rect 403398 244170 582970 244226
rect 583026 244170 583094 244226
rect 583150 244170 583218 244226
rect 583274 244170 583342 244226
rect 583398 244170 597456 244226
rect 597512 244170 597580 244226
rect 597636 244170 597704 244226
rect 597760 244170 597828 244226
rect 597884 244170 597980 244226
rect -1916 244102 597980 244170
rect -1916 244046 -1820 244102
rect -1764 244046 -1696 244102
rect -1640 244046 -1572 244102
rect -1516 244046 -1448 244102
rect -1392 244046 6970 244102
rect 7026 244046 7094 244102
rect 7150 244046 7218 244102
rect 7274 244046 7342 244102
rect 7398 244046 204970 244102
rect 205026 244046 205094 244102
rect 205150 244046 205218 244102
rect 205274 244046 205342 244102
rect 205398 244046 384970 244102
rect 385026 244046 385094 244102
rect 385150 244046 385218 244102
rect 385274 244046 385342 244102
rect 385398 244046 402970 244102
rect 403026 244046 403094 244102
rect 403150 244046 403218 244102
rect 403274 244046 403342 244102
rect 403398 244046 582970 244102
rect 583026 244046 583094 244102
rect 583150 244046 583218 244102
rect 583274 244046 583342 244102
rect 583398 244046 597456 244102
rect 597512 244046 597580 244102
rect 597636 244046 597704 244102
rect 597760 244046 597828 244102
rect 597884 244046 597980 244102
rect -1916 243978 597980 244046
rect -1916 243922 -1820 243978
rect -1764 243922 -1696 243978
rect -1640 243922 -1572 243978
rect -1516 243922 -1448 243978
rect -1392 243922 6970 243978
rect 7026 243922 7094 243978
rect 7150 243922 7218 243978
rect 7274 243922 7342 243978
rect 7398 243922 204970 243978
rect 205026 243922 205094 243978
rect 205150 243922 205218 243978
rect 205274 243922 205342 243978
rect 205398 243922 384970 243978
rect 385026 243922 385094 243978
rect 385150 243922 385218 243978
rect 385274 243922 385342 243978
rect 385398 243922 402970 243978
rect 403026 243922 403094 243978
rect 403150 243922 403218 243978
rect 403274 243922 403342 243978
rect 403398 243922 582970 243978
rect 583026 243922 583094 243978
rect 583150 243922 583218 243978
rect 583274 243922 583342 243978
rect 583398 243922 597456 243978
rect 597512 243922 597580 243978
rect 597636 243922 597704 243978
rect 597760 243922 597828 243978
rect 597884 243922 597980 243978
rect -1916 243826 597980 243922
rect -1916 238350 597980 238446
rect -1916 238294 -860 238350
rect -804 238294 -736 238350
rect -680 238294 -612 238350
rect -556 238294 -488 238350
rect -432 238294 3250 238350
rect 3306 238294 3374 238350
rect 3430 238294 3498 238350
rect 3554 238294 3622 238350
rect 3678 238294 201250 238350
rect 201306 238294 201374 238350
rect 201430 238294 201498 238350
rect 201554 238294 201622 238350
rect 201678 238294 381250 238350
rect 381306 238294 381374 238350
rect 381430 238294 381498 238350
rect 381554 238294 381622 238350
rect 381678 238294 399250 238350
rect 399306 238294 399374 238350
rect 399430 238294 399498 238350
rect 399554 238294 399622 238350
rect 399678 238294 579250 238350
rect 579306 238294 579374 238350
rect 579430 238294 579498 238350
rect 579554 238294 579622 238350
rect 579678 238294 596496 238350
rect 596552 238294 596620 238350
rect 596676 238294 596744 238350
rect 596800 238294 596868 238350
rect 596924 238294 597980 238350
rect -1916 238226 597980 238294
rect -1916 238170 -860 238226
rect -804 238170 -736 238226
rect -680 238170 -612 238226
rect -556 238170 -488 238226
rect -432 238170 3250 238226
rect 3306 238170 3374 238226
rect 3430 238170 3498 238226
rect 3554 238170 3622 238226
rect 3678 238170 201250 238226
rect 201306 238170 201374 238226
rect 201430 238170 201498 238226
rect 201554 238170 201622 238226
rect 201678 238170 381250 238226
rect 381306 238170 381374 238226
rect 381430 238170 381498 238226
rect 381554 238170 381622 238226
rect 381678 238170 399250 238226
rect 399306 238170 399374 238226
rect 399430 238170 399498 238226
rect 399554 238170 399622 238226
rect 399678 238170 579250 238226
rect 579306 238170 579374 238226
rect 579430 238170 579498 238226
rect 579554 238170 579622 238226
rect 579678 238170 596496 238226
rect 596552 238170 596620 238226
rect 596676 238170 596744 238226
rect 596800 238170 596868 238226
rect 596924 238170 597980 238226
rect -1916 238102 597980 238170
rect -1916 238046 -860 238102
rect -804 238046 -736 238102
rect -680 238046 -612 238102
rect -556 238046 -488 238102
rect -432 238046 3250 238102
rect 3306 238046 3374 238102
rect 3430 238046 3498 238102
rect 3554 238046 3622 238102
rect 3678 238046 201250 238102
rect 201306 238046 201374 238102
rect 201430 238046 201498 238102
rect 201554 238046 201622 238102
rect 201678 238046 381250 238102
rect 381306 238046 381374 238102
rect 381430 238046 381498 238102
rect 381554 238046 381622 238102
rect 381678 238046 399250 238102
rect 399306 238046 399374 238102
rect 399430 238046 399498 238102
rect 399554 238046 399622 238102
rect 399678 238046 579250 238102
rect 579306 238046 579374 238102
rect 579430 238046 579498 238102
rect 579554 238046 579622 238102
rect 579678 238046 596496 238102
rect 596552 238046 596620 238102
rect 596676 238046 596744 238102
rect 596800 238046 596868 238102
rect 596924 238046 597980 238102
rect -1916 237978 597980 238046
rect -1916 237922 -860 237978
rect -804 237922 -736 237978
rect -680 237922 -612 237978
rect -556 237922 -488 237978
rect -432 237922 3250 237978
rect 3306 237922 3374 237978
rect 3430 237922 3498 237978
rect 3554 237922 3622 237978
rect 3678 237922 201250 237978
rect 201306 237922 201374 237978
rect 201430 237922 201498 237978
rect 201554 237922 201622 237978
rect 201678 237922 381250 237978
rect 381306 237922 381374 237978
rect 381430 237922 381498 237978
rect 381554 237922 381622 237978
rect 381678 237922 399250 237978
rect 399306 237922 399374 237978
rect 399430 237922 399498 237978
rect 399554 237922 399622 237978
rect 399678 237922 579250 237978
rect 579306 237922 579374 237978
rect 579430 237922 579498 237978
rect 579554 237922 579622 237978
rect 579678 237922 596496 237978
rect 596552 237922 596620 237978
rect 596676 237922 596744 237978
rect 596800 237922 596868 237978
rect 596924 237922 597980 237978
rect -1916 237826 597980 237922
rect -1916 226350 597980 226446
rect -1916 226294 -1820 226350
rect -1764 226294 -1696 226350
rect -1640 226294 -1572 226350
rect -1516 226294 -1448 226350
rect -1392 226294 6970 226350
rect 7026 226294 7094 226350
rect 7150 226294 7218 226350
rect 7274 226294 7342 226350
rect 7398 226294 204970 226350
rect 205026 226294 205094 226350
rect 205150 226294 205218 226350
rect 205274 226294 205342 226350
rect 205398 226294 384970 226350
rect 385026 226294 385094 226350
rect 385150 226294 385218 226350
rect 385274 226294 385342 226350
rect 385398 226294 402970 226350
rect 403026 226294 403094 226350
rect 403150 226294 403218 226350
rect 403274 226294 403342 226350
rect 403398 226294 582970 226350
rect 583026 226294 583094 226350
rect 583150 226294 583218 226350
rect 583274 226294 583342 226350
rect 583398 226294 597456 226350
rect 597512 226294 597580 226350
rect 597636 226294 597704 226350
rect 597760 226294 597828 226350
rect 597884 226294 597980 226350
rect -1916 226226 597980 226294
rect -1916 226170 -1820 226226
rect -1764 226170 -1696 226226
rect -1640 226170 -1572 226226
rect -1516 226170 -1448 226226
rect -1392 226170 6970 226226
rect 7026 226170 7094 226226
rect 7150 226170 7218 226226
rect 7274 226170 7342 226226
rect 7398 226170 204970 226226
rect 205026 226170 205094 226226
rect 205150 226170 205218 226226
rect 205274 226170 205342 226226
rect 205398 226170 384970 226226
rect 385026 226170 385094 226226
rect 385150 226170 385218 226226
rect 385274 226170 385342 226226
rect 385398 226170 402970 226226
rect 403026 226170 403094 226226
rect 403150 226170 403218 226226
rect 403274 226170 403342 226226
rect 403398 226170 582970 226226
rect 583026 226170 583094 226226
rect 583150 226170 583218 226226
rect 583274 226170 583342 226226
rect 583398 226170 597456 226226
rect 597512 226170 597580 226226
rect 597636 226170 597704 226226
rect 597760 226170 597828 226226
rect 597884 226170 597980 226226
rect -1916 226102 597980 226170
rect -1916 226046 -1820 226102
rect -1764 226046 -1696 226102
rect -1640 226046 -1572 226102
rect -1516 226046 -1448 226102
rect -1392 226046 6970 226102
rect 7026 226046 7094 226102
rect 7150 226046 7218 226102
rect 7274 226046 7342 226102
rect 7398 226046 204970 226102
rect 205026 226046 205094 226102
rect 205150 226046 205218 226102
rect 205274 226046 205342 226102
rect 205398 226046 384970 226102
rect 385026 226046 385094 226102
rect 385150 226046 385218 226102
rect 385274 226046 385342 226102
rect 385398 226046 402970 226102
rect 403026 226046 403094 226102
rect 403150 226046 403218 226102
rect 403274 226046 403342 226102
rect 403398 226046 582970 226102
rect 583026 226046 583094 226102
rect 583150 226046 583218 226102
rect 583274 226046 583342 226102
rect 583398 226046 597456 226102
rect 597512 226046 597580 226102
rect 597636 226046 597704 226102
rect 597760 226046 597828 226102
rect 597884 226046 597980 226102
rect -1916 225978 597980 226046
rect -1916 225922 -1820 225978
rect -1764 225922 -1696 225978
rect -1640 225922 -1572 225978
rect -1516 225922 -1448 225978
rect -1392 225922 6970 225978
rect 7026 225922 7094 225978
rect 7150 225922 7218 225978
rect 7274 225922 7342 225978
rect 7398 225922 204970 225978
rect 205026 225922 205094 225978
rect 205150 225922 205218 225978
rect 205274 225922 205342 225978
rect 205398 225922 384970 225978
rect 385026 225922 385094 225978
rect 385150 225922 385218 225978
rect 385274 225922 385342 225978
rect 385398 225922 402970 225978
rect 403026 225922 403094 225978
rect 403150 225922 403218 225978
rect 403274 225922 403342 225978
rect 403398 225922 582970 225978
rect 583026 225922 583094 225978
rect 583150 225922 583218 225978
rect 583274 225922 583342 225978
rect 583398 225922 597456 225978
rect 597512 225922 597580 225978
rect 597636 225922 597704 225978
rect 597760 225922 597828 225978
rect 597884 225922 597980 225978
rect -1916 225826 597980 225922
rect -1916 220350 597980 220446
rect -1916 220294 -860 220350
rect -804 220294 -736 220350
rect -680 220294 -612 220350
rect -556 220294 -488 220350
rect -432 220294 3250 220350
rect 3306 220294 3374 220350
rect 3430 220294 3498 220350
rect 3554 220294 3622 220350
rect 3678 220294 201250 220350
rect 201306 220294 201374 220350
rect 201430 220294 201498 220350
rect 201554 220294 201622 220350
rect 201678 220294 381250 220350
rect 381306 220294 381374 220350
rect 381430 220294 381498 220350
rect 381554 220294 381622 220350
rect 381678 220294 399250 220350
rect 399306 220294 399374 220350
rect 399430 220294 399498 220350
rect 399554 220294 399622 220350
rect 399678 220294 579250 220350
rect 579306 220294 579374 220350
rect 579430 220294 579498 220350
rect 579554 220294 579622 220350
rect 579678 220294 596496 220350
rect 596552 220294 596620 220350
rect 596676 220294 596744 220350
rect 596800 220294 596868 220350
rect 596924 220294 597980 220350
rect -1916 220226 597980 220294
rect -1916 220170 -860 220226
rect -804 220170 -736 220226
rect -680 220170 -612 220226
rect -556 220170 -488 220226
rect -432 220170 3250 220226
rect 3306 220170 3374 220226
rect 3430 220170 3498 220226
rect 3554 220170 3622 220226
rect 3678 220170 201250 220226
rect 201306 220170 201374 220226
rect 201430 220170 201498 220226
rect 201554 220170 201622 220226
rect 201678 220170 381250 220226
rect 381306 220170 381374 220226
rect 381430 220170 381498 220226
rect 381554 220170 381622 220226
rect 381678 220170 399250 220226
rect 399306 220170 399374 220226
rect 399430 220170 399498 220226
rect 399554 220170 399622 220226
rect 399678 220170 579250 220226
rect 579306 220170 579374 220226
rect 579430 220170 579498 220226
rect 579554 220170 579622 220226
rect 579678 220170 596496 220226
rect 596552 220170 596620 220226
rect 596676 220170 596744 220226
rect 596800 220170 596868 220226
rect 596924 220170 597980 220226
rect -1916 220102 597980 220170
rect -1916 220046 -860 220102
rect -804 220046 -736 220102
rect -680 220046 -612 220102
rect -556 220046 -488 220102
rect -432 220046 3250 220102
rect 3306 220046 3374 220102
rect 3430 220046 3498 220102
rect 3554 220046 3622 220102
rect 3678 220046 201250 220102
rect 201306 220046 201374 220102
rect 201430 220046 201498 220102
rect 201554 220046 201622 220102
rect 201678 220046 381250 220102
rect 381306 220046 381374 220102
rect 381430 220046 381498 220102
rect 381554 220046 381622 220102
rect 381678 220046 399250 220102
rect 399306 220046 399374 220102
rect 399430 220046 399498 220102
rect 399554 220046 399622 220102
rect 399678 220046 579250 220102
rect 579306 220046 579374 220102
rect 579430 220046 579498 220102
rect 579554 220046 579622 220102
rect 579678 220046 596496 220102
rect 596552 220046 596620 220102
rect 596676 220046 596744 220102
rect 596800 220046 596868 220102
rect 596924 220046 597980 220102
rect -1916 219978 597980 220046
rect -1916 219922 -860 219978
rect -804 219922 -736 219978
rect -680 219922 -612 219978
rect -556 219922 -488 219978
rect -432 219922 3250 219978
rect 3306 219922 3374 219978
rect 3430 219922 3498 219978
rect 3554 219922 3622 219978
rect 3678 219922 201250 219978
rect 201306 219922 201374 219978
rect 201430 219922 201498 219978
rect 201554 219922 201622 219978
rect 201678 219922 381250 219978
rect 381306 219922 381374 219978
rect 381430 219922 381498 219978
rect 381554 219922 381622 219978
rect 381678 219922 399250 219978
rect 399306 219922 399374 219978
rect 399430 219922 399498 219978
rect 399554 219922 399622 219978
rect 399678 219922 579250 219978
rect 579306 219922 579374 219978
rect 579430 219922 579498 219978
rect 579554 219922 579622 219978
rect 579678 219922 596496 219978
rect 596552 219922 596620 219978
rect 596676 219922 596744 219978
rect 596800 219922 596868 219978
rect 596924 219922 597980 219978
rect -1916 219826 597980 219922
rect -1916 208350 597980 208446
rect -1916 208294 -1820 208350
rect -1764 208294 -1696 208350
rect -1640 208294 -1572 208350
rect -1516 208294 -1448 208350
rect -1392 208294 6970 208350
rect 7026 208294 7094 208350
rect 7150 208294 7218 208350
rect 7274 208294 7342 208350
rect 7398 208294 204970 208350
rect 205026 208294 205094 208350
rect 205150 208294 205218 208350
rect 205274 208294 205342 208350
rect 205398 208294 384970 208350
rect 385026 208294 385094 208350
rect 385150 208294 385218 208350
rect 385274 208294 385342 208350
rect 385398 208294 402970 208350
rect 403026 208294 403094 208350
rect 403150 208294 403218 208350
rect 403274 208294 403342 208350
rect 403398 208294 582970 208350
rect 583026 208294 583094 208350
rect 583150 208294 583218 208350
rect 583274 208294 583342 208350
rect 583398 208294 597456 208350
rect 597512 208294 597580 208350
rect 597636 208294 597704 208350
rect 597760 208294 597828 208350
rect 597884 208294 597980 208350
rect -1916 208226 597980 208294
rect -1916 208170 -1820 208226
rect -1764 208170 -1696 208226
rect -1640 208170 -1572 208226
rect -1516 208170 -1448 208226
rect -1392 208170 6970 208226
rect 7026 208170 7094 208226
rect 7150 208170 7218 208226
rect 7274 208170 7342 208226
rect 7398 208170 204970 208226
rect 205026 208170 205094 208226
rect 205150 208170 205218 208226
rect 205274 208170 205342 208226
rect 205398 208170 384970 208226
rect 385026 208170 385094 208226
rect 385150 208170 385218 208226
rect 385274 208170 385342 208226
rect 385398 208170 402970 208226
rect 403026 208170 403094 208226
rect 403150 208170 403218 208226
rect 403274 208170 403342 208226
rect 403398 208170 582970 208226
rect 583026 208170 583094 208226
rect 583150 208170 583218 208226
rect 583274 208170 583342 208226
rect 583398 208170 597456 208226
rect 597512 208170 597580 208226
rect 597636 208170 597704 208226
rect 597760 208170 597828 208226
rect 597884 208170 597980 208226
rect -1916 208102 597980 208170
rect -1916 208046 -1820 208102
rect -1764 208046 -1696 208102
rect -1640 208046 -1572 208102
rect -1516 208046 -1448 208102
rect -1392 208046 6970 208102
rect 7026 208046 7094 208102
rect 7150 208046 7218 208102
rect 7274 208046 7342 208102
rect 7398 208046 204970 208102
rect 205026 208046 205094 208102
rect 205150 208046 205218 208102
rect 205274 208046 205342 208102
rect 205398 208046 384970 208102
rect 385026 208046 385094 208102
rect 385150 208046 385218 208102
rect 385274 208046 385342 208102
rect 385398 208046 402970 208102
rect 403026 208046 403094 208102
rect 403150 208046 403218 208102
rect 403274 208046 403342 208102
rect 403398 208046 582970 208102
rect 583026 208046 583094 208102
rect 583150 208046 583218 208102
rect 583274 208046 583342 208102
rect 583398 208046 597456 208102
rect 597512 208046 597580 208102
rect 597636 208046 597704 208102
rect 597760 208046 597828 208102
rect 597884 208046 597980 208102
rect -1916 207978 597980 208046
rect -1916 207922 -1820 207978
rect -1764 207922 -1696 207978
rect -1640 207922 -1572 207978
rect -1516 207922 -1448 207978
rect -1392 207922 6970 207978
rect 7026 207922 7094 207978
rect 7150 207922 7218 207978
rect 7274 207922 7342 207978
rect 7398 207922 204970 207978
rect 205026 207922 205094 207978
rect 205150 207922 205218 207978
rect 205274 207922 205342 207978
rect 205398 207922 384970 207978
rect 385026 207922 385094 207978
rect 385150 207922 385218 207978
rect 385274 207922 385342 207978
rect 385398 207922 402970 207978
rect 403026 207922 403094 207978
rect 403150 207922 403218 207978
rect 403274 207922 403342 207978
rect 403398 207922 582970 207978
rect 583026 207922 583094 207978
rect 583150 207922 583218 207978
rect 583274 207922 583342 207978
rect 583398 207922 597456 207978
rect 597512 207922 597580 207978
rect 597636 207922 597704 207978
rect 597760 207922 597828 207978
rect 597884 207922 597980 207978
rect -1916 207826 597980 207922
rect -1916 202350 597980 202446
rect -1916 202294 -860 202350
rect -804 202294 -736 202350
rect -680 202294 -612 202350
rect -556 202294 -488 202350
rect -432 202294 3250 202350
rect 3306 202294 3374 202350
rect 3430 202294 3498 202350
rect 3554 202294 3622 202350
rect 3678 202294 201250 202350
rect 201306 202294 201374 202350
rect 201430 202294 201498 202350
rect 201554 202294 201622 202350
rect 201678 202294 381250 202350
rect 381306 202294 381374 202350
rect 381430 202294 381498 202350
rect 381554 202294 381622 202350
rect 381678 202294 399250 202350
rect 399306 202294 399374 202350
rect 399430 202294 399498 202350
rect 399554 202294 399622 202350
rect 399678 202294 579250 202350
rect 579306 202294 579374 202350
rect 579430 202294 579498 202350
rect 579554 202294 579622 202350
rect 579678 202294 596496 202350
rect 596552 202294 596620 202350
rect 596676 202294 596744 202350
rect 596800 202294 596868 202350
rect 596924 202294 597980 202350
rect -1916 202226 597980 202294
rect -1916 202170 -860 202226
rect -804 202170 -736 202226
rect -680 202170 -612 202226
rect -556 202170 -488 202226
rect -432 202170 3250 202226
rect 3306 202170 3374 202226
rect 3430 202170 3498 202226
rect 3554 202170 3622 202226
rect 3678 202170 201250 202226
rect 201306 202170 201374 202226
rect 201430 202170 201498 202226
rect 201554 202170 201622 202226
rect 201678 202170 381250 202226
rect 381306 202170 381374 202226
rect 381430 202170 381498 202226
rect 381554 202170 381622 202226
rect 381678 202170 399250 202226
rect 399306 202170 399374 202226
rect 399430 202170 399498 202226
rect 399554 202170 399622 202226
rect 399678 202170 579250 202226
rect 579306 202170 579374 202226
rect 579430 202170 579498 202226
rect 579554 202170 579622 202226
rect 579678 202170 596496 202226
rect 596552 202170 596620 202226
rect 596676 202170 596744 202226
rect 596800 202170 596868 202226
rect 596924 202170 597980 202226
rect -1916 202102 597980 202170
rect -1916 202046 -860 202102
rect -804 202046 -736 202102
rect -680 202046 -612 202102
rect -556 202046 -488 202102
rect -432 202046 3250 202102
rect 3306 202046 3374 202102
rect 3430 202046 3498 202102
rect 3554 202046 3622 202102
rect 3678 202046 201250 202102
rect 201306 202046 201374 202102
rect 201430 202046 201498 202102
rect 201554 202046 201622 202102
rect 201678 202046 381250 202102
rect 381306 202046 381374 202102
rect 381430 202046 381498 202102
rect 381554 202046 381622 202102
rect 381678 202046 399250 202102
rect 399306 202046 399374 202102
rect 399430 202046 399498 202102
rect 399554 202046 399622 202102
rect 399678 202046 579250 202102
rect 579306 202046 579374 202102
rect 579430 202046 579498 202102
rect 579554 202046 579622 202102
rect 579678 202046 596496 202102
rect 596552 202046 596620 202102
rect 596676 202046 596744 202102
rect 596800 202046 596868 202102
rect 596924 202046 597980 202102
rect -1916 201978 597980 202046
rect -1916 201922 -860 201978
rect -804 201922 -736 201978
rect -680 201922 -612 201978
rect -556 201922 -488 201978
rect -432 201922 3250 201978
rect 3306 201922 3374 201978
rect 3430 201922 3498 201978
rect 3554 201922 3622 201978
rect 3678 201922 201250 201978
rect 201306 201922 201374 201978
rect 201430 201922 201498 201978
rect 201554 201922 201622 201978
rect 201678 201922 381250 201978
rect 381306 201922 381374 201978
rect 381430 201922 381498 201978
rect 381554 201922 381622 201978
rect 381678 201922 399250 201978
rect 399306 201922 399374 201978
rect 399430 201922 399498 201978
rect 399554 201922 399622 201978
rect 399678 201922 579250 201978
rect 579306 201922 579374 201978
rect 579430 201922 579498 201978
rect 579554 201922 579622 201978
rect 579678 201922 596496 201978
rect 596552 201922 596620 201978
rect 596676 201922 596744 201978
rect 596800 201922 596868 201978
rect 596924 201922 597980 201978
rect -1916 201826 597980 201922
rect -1916 190350 597980 190446
rect -1916 190294 -1820 190350
rect -1764 190294 -1696 190350
rect -1640 190294 -1572 190350
rect -1516 190294 -1448 190350
rect -1392 190294 6970 190350
rect 7026 190294 7094 190350
rect 7150 190294 7218 190350
rect 7274 190294 7342 190350
rect 7398 190294 204970 190350
rect 205026 190294 205094 190350
rect 205150 190294 205218 190350
rect 205274 190294 205342 190350
rect 205398 190294 384970 190350
rect 385026 190294 385094 190350
rect 385150 190294 385218 190350
rect 385274 190294 385342 190350
rect 385398 190294 402970 190350
rect 403026 190294 403094 190350
rect 403150 190294 403218 190350
rect 403274 190294 403342 190350
rect 403398 190294 582970 190350
rect 583026 190294 583094 190350
rect 583150 190294 583218 190350
rect 583274 190294 583342 190350
rect 583398 190294 597456 190350
rect 597512 190294 597580 190350
rect 597636 190294 597704 190350
rect 597760 190294 597828 190350
rect 597884 190294 597980 190350
rect -1916 190226 597980 190294
rect -1916 190170 -1820 190226
rect -1764 190170 -1696 190226
rect -1640 190170 -1572 190226
rect -1516 190170 -1448 190226
rect -1392 190170 6970 190226
rect 7026 190170 7094 190226
rect 7150 190170 7218 190226
rect 7274 190170 7342 190226
rect 7398 190170 204970 190226
rect 205026 190170 205094 190226
rect 205150 190170 205218 190226
rect 205274 190170 205342 190226
rect 205398 190170 384970 190226
rect 385026 190170 385094 190226
rect 385150 190170 385218 190226
rect 385274 190170 385342 190226
rect 385398 190170 402970 190226
rect 403026 190170 403094 190226
rect 403150 190170 403218 190226
rect 403274 190170 403342 190226
rect 403398 190170 582970 190226
rect 583026 190170 583094 190226
rect 583150 190170 583218 190226
rect 583274 190170 583342 190226
rect 583398 190170 597456 190226
rect 597512 190170 597580 190226
rect 597636 190170 597704 190226
rect 597760 190170 597828 190226
rect 597884 190170 597980 190226
rect -1916 190102 597980 190170
rect -1916 190046 -1820 190102
rect -1764 190046 -1696 190102
rect -1640 190046 -1572 190102
rect -1516 190046 -1448 190102
rect -1392 190046 6970 190102
rect 7026 190046 7094 190102
rect 7150 190046 7218 190102
rect 7274 190046 7342 190102
rect 7398 190046 204970 190102
rect 205026 190046 205094 190102
rect 205150 190046 205218 190102
rect 205274 190046 205342 190102
rect 205398 190046 384970 190102
rect 385026 190046 385094 190102
rect 385150 190046 385218 190102
rect 385274 190046 385342 190102
rect 385398 190046 402970 190102
rect 403026 190046 403094 190102
rect 403150 190046 403218 190102
rect 403274 190046 403342 190102
rect 403398 190046 582970 190102
rect 583026 190046 583094 190102
rect 583150 190046 583218 190102
rect 583274 190046 583342 190102
rect 583398 190046 597456 190102
rect 597512 190046 597580 190102
rect 597636 190046 597704 190102
rect 597760 190046 597828 190102
rect 597884 190046 597980 190102
rect -1916 189978 597980 190046
rect -1916 189922 -1820 189978
rect -1764 189922 -1696 189978
rect -1640 189922 -1572 189978
rect -1516 189922 -1448 189978
rect -1392 189922 6970 189978
rect 7026 189922 7094 189978
rect 7150 189922 7218 189978
rect 7274 189922 7342 189978
rect 7398 189922 204970 189978
rect 205026 189922 205094 189978
rect 205150 189922 205218 189978
rect 205274 189922 205342 189978
rect 205398 189922 384970 189978
rect 385026 189922 385094 189978
rect 385150 189922 385218 189978
rect 385274 189922 385342 189978
rect 385398 189922 402970 189978
rect 403026 189922 403094 189978
rect 403150 189922 403218 189978
rect 403274 189922 403342 189978
rect 403398 189922 582970 189978
rect 583026 189922 583094 189978
rect 583150 189922 583218 189978
rect 583274 189922 583342 189978
rect 583398 189922 597456 189978
rect 597512 189922 597580 189978
rect 597636 189922 597704 189978
rect 597760 189922 597828 189978
rect 597884 189922 597980 189978
rect -1916 189826 597980 189922
rect -1916 184350 597980 184446
rect -1916 184294 -860 184350
rect -804 184294 -736 184350
rect -680 184294 -612 184350
rect -556 184294 -488 184350
rect -432 184294 3250 184350
rect 3306 184294 3374 184350
rect 3430 184294 3498 184350
rect 3554 184294 3622 184350
rect 3678 184294 201250 184350
rect 201306 184294 201374 184350
rect 201430 184294 201498 184350
rect 201554 184294 201622 184350
rect 201678 184294 381250 184350
rect 381306 184294 381374 184350
rect 381430 184294 381498 184350
rect 381554 184294 381622 184350
rect 381678 184294 399250 184350
rect 399306 184294 399374 184350
rect 399430 184294 399498 184350
rect 399554 184294 399622 184350
rect 399678 184294 579250 184350
rect 579306 184294 579374 184350
rect 579430 184294 579498 184350
rect 579554 184294 579622 184350
rect 579678 184294 596496 184350
rect 596552 184294 596620 184350
rect 596676 184294 596744 184350
rect 596800 184294 596868 184350
rect 596924 184294 597980 184350
rect -1916 184226 597980 184294
rect -1916 184170 -860 184226
rect -804 184170 -736 184226
rect -680 184170 -612 184226
rect -556 184170 -488 184226
rect -432 184170 3250 184226
rect 3306 184170 3374 184226
rect 3430 184170 3498 184226
rect 3554 184170 3622 184226
rect 3678 184170 201250 184226
rect 201306 184170 201374 184226
rect 201430 184170 201498 184226
rect 201554 184170 201622 184226
rect 201678 184170 381250 184226
rect 381306 184170 381374 184226
rect 381430 184170 381498 184226
rect 381554 184170 381622 184226
rect 381678 184170 399250 184226
rect 399306 184170 399374 184226
rect 399430 184170 399498 184226
rect 399554 184170 399622 184226
rect 399678 184170 579250 184226
rect 579306 184170 579374 184226
rect 579430 184170 579498 184226
rect 579554 184170 579622 184226
rect 579678 184170 596496 184226
rect 596552 184170 596620 184226
rect 596676 184170 596744 184226
rect 596800 184170 596868 184226
rect 596924 184170 597980 184226
rect -1916 184102 597980 184170
rect -1916 184046 -860 184102
rect -804 184046 -736 184102
rect -680 184046 -612 184102
rect -556 184046 -488 184102
rect -432 184046 3250 184102
rect 3306 184046 3374 184102
rect 3430 184046 3498 184102
rect 3554 184046 3622 184102
rect 3678 184046 201250 184102
rect 201306 184046 201374 184102
rect 201430 184046 201498 184102
rect 201554 184046 201622 184102
rect 201678 184046 381250 184102
rect 381306 184046 381374 184102
rect 381430 184046 381498 184102
rect 381554 184046 381622 184102
rect 381678 184046 399250 184102
rect 399306 184046 399374 184102
rect 399430 184046 399498 184102
rect 399554 184046 399622 184102
rect 399678 184046 579250 184102
rect 579306 184046 579374 184102
rect 579430 184046 579498 184102
rect 579554 184046 579622 184102
rect 579678 184046 596496 184102
rect 596552 184046 596620 184102
rect 596676 184046 596744 184102
rect 596800 184046 596868 184102
rect 596924 184046 597980 184102
rect -1916 183978 597980 184046
rect -1916 183922 -860 183978
rect -804 183922 -736 183978
rect -680 183922 -612 183978
rect -556 183922 -488 183978
rect -432 183922 3250 183978
rect 3306 183922 3374 183978
rect 3430 183922 3498 183978
rect 3554 183922 3622 183978
rect 3678 183922 201250 183978
rect 201306 183922 201374 183978
rect 201430 183922 201498 183978
rect 201554 183922 201622 183978
rect 201678 183922 381250 183978
rect 381306 183922 381374 183978
rect 381430 183922 381498 183978
rect 381554 183922 381622 183978
rect 381678 183922 399250 183978
rect 399306 183922 399374 183978
rect 399430 183922 399498 183978
rect 399554 183922 399622 183978
rect 399678 183922 579250 183978
rect 579306 183922 579374 183978
rect 579430 183922 579498 183978
rect 579554 183922 579622 183978
rect 579678 183922 596496 183978
rect 596552 183922 596620 183978
rect 596676 183922 596744 183978
rect 596800 183922 596868 183978
rect 596924 183922 597980 183978
rect -1916 183826 597980 183922
rect -1916 172350 597980 172446
rect -1916 172294 -1820 172350
rect -1764 172294 -1696 172350
rect -1640 172294 -1572 172350
rect -1516 172294 -1448 172350
rect -1392 172294 6970 172350
rect 7026 172294 7094 172350
rect 7150 172294 7218 172350
rect 7274 172294 7342 172350
rect 7398 172294 204970 172350
rect 205026 172294 205094 172350
rect 205150 172294 205218 172350
rect 205274 172294 205342 172350
rect 205398 172294 384970 172350
rect 385026 172294 385094 172350
rect 385150 172294 385218 172350
rect 385274 172294 385342 172350
rect 385398 172294 402970 172350
rect 403026 172294 403094 172350
rect 403150 172294 403218 172350
rect 403274 172294 403342 172350
rect 403398 172294 582970 172350
rect 583026 172294 583094 172350
rect 583150 172294 583218 172350
rect 583274 172294 583342 172350
rect 583398 172294 597456 172350
rect 597512 172294 597580 172350
rect 597636 172294 597704 172350
rect 597760 172294 597828 172350
rect 597884 172294 597980 172350
rect -1916 172226 597980 172294
rect -1916 172170 -1820 172226
rect -1764 172170 -1696 172226
rect -1640 172170 -1572 172226
rect -1516 172170 -1448 172226
rect -1392 172170 6970 172226
rect 7026 172170 7094 172226
rect 7150 172170 7218 172226
rect 7274 172170 7342 172226
rect 7398 172170 204970 172226
rect 205026 172170 205094 172226
rect 205150 172170 205218 172226
rect 205274 172170 205342 172226
rect 205398 172170 384970 172226
rect 385026 172170 385094 172226
rect 385150 172170 385218 172226
rect 385274 172170 385342 172226
rect 385398 172170 402970 172226
rect 403026 172170 403094 172226
rect 403150 172170 403218 172226
rect 403274 172170 403342 172226
rect 403398 172170 582970 172226
rect 583026 172170 583094 172226
rect 583150 172170 583218 172226
rect 583274 172170 583342 172226
rect 583398 172170 597456 172226
rect 597512 172170 597580 172226
rect 597636 172170 597704 172226
rect 597760 172170 597828 172226
rect 597884 172170 597980 172226
rect -1916 172102 597980 172170
rect -1916 172046 -1820 172102
rect -1764 172046 -1696 172102
rect -1640 172046 -1572 172102
rect -1516 172046 -1448 172102
rect -1392 172046 6970 172102
rect 7026 172046 7094 172102
rect 7150 172046 7218 172102
rect 7274 172046 7342 172102
rect 7398 172046 204970 172102
rect 205026 172046 205094 172102
rect 205150 172046 205218 172102
rect 205274 172046 205342 172102
rect 205398 172046 384970 172102
rect 385026 172046 385094 172102
rect 385150 172046 385218 172102
rect 385274 172046 385342 172102
rect 385398 172046 402970 172102
rect 403026 172046 403094 172102
rect 403150 172046 403218 172102
rect 403274 172046 403342 172102
rect 403398 172046 582970 172102
rect 583026 172046 583094 172102
rect 583150 172046 583218 172102
rect 583274 172046 583342 172102
rect 583398 172046 597456 172102
rect 597512 172046 597580 172102
rect 597636 172046 597704 172102
rect 597760 172046 597828 172102
rect 597884 172046 597980 172102
rect -1916 171978 597980 172046
rect -1916 171922 -1820 171978
rect -1764 171922 -1696 171978
rect -1640 171922 -1572 171978
rect -1516 171922 -1448 171978
rect -1392 171922 6970 171978
rect 7026 171922 7094 171978
rect 7150 171922 7218 171978
rect 7274 171922 7342 171978
rect 7398 171922 204970 171978
rect 205026 171922 205094 171978
rect 205150 171922 205218 171978
rect 205274 171922 205342 171978
rect 205398 171922 384970 171978
rect 385026 171922 385094 171978
rect 385150 171922 385218 171978
rect 385274 171922 385342 171978
rect 385398 171922 402970 171978
rect 403026 171922 403094 171978
rect 403150 171922 403218 171978
rect 403274 171922 403342 171978
rect 403398 171922 582970 171978
rect 583026 171922 583094 171978
rect 583150 171922 583218 171978
rect 583274 171922 583342 171978
rect 583398 171922 597456 171978
rect 597512 171922 597580 171978
rect 597636 171922 597704 171978
rect 597760 171922 597828 171978
rect 597884 171922 597980 171978
rect -1916 171826 597980 171922
rect -1916 166350 597980 166446
rect -1916 166294 -860 166350
rect -804 166294 -736 166350
rect -680 166294 -612 166350
rect -556 166294 -488 166350
rect -432 166294 3250 166350
rect 3306 166294 3374 166350
rect 3430 166294 3498 166350
rect 3554 166294 3622 166350
rect 3678 166294 201250 166350
rect 201306 166294 201374 166350
rect 201430 166294 201498 166350
rect 201554 166294 201622 166350
rect 201678 166294 381250 166350
rect 381306 166294 381374 166350
rect 381430 166294 381498 166350
rect 381554 166294 381622 166350
rect 381678 166294 399250 166350
rect 399306 166294 399374 166350
rect 399430 166294 399498 166350
rect 399554 166294 399622 166350
rect 399678 166294 579250 166350
rect 579306 166294 579374 166350
rect 579430 166294 579498 166350
rect 579554 166294 579622 166350
rect 579678 166294 596496 166350
rect 596552 166294 596620 166350
rect 596676 166294 596744 166350
rect 596800 166294 596868 166350
rect 596924 166294 597980 166350
rect -1916 166226 597980 166294
rect -1916 166170 -860 166226
rect -804 166170 -736 166226
rect -680 166170 -612 166226
rect -556 166170 -488 166226
rect -432 166170 3250 166226
rect 3306 166170 3374 166226
rect 3430 166170 3498 166226
rect 3554 166170 3622 166226
rect 3678 166170 201250 166226
rect 201306 166170 201374 166226
rect 201430 166170 201498 166226
rect 201554 166170 201622 166226
rect 201678 166170 381250 166226
rect 381306 166170 381374 166226
rect 381430 166170 381498 166226
rect 381554 166170 381622 166226
rect 381678 166170 399250 166226
rect 399306 166170 399374 166226
rect 399430 166170 399498 166226
rect 399554 166170 399622 166226
rect 399678 166170 579250 166226
rect 579306 166170 579374 166226
rect 579430 166170 579498 166226
rect 579554 166170 579622 166226
rect 579678 166170 596496 166226
rect 596552 166170 596620 166226
rect 596676 166170 596744 166226
rect 596800 166170 596868 166226
rect 596924 166170 597980 166226
rect -1916 166102 597980 166170
rect -1916 166046 -860 166102
rect -804 166046 -736 166102
rect -680 166046 -612 166102
rect -556 166046 -488 166102
rect -432 166046 3250 166102
rect 3306 166046 3374 166102
rect 3430 166046 3498 166102
rect 3554 166046 3622 166102
rect 3678 166046 201250 166102
rect 201306 166046 201374 166102
rect 201430 166046 201498 166102
rect 201554 166046 201622 166102
rect 201678 166046 381250 166102
rect 381306 166046 381374 166102
rect 381430 166046 381498 166102
rect 381554 166046 381622 166102
rect 381678 166046 399250 166102
rect 399306 166046 399374 166102
rect 399430 166046 399498 166102
rect 399554 166046 399622 166102
rect 399678 166046 579250 166102
rect 579306 166046 579374 166102
rect 579430 166046 579498 166102
rect 579554 166046 579622 166102
rect 579678 166046 596496 166102
rect 596552 166046 596620 166102
rect 596676 166046 596744 166102
rect 596800 166046 596868 166102
rect 596924 166046 597980 166102
rect -1916 165978 597980 166046
rect -1916 165922 -860 165978
rect -804 165922 -736 165978
rect -680 165922 -612 165978
rect -556 165922 -488 165978
rect -432 165922 3250 165978
rect 3306 165922 3374 165978
rect 3430 165922 3498 165978
rect 3554 165922 3622 165978
rect 3678 165922 201250 165978
rect 201306 165922 201374 165978
rect 201430 165922 201498 165978
rect 201554 165922 201622 165978
rect 201678 165922 381250 165978
rect 381306 165922 381374 165978
rect 381430 165922 381498 165978
rect 381554 165922 381622 165978
rect 381678 165922 399250 165978
rect 399306 165922 399374 165978
rect 399430 165922 399498 165978
rect 399554 165922 399622 165978
rect 399678 165922 579250 165978
rect 579306 165922 579374 165978
rect 579430 165922 579498 165978
rect 579554 165922 579622 165978
rect 579678 165922 596496 165978
rect 596552 165922 596620 165978
rect 596676 165922 596744 165978
rect 596800 165922 596868 165978
rect 596924 165922 597980 165978
rect -1916 165826 597980 165922
rect -1916 154350 597980 154446
rect -1916 154294 -1820 154350
rect -1764 154294 -1696 154350
rect -1640 154294 -1572 154350
rect -1516 154294 -1448 154350
rect -1392 154294 6970 154350
rect 7026 154294 7094 154350
rect 7150 154294 7218 154350
rect 7274 154294 7342 154350
rect 7398 154294 24970 154350
rect 25026 154294 25094 154350
rect 25150 154294 25218 154350
rect 25274 154294 25342 154350
rect 25398 154294 42970 154350
rect 43026 154294 43094 154350
rect 43150 154294 43218 154350
rect 43274 154294 43342 154350
rect 43398 154294 60970 154350
rect 61026 154294 61094 154350
rect 61150 154294 61218 154350
rect 61274 154294 61342 154350
rect 61398 154294 78970 154350
rect 79026 154294 79094 154350
rect 79150 154294 79218 154350
rect 79274 154294 79342 154350
rect 79398 154294 96970 154350
rect 97026 154294 97094 154350
rect 97150 154294 97218 154350
rect 97274 154294 97342 154350
rect 97398 154294 114970 154350
rect 115026 154294 115094 154350
rect 115150 154294 115218 154350
rect 115274 154294 115342 154350
rect 115398 154294 132970 154350
rect 133026 154294 133094 154350
rect 133150 154294 133218 154350
rect 133274 154294 133342 154350
rect 133398 154294 150970 154350
rect 151026 154294 151094 154350
rect 151150 154294 151218 154350
rect 151274 154294 151342 154350
rect 151398 154294 168970 154350
rect 169026 154294 169094 154350
rect 169150 154294 169218 154350
rect 169274 154294 169342 154350
rect 169398 154294 186970 154350
rect 187026 154294 187094 154350
rect 187150 154294 187218 154350
rect 187274 154294 187342 154350
rect 187398 154294 204970 154350
rect 205026 154294 205094 154350
rect 205150 154294 205218 154350
rect 205274 154294 205342 154350
rect 205398 154294 222970 154350
rect 223026 154294 223094 154350
rect 223150 154294 223218 154350
rect 223274 154294 223342 154350
rect 223398 154294 240970 154350
rect 241026 154294 241094 154350
rect 241150 154294 241218 154350
rect 241274 154294 241342 154350
rect 241398 154294 258970 154350
rect 259026 154294 259094 154350
rect 259150 154294 259218 154350
rect 259274 154294 259342 154350
rect 259398 154294 276970 154350
rect 277026 154294 277094 154350
rect 277150 154294 277218 154350
rect 277274 154294 277342 154350
rect 277398 154294 294970 154350
rect 295026 154294 295094 154350
rect 295150 154294 295218 154350
rect 295274 154294 295342 154350
rect 295398 154294 312970 154350
rect 313026 154294 313094 154350
rect 313150 154294 313218 154350
rect 313274 154294 313342 154350
rect 313398 154294 330970 154350
rect 331026 154294 331094 154350
rect 331150 154294 331218 154350
rect 331274 154294 331342 154350
rect 331398 154294 348970 154350
rect 349026 154294 349094 154350
rect 349150 154294 349218 154350
rect 349274 154294 349342 154350
rect 349398 154294 366970 154350
rect 367026 154294 367094 154350
rect 367150 154294 367218 154350
rect 367274 154294 367342 154350
rect 367398 154294 384970 154350
rect 385026 154294 385094 154350
rect 385150 154294 385218 154350
rect 385274 154294 385342 154350
rect 385398 154294 402970 154350
rect 403026 154294 403094 154350
rect 403150 154294 403218 154350
rect 403274 154294 403342 154350
rect 403398 154294 420970 154350
rect 421026 154294 421094 154350
rect 421150 154294 421218 154350
rect 421274 154294 421342 154350
rect 421398 154294 438970 154350
rect 439026 154294 439094 154350
rect 439150 154294 439218 154350
rect 439274 154294 439342 154350
rect 439398 154294 456970 154350
rect 457026 154294 457094 154350
rect 457150 154294 457218 154350
rect 457274 154294 457342 154350
rect 457398 154294 474970 154350
rect 475026 154294 475094 154350
rect 475150 154294 475218 154350
rect 475274 154294 475342 154350
rect 475398 154294 492970 154350
rect 493026 154294 493094 154350
rect 493150 154294 493218 154350
rect 493274 154294 493342 154350
rect 493398 154294 510970 154350
rect 511026 154294 511094 154350
rect 511150 154294 511218 154350
rect 511274 154294 511342 154350
rect 511398 154294 528970 154350
rect 529026 154294 529094 154350
rect 529150 154294 529218 154350
rect 529274 154294 529342 154350
rect 529398 154294 546970 154350
rect 547026 154294 547094 154350
rect 547150 154294 547218 154350
rect 547274 154294 547342 154350
rect 547398 154294 564970 154350
rect 565026 154294 565094 154350
rect 565150 154294 565218 154350
rect 565274 154294 565342 154350
rect 565398 154294 582970 154350
rect 583026 154294 583094 154350
rect 583150 154294 583218 154350
rect 583274 154294 583342 154350
rect 583398 154294 597456 154350
rect 597512 154294 597580 154350
rect 597636 154294 597704 154350
rect 597760 154294 597828 154350
rect 597884 154294 597980 154350
rect -1916 154226 597980 154294
rect -1916 154170 -1820 154226
rect -1764 154170 -1696 154226
rect -1640 154170 -1572 154226
rect -1516 154170 -1448 154226
rect -1392 154170 6970 154226
rect 7026 154170 7094 154226
rect 7150 154170 7218 154226
rect 7274 154170 7342 154226
rect 7398 154170 24970 154226
rect 25026 154170 25094 154226
rect 25150 154170 25218 154226
rect 25274 154170 25342 154226
rect 25398 154170 42970 154226
rect 43026 154170 43094 154226
rect 43150 154170 43218 154226
rect 43274 154170 43342 154226
rect 43398 154170 60970 154226
rect 61026 154170 61094 154226
rect 61150 154170 61218 154226
rect 61274 154170 61342 154226
rect 61398 154170 78970 154226
rect 79026 154170 79094 154226
rect 79150 154170 79218 154226
rect 79274 154170 79342 154226
rect 79398 154170 96970 154226
rect 97026 154170 97094 154226
rect 97150 154170 97218 154226
rect 97274 154170 97342 154226
rect 97398 154170 114970 154226
rect 115026 154170 115094 154226
rect 115150 154170 115218 154226
rect 115274 154170 115342 154226
rect 115398 154170 132970 154226
rect 133026 154170 133094 154226
rect 133150 154170 133218 154226
rect 133274 154170 133342 154226
rect 133398 154170 150970 154226
rect 151026 154170 151094 154226
rect 151150 154170 151218 154226
rect 151274 154170 151342 154226
rect 151398 154170 168970 154226
rect 169026 154170 169094 154226
rect 169150 154170 169218 154226
rect 169274 154170 169342 154226
rect 169398 154170 186970 154226
rect 187026 154170 187094 154226
rect 187150 154170 187218 154226
rect 187274 154170 187342 154226
rect 187398 154170 204970 154226
rect 205026 154170 205094 154226
rect 205150 154170 205218 154226
rect 205274 154170 205342 154226
rect 205398 154170 222970 154226
rect 223026 154170 223094 154226
rect 223150 154170 223218 154226
rect 223274 154170 223342 154226
rect 223398 154170 240970 154226
rect 241026 154170 241094 154226
rect 241150 154170 241218 154226
rect 241274 154170 241342 154226
rect 241398 154170 258970 154226
rect 259026 154170 259094 154226
rect 259150 154170 259218 154226
rect 259274 154170 259342 154226
rect 259398 154170 276970 154226
rect 277026 154170 277094 154226
rect 277150 154170 277218 154226
rect 277274 154170 277342 154226
rect 277398 154170 294970 154226
rect 295026 154170 295094 154226
rect 295150 154170 295218 154226
rect 295274 154170 295342 154226
rect 295398 154170 312970 154226
rect 313026 154170 313094 154226
rect 313150 154170 313218 154226
rect 313274 154170 313342 154226
rect 313398 154170 330970 154226
rect 331026 154170 331094 154226
rect 331150 154170 331218 154226
rect 331274 154170 331342 154226
rect 331398 154170 348970 154226
rect 349026 154170 349094 154226
rect 349150 154170 349218 154226
rect 349274 154170 349342 154226
rect 349398 154170 366970 154226
rect 367026 154170 367094 154226
rect 367150 154170 367218 154226
rect 367274 154170 367342 154226
rect 367398 154170 384970 154226
rect 385026 154170 385094 154226
rect 385150 154170 385218 154226
rect 385274 154170 385342 154226
rect 385398 154170 402970 154226
rect 403026 154170 403094 154226
rect 403150 154170 403218 154226
rect 403274 154170 403342 154226
rect 403398 154170 420970 154226
rect 421026 154170 421094 154226
rect 421150 154170 421218 154226
rect 421274 154170 421342 154226
rect 421398 154170 438970 154226
rect 439026 154170 439094 154226
rect 439150 154170 439218 154226
rect 439274 154170 439342 154226
rect 439398 154170 456970 154226
rect 457026 154170 457094 154226
rect 457150 154170 457218 154226
rect 457274 154170 457342 154226
rect 457398 154170 474970 154226
rect 475026 154170 475094 154226
rect 475150 154170 475218 154226
rect 475274 154170 475342 154226
rect 475398 154170 492970 154226
rect 493026 154170 493094 154226
rect 493150 154170 493218 154226
rect 493274 154170 493342 154226
rect 493398 154170 510970 154226
rect 511026 154170 511094 154226
rect 511150 154170 511218 154226
rect 511274 154170 511342 154226
rect 511398 154170 528970 154226
rect 529026 154170 529094 154226
rect 529150 154170 529218 154226
rect 529274 154170 529342 154226
rect 529398 154170 546970 154226
rect 547026 154170 547094 154226
rect 547150 154170 547218 154226
rect 547274 154170 547342 154226
rect 547398 154170 564970 154226
rect 565026 154170 565094 154226
rect 565150 154170 565218 154226
rect 565274 154170 565342 154226
rect 565398 154170 582970 154226
rect 583026 154170 583094 154226
rect 583150 154170 583218 154226
rect 583274 154170 583342 154226
rect 583398 154170 597456 154226
rect 597512 154170 597580 154226
rect 597636 154170 597704 154226
rect 597760 154170 597828 154226
rect 597884 154170 597980 154226
rect -1916 154102 597980 154170
rect -1916 154046 -1820 154102
rect -1764 154046 -1696 154102
rect -1640 154046 -1572 154102
rect -1516 154046 -1448 154102
rect -1392 154046 6970 154102
rect 7026 154046 7094 154102
rect 7150 154046 7218 154102
rect 7274 154046 7342 154102
rect 7398 154046 24970 154102
rect 25026 154046 25094 154102
rect 25150 154046 25218 154102
rect 25274 154046 25342 154102
rect 25398 154046 42970 154102
rect 43026 154046 43094 154102
rect 43150 154046 43218 154102
rect 43274 154046 43342 154102
rect 43398 154046 60970 154102
rect 61026 154046 61094 154102
rect 61150 154046 61218 154102
rect 61274 154046 61342 154102
rect 61398 154046 78970 154102
rect 79026 154046 79094 154102
rect 79150 154046 79218 154102
rect 79274 154046 79342 154102
rect 79398 154046 96970 154102
rect 97026 154046 97094 154102
rect 97150 154046 97218 154102
rect 97274 154046 97342 154102
rect 97398 154046 114970 154102
rect 115026 154046 115094 154102
rect 115150 154046 115218 154102
rect 115274 154046 115342 154102
rect 115398 154046 132970 154102
rect 133026 154046 133094 154102
rect 133150 154046 133218 154102
rect 133274 154046 133342 154102
rect 133398 154046 150970 154102
rect 151026 154046 151094 154102
rect 151150 154046 151218 154102
rect 151274 154046 151342 154102
rect 151398 154046 168970 154102
rect 169026 154046 169094 154102
rect 169150 154046 169218 154102
rect 169274 154046 169342 154102
rect 169398 154046 186970 154102
rect 187026 154046 187094 154102
rect 187150 154046 187218 154102
rect 187274 154046 187342 154102
rect 187398 154046 204970 154102
rect 205026 154046 205094 154102
rect 205150 154046 205218 154102
rect 205274 154046 205342 154102
rect 205398 154046 222970 154102
rect 223026 154046 223094 154102
rect 223150 154046 223218 154102
rect 223274 154046 223342 154102
rect 223398 154046 240970 154102
rect 241026 154046 241094 154102
rect 241150 154046 241218 154102
rect 241274 154046 241342 154102
rect 241398 154046 258970 154102
rect 259026 154046 259094 154102
rect 259150 154046 259218 154102
rect 259274 154046 259342 154102
rect 259398 154046 276970 154102
rect 277026 154046 277094 154102
rect 277150 154046 277218 154102
rect 277274 154046 277342 154102
rect 277398 154046 294970 154102
rect 295026 154046 295094 154102
rect 295150 154046 295218 154102
rect 295274 154046 295342 154102
rect 295398 154046 312970 154102
rect 313026 154046 313094 154102
rect 313150 154046 313218 154102
rect 313274 154046 313342 154102
rect 313398 154046 330970 154102
rect 331026 154046 331094 154102
rect 331150 154046 331218 154102
rect 331274 154046 331342 154102
rect 331398 154046 348970 154102
rect 349026 154046 349094 154102
rect 349150 154046 349218 154102
rect 349274 154046 349342 154102
rect 349398 154046 366970 154102
rect 367026 154046 367094 154102
rect 367150 154046 367218 154102
rect 367274 154046 367342 154102
rect 367398 154046 384970 154102
rect 385026 154046 385094 154102
rect 385150 154046 385218 154102
rect 385274 154046 385342 154102
rect 385398 154046 402970 154102
rect 403026 154046 403094 154102
rect 403150 154046 403218 154102
rect 403274 154046 403342 154102
rect 403398 154046 420970 154102
rect 421026 154046 421094 154102
rect 421150 154046 421218 154102
rect 421274 154046 421342 154102
rect 421398 154046 438970 154102
rect 439026 154046 439094 154102
rect 439150 154046 439218 154102
rect 439274 154046 439342 154102
rect 439398 154046 456970 154102
rect 457026 154046 457094 154102
rect 457150 154046 457218 154102
rect 457274 154046 457342 154102
rect 457398 154046 474970 154102
rect 475026 154046 475094 154102
rect 475150 154046 475218 154102
rect 475274 154046 475342 154102
rect 475398 154046 492970 154102
rect 493026 154046 493094 154102
rect 493150 154046 493218 154102
rect 493274 154046 493342 154102
rect 493398 154046 510970 154102
rect 511026 154046 511094 154102
rect 511150 154046 511218 154102
rect 511274 154046 511342 154102
rect 511398 154046 528970 154102
rect 529026 154046 529094 154102
rect 529150 154046 529218 154102
rect 529274 154046 529342 154102
rect 529398 154046 546970 154102
rect 547026 154046 547094 154102
rect 547150 154046 547218 154102
rect 547274 154046 547342 154102
rect 547398 154046 564970 154102
rect 565026 154046 565094 154102
rect 565150 154046 565218 154102
rect 565274 154046 565342 154102
rect 565398 154046 582970 154102
rect 583026 154046 583094 154102
rect 583150 154046 583218 154102
rect 583274 154046 583342 154102
rect 583398 154046 597456 154102
rect 597512 154046 597580 154102
rect 597636 154046 597704 154102
rect 597760 154046 597828 154102
rect 597884 154046 597980 154102
rect -1916 153978 597980 154046
rect -1916 153922 -1820 153978
rect -1764 153922 -1696 153978
rect -1640 153922 -1572 153978
rect -1516 153922 -1448 153978
rect -1392 153922 6970 153978
rect 7026 153922 7094 153978
rect 7150 153922 7218 153978
rect 7274 153922 7342 153978
rect 7398 153922 24970 153978
rect 25026 153922 25094 153978
rect 25150 153922 25218 153978
rect 25274 153922 25342 153978
rect 25398 153922 42970 153978
rect 43026 153922 43094 153978
rect 43150 153922 43218 153978
rect 43274 153922 43342 153978
rect 43398 153922 60970 153978
rect 61026 153922 61094 153978
rect 61150 153922 61218 153978
rect 61274 153922 61342 153978
rect 61398 153922 78970 153978
rect 79026 153922 79094 153978
rect 79150 153922 79218 153978
rect 79274 153922 79342 153978
rect 79398 153922 96970 153978
rect 97026 153922 97094 153978
rect 97150 153922 97218 153978
rect 97274 153922 97342 153978
rect 97398 153922 114970 153978
rect 115026 153922 115094 153978
rect 115150 153922 115218 153978
rect 115274 153922 115342 153978
rect 115398 153922 132970 153978
rect 133026 153922 133094 153978
rect 133150 153922 133218 153978
rect 133274 153922 133342 153978
rect 133398 153922 150970 153978
rect 151026 153922 151094 153978
rect 151150 153922 151218 153978
rect 151274 153922 151342 153978
rect 151398 153922 168970 153978
rect 169026 153922 169094 153978
rect 169150 153922 169218 153978
rect 169274 153922 169342 153978
rect 169398 153922 186970 153978
rect 187026 153922 187094 153978
rect 187150 153922 187218 153978
rect 187274 153922 187342 153978
rect 187398 153922 204970 153978
rect 205026 153922 205094 153978
rect 205150 153922 205218 153978
rect 205274 153922 205342 153978
rect 205398 153922 222970 153978
rect 223026 153922 223094 153978
rect 223150 153922 223218 153978
rect 223274 153922 223342 153978
rect 223398 153922 240970 153978
rect 241026 153922 241094 153978
rect 241150 153922 241218 153978
rect 241274 153922 241342 153978
rect 241398 153922 258970 153978
rect 259026 153922 259094 153978
rect 259150 153922 259218 153978
rect 259274 153922 259342 153978
rect 259398 153922 276970 153978
rect 277026 153922 277094 153978
rect 277150 153922 277218 153978
rect 277274 153922 277342 153978
rect 277398 153922 294970 153978
rect 295026 153922 295094 153978
rect 295150 153922 295218 153978
rect 295274 153922 295342 153978
rect 295398 153922 312970 153978
rect 313026 153922 313094 153978
rect 313150 153922 313218 153978
rect 313274 153922 313342 153978
rect 313398 153922 330970 153978
rect 331026 153922 331094 153978
rect 331150 153922 331218 153978
rect 331274 153922 331342 153978
rect 331398 153922 348970 153978
rect 349026 153922 349094 153978
rect 349150 153922 349218 153978
rect 349274 153922 349342 153978
rect 349398 153922 366970 153978
rect 367026 153922 367094 153978
rect 367150 153922 367218 153978
rect 367274 153922 367342 153978
rect 367398 153922 384970 153978
rect 385026 153922 385094 153978
rect 385150 153922 385218 153978
rect 385274 153922 385342 153978
rect 385398 153922 402970 153978
rect 403026 153922 403094 153978
rect 403150 153922 403218 153978
rect 403274 153922 403342 153978
rect 403398 153922 420970 153978
rect 421026 153922 421094 153978
rect 421150 153922 421218 153978
rect 421274 153922 421342 153978
rect 421398 153922 438970 153978
rect 439026 153922 439094 153978
rect 439150 153922 439218 153978
rect 439274 153922 439342 153978
rect 439398 153922 456970 153978
rect 457026 153922 457094 153978
rect 457150 153922 457218 153978
rect 457274 153922 457342 153978
rect 457398 153922 474970 153978
rect 475026 153922 475094 153978
rect 475150 153922 475218 153978
rect 475274 153922 475342 153978
rect 475398 153922 492970 153978
rect 493026 153922 493094 153978
rect 493150 153922 493218 153978
rect 493274 153922 493342 153978
rect 493398 153922 510970 153978
rect 511026 153922 511094 153978
rect 511150 153922 511218 153978
rect 511274 153922 511342 153978
rect 511398 153922 528970 153978
rect 529026 153922 529094 153978
rect 529150 153922 529218 153978
rect 529274 153922 529342 153978
rect 529398 153922 546970 153978
rect 547026 153922 547094 153978
rect 547150 153922 547218 153978
rect 547274 153922 547342 153978
rect 547398 153922 564970 153978
rect 565026 153922 565094 153978
rect 565150 153922 565218 153978
rect 565274 153922 565342 153978
rect 565398 153922 582970 153978
rect 583026 153922 583094 153978
rect 583150 153922 583218 153978
rect 583274 153922 583342 153978
rect 583398 153922 597456 153978
rect 597512 153922 597580 153978
rect 597636 153922 597704 153978
rect 597760 153922 597828 153978
rect 597884 153922 597980 153978
rect -1916 153826 597980 153922
rect -1916 148422 597980 148446
rect -1916 148366 219250 148422
rect 219306 148366 219374 148422
rect 219430 148366 219498 148422
rect 219554 148366 219622 148422
rect 219678 148366 237250 148422
rect 237306 148366 237374 148422
rect 237430 148366 237498 148422
rect 237554 148366 237622 148422
rect 237678 148366 255250 148422
rect 255306 148366 255374 148422
rect 255430 148366 255498 148422
rect 255554 148366 255622 148422
rect 255678 148366 273250 148422
rect 273306 148366 273374 148422
rect 273430 148366 273498 148422
rect 273554 148366 273622 148422
rect 273678 148366 291250 148422
rect 291306 148366 291374 148422
rect 291430 148366 291498 148422
rect 291554 148366 291622 148422
rect 291678 148366 309250 148422
rect 309306 148366 309374 148422
rect 309430 148366 309498 148422
rect 309554 148366 309622 148422
rect 309678 148366 327250 148422
rect 327306 148366 327374 148422
rect 327430 148366 327498 148422
rect 327554 148366 327622 148422
rect 327678 148366 345250 148422
rect 345306 148366 345374 148422
rect 345430 148366 345498 148422
rect 345554 148366 345622 148422
rect 345678 148366 363250 148422
rect 363306 148366 363374 148422
rect 363430 148366 363498 148422
rect 363554 148366 363622 148422
rect 363678 148366 597980 148422
rect -1916 148350 597980 148366
rect -1916 148294 -860 148350
rect -804 148294 -736 148350
rect -680 148294 -612 148350
rect -556 148294 -488 148350
rect -432 148294 3250 148350
rect 3306 148294 3374 148350
rect 3430 148294 3498 148350
rect 3554 148294 3622 148350
rect 3678 148294 21250 148350
rect 21306 148294 21374 148350
rect 21430 148294 21498 148350
rect 21554 148294 21622 148350
rect 21678 148294 39250 148350
rect 39306 148294 39374 148350
rect 39430 148294 39498 148350
rect 39554 148294 39622 148350
rect 39678 148294 57250 148350
rect 57306 148294 57374 148350
rect 57430 148294 57498 148350
rect 57554 148294 57622 148350
rect 57678 148294 75250 148350
rect 75306 148294 75374 148350
rect 75430 148294 75498 148350
rect 75554 148294 75622 148350
rect 75678 148294 93250 148350
rect 93306 148294 93374 148350
rect 93430 148294 93498 148350
rect 93554 148294 93622 148350
rect 93678 148294 111250 148350
rect 111306 148294 111374 148350
rect 111430 148294 111498 148350
rect 111554 148294 111622 148350
rect 111678 148294 129250 148350
rect 129306 148294 129374 148350
rect 129430 148294 129498 148350
rect 129554 148294 129622 148350
rect 129678 148294 147250 148350
rect 147306 148294 147374 148350
rect 147430 148294 147498 148350
rect 147554 148294 147622 148350
rect 147678 148294 165250 148350
rect 165306 148294 165374 148350
rect 165430 148294 165498 148350
rect 165554 148294 165622 148350
rect 165678 148294 183250 148350
rect 183306 148294 183374 148350
rect 183430 148294 183498 148350
rect 183554 148294 183622 148350
rect 183678 148294 201250 148350
rect 201306 148294 201374 148350
rect 201430 148294 201498 148350
rect 201554 148294 201622 148350
rect 201678 148294 381250 148350
rect 381306 148294 381374 148350
rect 381430 148294 381498 148350
rect 381554 148294 381622 148350
rect 381678 148294 399250 148350
rect 399306 148294 399374 148350
rect 399430 148294 399498 148350
rect 399554 148294 399622 148350
rect 399678 148294 417250 148350
rect 417306 148294 417374 148350
rect 417430 148294 417498 148350
rect 417554 148294 417622 148350
rect 417678 148294 435250 148350
rect 435306 148294 435374 148350
rect 435430 148294 435498 148350
rect 435554 148294 435622 148350
rect 435678 148294 453250 148350
rect 453306 148294 453374 148350
rect 453430 148294 453498 148350
rect 453554 148294 453622 148350
rect 453678 148294 471250 148350
rect 471306 148294 471374 148350
rect 471430 148294 471498 148350
rect 471554 148294 471622 148350
rect 471678 148294 489250 148350
rect 489306 148294 489374 148350
rect 489430 148294 489498 148350
rect 489554 148294 489622 148350
rect 489678 148294 507250 148350
rect 507306 148294 507374 148350
rect 507430 148294 507498 148350
rect 507554 148294 507622 148350
rect 507678 148294 525250 148350
rect 525306 148294 525374 148350
rect 525430 148294 525498 148350
rect 525554 148294 525622 148350
rect 525678 148294 543250 148350
rect 543306 148294 543374 148350
rect 543430 148294 543498 148350
rect 543554 148294 543622 148350
rect 543678 148294 561250 148350
rect 561306 148294 561374 148350
rect 561430 148294 561498 148350
rect 561554 148294 561622 148350
rect 561678 148294 579250 148350
rect 579306 148294 579374 148350
rect 579430 148294 579498 148350
rect 579554 148294 579622 148350
rect 579678 148294 596496 148350
rect 596552 148294 596620 148350
rect 596676 148294 596744 148350
rect 596800 148294 596868 148350
rect 596924 148294 597980 148350
rect -1916 148226 597980 148294
rect -1916 148170 -860 148226
rect -804 148170 -736 148226
rect -680 148170 -612 148226
rect -556 148170 -488 148226
rect -432 148170 3250 148226
rect 3306 148170 3374 148226
rect 3430 148170 3498 148226
rect 3554 148170 3622 148226
rect 3678 148170 21250 148226
rect 21306 148170 21374 148226
rect 21430 148170 21498 148226
rect 21554 148170 21622 148226
rect 21678 148170 39250 148226
rect 39306 148170 39374 148226
rect 39430 148170 39498 148226
rect 39554 148170 39622 148226
rect 39678 148170 57250 148226
rect 57306 148170 57374 148226
rect 57430 148170 57498 148226
rect 57554 148170 57622 148226
rect 57678 148170 75250 148226
rect 75306 148170 75374 148226
rect 75430 148170 75498 148226
rect 75554 148170 75622 148226
rect 75678 148170 93250 148226
rect 93306 148170 93374 148226
rect 93430 148170 93498 148226
rect 93554 148170 93622 148226
rect 93678 148170 111250 148226
rect 111306 148170 111374 148226
rect 111430 148170 111498 148226
rect 111554 148170 111622 148226
rect 111678 148170 129250 148226
rect 129306 148170 129374 148226
rect 129430 148170 129498 148226
rect 129554 148170 129622 148226
rect 129678 148170 147250 148226
rect 147306 148170 147374 148226
rect 147430 148170 147498 148226
rect 147554 148170 147622 148226
rect 147678 148170 165250 148226
rect 165306 148170 165374 148226
rect 165430 148170 165498 148226
rect 165554 148170 165622 148226
rect 165678 148170 183250 148226
rect 183306 148170 183374 148226
rect 183430 148170 183498 148226
rect 183554 148170 183622 148226
rect 183678 148170 201250 148226
rect 201306 148170 201374 148226
rect 201430 148170 201498 148226
rect 201554 148170 201622 148226
rect 201678 148170 381250 148226
rect 381306 148170 381374 148226
rect 381430 148170 381498 148226
rect 381554 148170 381622 148226
rect 381678 148170 399250 148226
rect 399306 148170 399374 148226
rect 399430 148170 399498 148226
rect 399554 148170 399622 148226
rect 399678 148170 417250 148226
rect 417306 148170 417374 148226
rect 417430 148170 417498 148226
rect 417554 148170 417622 148226
rect 417678 148170 435250 148226
rect 435306 148170 435374 148226
rect 435430 148170 435498 148226
rect 435554 148170 435622 148226
rect 435678 148170 453250 148226
rect 453306 148170 453374 148226
rect 453430 148170 453498 148226
rect 453554 148170 453622 148226
rect 453678 148170 471250 148226
rect 471306 148170 471374 148226
rect 471430 148170 471498 148226
rect 471554 148170 471622 148226
rect 471678 148170 489250 148226
rect 489306 148170 489374 148226
rect 489430 148170 489498 148226
rect 489554 148170 489622 148226
rect 489678 148170 507250 148226
rect 507306 148170 507374 148226
rect 507430 148170 507498 148226
rect 507554 148170 507622 148226
rect 507678 148170 525250 148226
rect 525306 148170 525374 148226
rect 525430 148170 525498 148226
rect 525554 148170 525622 148226
rect 525678 148170 543250 148226
rect 543306 148170 543374 148226
rect 543430 148170 543498 148226
rect 543554 148170 543622 148226
rect 543678 148170 561250 148226
rect 561306 148170 561374 148226
rect 561430 148170 561498 148226
rect 561554 148170 561622 148226
rect 561678 148170 579250 148226
rect 579306 148170 579374 148226
rect 579430 148170 579498 148226
rect 579554 148170 579622 148226
rect 579678 148170 596496 148226
rect 596552 148170 596620 148226
rect 596676 148170 596744 148226
rect 596800 148170 596868 148226
rect 596924 148170 597980 148226
rect -1916 148102 597980 148170
rect -1916 148046 -860 148102
rect -804 148046 -736 148102
rect -680 148046 -612 148102
rect -556 148046 -488 148102
rect -432 148046 3250 148102
rect 3306 148046 3374 148102
rect 3430 148046 3498 148102
rect 3554 148046 3622 148102
rect 3678 148046 21250 148102
rect 21306 148046 21374 148102
rect 21430 148046 21498 148102
rect 21554 148046 21622 148102
rect 21678 148046 39250 148102
rect 39306 148046 39374 148102
rect 39430 148046 39498 148102
rect 39554 148046 39622 148102
rect 39678 148046 57250 148102
rect 57306 148046 57374 148102
rect 57430 148046 57498 148102
rect 57554 148046 57622 148102
rect 57678 148046 75250 148102
rect 75306 148046 75374 148102
rect 75430 148046 75498 148102
rect 75554 148046 75622 148102
rect 75678 148046 93250 148102
rect 93306 148046 93374 148102
rect 93430 148046 93498 148102
rect 93554 148046 93622 148102
rect 93678 148046 111250 148102
rect 111306 148046 111374 148102
rect 111430 148046 111498 148102
rect 111554 148046 111622 148102
rect 111678 148046 129250 148102
rect 129306 148046 129374 148102
rect 129430 148046 129498 148102
rect 129554 148046 129622 148102
rect 129678 148046 147250 148102
rect 147306 148046 147374 148102
rect 147430 148046 147498 148102
rect 147554 148046 147622 148102
rect 147678 148046 165250 148102
rect 165306 148046 165374 148102
rect 165430 148046 165498 148102
rect 165554 148046 165622 148102
rect 165678 148046 183250 148102
rect 183306 148046 183374 148102
rect 183430 148046 183498 148102
rect 183554 148046 183622 148102
rect 183678 148046 201250 148102
rect 201306 148046 201374 148102
rect 201430 148046 201498 148102
rect 201554 148046 201622 148102
rect 201678 148046 381250 148102
rect 381306 148046 381374 148102
rect 381430 148046 381498 148102
rect 381554 148046 381622 148102
rect 381678 148046 399250 148102
rect 399306 148046 399374 148102
rect 399430 148046 399498 148102
rect 399554 148046 399622 148102
rect 399678 148046 417250 148102
rect 417306 148046 417374 148102
rect 417430 148046 417498 148102
rect 417554 148046 417622 148102
rect 417678 148046 435250 148102
rect 435306 148046 435374 148102
rect 435430 148046 435498 148102
rect 435554 148046 435622 148102
rect 435678 148046 453250 148102
rect 453306 148046 453374 148102
rect 453430 148046 453498 148102
rect 453554 148046 453622 148102
rect 453678 148046 471250 148102
rect 471306 148046 471374 148102
rect 471430 148046 471498 148102
rect 471554 148046 471622 148102
rect 471678 148046 489250 148102
rect 489306 148046 489374 148102
rect 489430 148046 489498 148102
rect 489554 148046 489622 148102
rect 489678 148046 507250 148102
rect 507306 148046 507374 148102
rect 507430 148046 507498 148102
rect 507554 148046 507622 148102
rect 507678 148046 525250 148102
rect 525306 148046 525374 148102
rect 525430 148046 525498 148102
rect 525554 148046 525622 148102
rect 525678 148046 543250 148102
rect 543306 148046 543374 148102
rect 543430 148046 543498 148102
rect 543554 148046 543622 148102
rect 543678 148046 561250 148102
rect 561306 148046 561374 148102
rect 561430 148046 561498 148102
rect 561554 148046 561622 148102
rect 561678 148046 579250 148102
rect 579306 148046 579374 148102
rect 579430 148046 579498 148102
rect 579554 148046 579622 148102
rect 579678 148046 596496 148102
rect 596552 148046 596620 148102
rect 596676 148046 596744 148102
rect 596800 148046 596868 148102
rect 596924 148046 597980 148102
rect -1916 147978 597980 148046
rect -1916 147922 -860 147978
rect -804 147922 -736 147978
rect -680 147922 -612 147978
rect -556 147922 -488 147978
rect -432 147922 3250 147978
rect 3306 147922 3374 147978
rect 3430 147922 3498 147978
rect 3554 147922 3622 147978
rect 3678 147922 21250 147978
rect 21306 147922 21374 147978
rect 21430 147922 21498 147978
rect 21554 147922 21622 147978
rect 21678 147922 39250 147978
rect 39306 147922 39374 147978
rect 39430 147922 39498 147978
rect 39554 147922 39622 147978
rect 39678 147922 57250 147978
rect 57306 147922 57374 147978
rect 57430 147922 57498 147978
rect 57554 147922 57622 147978
rect 57678 147922 75250 147978
rect 75306 147922 75374 147978
rect 75430 147922 75498 147978
rect 75554 147922 75622 147978
rect 75678 147922 93250 147978
rect 93306 147922 93374 147978
rect 93430 147922 93498 147978
rect 93554 147922 93622 147978
rect 93678 147922 111250 147978
rect 111306 147922 111374 147978
rect 111430 147922 111498 147978
rect 111554 147922 111622 147978
rect 111678 147922 129250 147978
rect 129306 147922 129374 147978
rect 129430 147922 129498 147978
rect 129554 147922 129622 147978
rect 129678 147922 147250 147978
rect 147306 147922 147374 147978
rect 147430 147922 147498 147978
rect 147554 147922 147622 147978
rect 147678 147922 165250 147978
rect 165306 147922 165374 147978
rect 165430 147922 165498 147978
rect 165554 147922 165622 147978
rect 165678 147922 183250 147978
rect 183306 147922 183374 147978
rect 183430 147922 183498 147978
rect 183554 147922 183622 147978
rect 183678 147922 201250 147978
rect 201306 147922 201374 147978
rect 201430 147922 201498 147978
rect 201554 147922 201622 147978
rect 201678 147922 381250 147978
rect 381306 147922 381374 147978
rect 381430 147922 381498 147978
rect 381554 147922 381622 147978
rect 381678 147922 399250 147978
rect 399306 147922 399374 147978
rect 399430 147922 399498 147978
rect 399554 147922 399622 147978
rect 399678 147922 417250 147978
rect 417306 147922 417374 147978
rect 417430 147922 417498 147978
rect 417554 147922 417622 147978
rect 417678 147922 435250 147978
rect 435306 147922 435374 147978
rect 435430 147922 435498 147978
rect 435554 147922 435622 147978
rect 435678 147922 453250 147978
rect 453306 147922 453374 147978
rect 453430 147922 453498 147978
rect 453554 147922 453622 147978
rect 453678 147922 471250 147978
rect 471306 147922 471374 147978
rect 471430 147922 471498 147978
rect 471554 147922 471622 147978
rect 471678 147922 489250 147978
rect 489306 147922 489374 147978
rect 489430 147922 489498 147978
rect 489554 147922 489622 147978
rect 489678 147922 507250 147978
rect 507306 147922 507374 147978
rect 507430 147922 507498 147978
rect 507554 147922 507622 147978
rect 507678 147922 525250 147978
rect 525306 147922 525374 147978
rect 525430 147922 525498 147978
rect 525554 147922 525622 147978
rect 525678 147922 543250 147978
rect 543306 147922 543374 147978
rect 543430 147922 543498 147978
rect 543554 147922 543622 147978
rect 543678 147922 561250 147978
rect 561306 147922 561374 147978
rect 561430 147922 561498 147978
rect 561554 147922 561622 147978
rect 561678 147922 579250 147978
rect 579306 147922 579374 147978
rect 579430 147922 579498 147978
rect 579554 147922 579622 147978
rect 579678 147922 596496 147978
rect 596552 147922 596620 147978
rect 596676 147922 596744 147978
rect 596800 147922 596868 147978
rect 596924 147922 597980 147978
rect -1916 147826 597980 147922
rect -1916 136350 597980 136446
rect -1916 136294 -1820 136350
rect -1764 136294 -1696 136350
rect -1640 136294 -1572 136350
rect -1516 136294 -1448 136350
rect -1392 136294 6970 136350
rect 7026 136294 7094 136350
rect 7150 136294 7218 136350
rect 7274 136294 7342 136350
rect 7398 136294 24970 136350
rect 25026 136294 25094 136350
rect 25150 136294 25218 136350
rect 25274 136294 25342 136350
rect 25398 136294 42970 136350
rect 43026 136294 43094 136350
rect 43150 136294 43218 136350
rect 43274 136294 43342 136350
rect 43398 136294 60970 136350
rect 61026 136294 61094 136350
rect 61150 136294 61218 136350
rect 61274 136294 61342 136350
rect 61398 136294 78970 136350
rect 79026 136294 79094 136350
rect 79150 136294 79218 136350
rect 79274 136294 79342 136350
rect 79398 136294 96970 136350
rect 97026 136294 97094 136350
rect 97150 136294 97218 136350
rect 97274 136294 97342 136350
rect 97398 136294 114970 136350
rect 115026 136294 115094 136350
rect 115150 136294 115218 136350
rect 115274 136294 115342 136350
rect 115398 136294 132970 136350
rect 133026 136294 133094 136350
rect 133150 136294 133218 136350
rect 133274 136294 133342 136350
rect 133398 136294 150970 136350
rect 151026 136294 151094 136350
rect 151150 136294 151218 136350
rect 151274 136294 151342 136350
rect 151398 136294 168970 136350
rect 169026 136294 169094 136350
rect 169150 136294 169218 136350
rect 169274 136294 169342 136350
rect 169398 136294 186970 136350
rect 187026 136294 187094 136350
rect 187150 136294 187218 136350
rect 187274 136294 187342 136350
rect 187398 136294 204970 136350
rect 205026 136294 205094 136350
rect 205150 136294 205218 136350
rect 205274 136294 205342 136350
rect 205398 136294 384970 136350
rect 385026 136294 385094 136350
rect 385150 136294 385218 136350
rect 385274 136294 385342 136350
rect 385398 136294 402970 136350
rect 403026 136294 403094 136350
rect 403150 136294 403218 136350
rect 403274 136294 403342 136350
rect 403398 136294 420970 136350
rect 421026 136294 421094 136350
rect 421150 136294 421218 136350
rect 421274 136294 421342 136350
rect 421398 136294 438970 136350
rect 439026 136294 439094 136350
rect 439150 136294 439218 136350
rect 439274 136294 439342 136350
rect 439398 136294 456970 136350
rect 457026 136294 457094 136350
rect 457150 136294 457218 136350
rect 457274 136294 457342 136350
rect 457398 136294 474970 136350
rect 475026 136294 475094 136350
rect 475150 136294 475218 136350
rect 475274 136294 475342 136350
rect 475398 136294 492970 136350
rect 493026 136294 493094 136350
rect 493150 136294 493218 136350
rect 493274 136294 493342 136350
rect 493398 136294 510970 136350
rect 511026 136294 511094 136350
rect 511150 136294 511218 136350
rect 511274 136294 511342 136350
rect 511398 136294 528970 136350
rect 529026 136294 529094 136350
rect 529150 136294 529218 136350
rect 529274 136294 529342 136350
rect 529398 136294 546970 136350
rect 547026 136294 547094 136350
rect 547150 136294 547218 136350
rect 547274 136294 547342 136350
rect 547398 136294 564970 136350
rect 565026 136294 565094 136350
rect 565150 136294 565218 136350
rect 565274 136294 565342 136350
rect 565398 136294 582970 136350
rect 583026 136294 583094 136350
rect 583150 136294 583218 136350
rect 583274 136294 583342 136350
rect 583398 136294 597456 136350
rect 597512 136294 597580 136350
rect 597636 136294 597704 136350
rect 597760 136294 597828 136350
rect 597884 136294 597980 136350
rect -1916 136226 597980 136294
rect -1916 136170 -1820 136226
rect -1764 136170 -1696 136226
rect -1640 136170 -1572 136226
rect -1516 136170 -1448 136226
rect -1392 136170 6970 136226
rect 7026 136170 7094 136226
rect 7150 136170 7218 136226
rect 7274 136170 7342 136226
rect 7398 136170 24970 136226
rect 25026 136170 25094 136226
rect 25150 136170 25218 136226
rect 25274 136170 25342 136226
rect 25398 136170 42970 136226
rect 43026 136170 43094 136226
rect 43150 136170 43218 136226
rect 43274 136170 43342 136226
rect 43398 136170 60970 136226
rect 61026 136170 61094 136226
rect 61150 136170 61218 136226
rect 61274 136170 61342 136226
rect 61398 136170 78970 136226
rect 79026 136170 79094 136226
rect 79150 136170 79218 136226
rect 79274 136170 79342 136226
rect 79398 136170 96970 136226
rect 97026 136170 97094 136226
rect 97150 136170 97218 136226
rect 97274 136170 97342 136226
rect 97398 136170 114970 136226
rect 115026 136170 115094 136226
rect 115150 136170 115218 136226
rect 115274 136170 115342 136226
rect 115398 136170 132970 136226
rect 133026 136170 133094 136226
rect 133150 136170 133218 136226
rect 133274 136170 133342 136226
rect 133398 136170 150970 136226
rect 151026 136170 151094 136226
rect 151150 136170 151218 136226
rect 151274 136170 151342 136226
rect 151398 136170 168970 136226
rect 169026 136170 169094 136226
rect 169150 136170 169218 136226
rect 169274 136170 169342 136226
rect 169398 136170 186970 136226
rect 187026 136170 187094 136226
rect 187150 136170 187218 136226
rect 187274 136170 187342 136226
rect 187398 136170 204970 136226
rect 205026 136170 205094 136226
rect 205150 136170 205218 136226
rect 205274 136170 205342 136226
rect 205398 136170 384970 136226
rect 385026 136170 385094 136226
rect 385150 136170 385218 136226
rect 385274 136170 385342 136226
rect 385398 136170 402970 136226
rect 403026 136170 403094 136226
rect 403150 136170 403218 136226
rect 403274 136170 403342 136226
rect 403398 136170 420970 136226
rect 421026 136170 421094 136226
rect 421150 136170 421218 136226
rect 421274 136170 421342 136226
rect 421398 136170 438970 136226
rect 439026 136170 439094 136226
rect 439150 136170 439218 136226
rect 439274 136170 439342 136226
rect 439398 136170 456970 136226
rect 457026 136170 457094 136226
rect 457150 136170 457218 136226
rect 457274 136170 457342 136226
rect 457398 136170 474970 136226
rect 475026 136170 475094 136226
rect 475150 136170 475218 136226
rect 475274 136170 475342 136226
rect 475398 136170 492970 136226
rect 493026 136170 493094 136226
rect 493150 136170 493218 136226
rect 493274 136170 493342 136226
rect 493398 136170 510970 136226
rect 511026 136170 511094 136226
rect 511150 136170 511218 136226
rect 511274 136170 511342 136226
rect 511398 136170 528970 136226
rect 529026 136170 529094 136226
rect 529150 136170 529218 136226
rect 529274 136170 529342 136226
rect 529398 136170 546970 136226
rect 547026 136170 547094 136226
rect 547150 136170 547218 136226
rect 547274 136170 547342 136226
rect 547398 136170 564970 136226
rect 565026 136170 565094 136226
rect 565150 136170 565218 136226
rect 565274 136170 565342 136226
rect 565398 136170 582970 136226
rect 583026 136170 583094 136226
rect 583150 136170 583218 136226
rect 583274 136170 583342 136226
rect 583398 136170 597456 136226
rect 597512 136170 597580 136226
rect 597636 136170 597704 136226
rect 597760 136170 597828 136226
rect 597884 136170 597980 136226
rect -1916 136102 597980 136170
rect -1916 136046 -1820 136102
rect -1764 136046 -1696 136102
rect -1640 136046 -1572 136102
rect -1516 136046 -1448 136102
rect -1392 136046 6970 136102
rect 7026 136046 7094 136102
rect 7150 136046 7218 136102
rect 7274 136046 7342 136102
rect 7398 136046 24970 136102
rect 25026 136046 25094 136102
rect 25150 136046 25218 136102
rect 25274 136046 25342 136102
rect 25398 136046 42970 136102
rect 43026 136046 43094 136102
rect 43150 136046 43218 136102
rect 43274 136046 43342 136102
rect 43398 136046 60970 136102
rect 61026 136046 61094 136102
rect 61150 136046 61218 136102
rect 61274 136046 61342 136102
rect 61398 136046 78970 136102
rect 79026 136046 79094 136102
rect 79150 136046 79218 136102
rect 79274 136046 79342 136102
rect 79398 136046 96970 136102
rect 97026 136046 97094 136102
rect 97150 136046 97218 136102
rect 97274 136046 97342 136102
rect 97398 136046 114970 136102
rect 115026 136046 115094 136102
rect 115150 136046 115218 136102
rect 115274 136046 115342 136102
rect 115398 136046 132970 136102
rect 133026 136046 133094 136102
rect 133150 136046 133218 136102
rect 133274 136046 133342 136102
rect 133398 136046 150970 136102
rect 151026 136046 151094 136102
rect 151150 136046 151218 136102
rect 151274 136046 151342 136102
rect 151398 136046 168970 136102
rect 169026 136046 169094 136102
rect 169150 136046 169218 136102
rect 169274 136046 169342 136102
rect 169398 136046 186970 136102
rect 187026 136046 187094 136102
rect 187150 136046 187218 136102
rect 187274 136046 187342 136102
rect 187398 136046 204970 136102
rect 205026 136046 205094 136102
rect 205150 136046 205218 136102
rect 205274 136046 205342 136102
rect 205398 136046 384970 136102
rect 385026 136046 385094 136102
rect 385150 136046 385218 136102
rect 385274 136046 385342 136102
rect 385398 136046 402970 136102
rect 403026 136046 403094 136102
rect 403150 136046 403218 136102
rect 403274 136046 403342 136102
rect 403398 136046 420970 136102
rect 421026 136046 421094 136102
rect 421150 136046 421218 136102
rect 421274 136046 421342 136102
rect 421398 136046 438970 136102
rect 439026 136046 439094 136102
rect 439150 136046 439218 136102
rect 439274 136046 439342 136102
rect 439398 136046 456970 136102
rect 457026 136046 457094 136102
rect 457150 136046 457218 136102
rect 457274 136046 457342 136102
rect 457398 136046 474970 136102
rect 475026 136046 475094 136102
rect 475150 136046 475218 136102
rect 475274 136046 475342 136102
rect 475398 136046 492970 136102
rect 493026 136046 493094 136102
rect 493150 136046 493218 136102
rect 493274 136046 493342 136102
rect 493398 136046 510970 136102
rect 511026 136046 511094 136102
rect 511150 136046 511218 136102
rect 511274 136046 511342 136102
rect 511398 136046 528970 136102
rect 529026 136046 529094 136102
rect 529150 136046 529218 136102
rect 529274 136046 529342 136102
rect 529398 136046 546970 136102
rect 547026 136046 547094 136102
rect 547150 136046 547218 136102
rect 547274 136046 547342 136102
rect 547398 136046 564970 136102
rect 565026 136046 565094 136102
rect 565150 136046 565218 136102
rect 565274 136046 565342 136102
rect 565398 136046 582970 136102
rect 583026 136046 583094 136102
rect 583150 136046 583218 136102
rect 583274 136046 583342 136102
rect 583398 136046 597456 136102
rect 597512 136046 597580 136102
rect 597636 136046 597704 136102
rect 597760 136046 597828 136102
rect 597884 136046 597980 136102
rect -1916 135978 597980 136046
rect -1916 135922 -1820 135978
rect -1764 135922 -1696 135978
rect -1640 135922 -1572 135978
rect -1516 135922 -1448 135978
rect -1392 135922 6970 135978
rect 7026 135922 7094 135978
rect 7150 135922 7218 135978
rect 7274 135922 7342 135978
rect 7398 135922 24970 135978
rect 25026 135922 25094 135978
rect 25150 135922 25218 135978
rect 25274 135922 25342 135978
rect 25398 135922 42970 135978
rect 43026 135922 43094 135978
rect 43150 135922 43218 135978
rect 43274 135922 43342 135978
rect 43398 135922 60970 135978
rect 61026 135922 61094 135978
rect 61150 135922 61218 135978
rect 61274 135922 61342 135978
rect 61398 135922 78970 135978
rect 79026 135922 79094 135978
rect 79150 135922 79218 135978
rect 79274 135922 79342 135978
rect 79398 135922 96970 135978
rect 97026 135922 97094 135978
rect 97150 135922 97218 135978
rect 97274 135922 97342 135978
rect 97398 135922 114970 135978
rect 115026 135922 115094 135978
rect 115150 135922 115218 135978
rect 115274 135922 115342 135978
rect 115398 135922 132970 135978
rect 133026 135922 133094 135978
rect 133150 135922 133218 135978
rect 133274 135922 133342 135978
rect 133398 135922 150970 135978
rect 151026 135922 151094 135978
rect 151150 135922 151218 135978
rect 151274 135922 151342 135978
rect 151398 135922 168970 135978
rect 169026 135922 169094 135978
rect 169150 135922 169218 135978
rect 169274 135922 169342 135978
rect 169398 135922 186970 135978
rect 187026 135922 187094 135978
rect 187150 135922 187218 135978
rect 187274 135922 187342 135978
rect 187398 135922 204970 135978
rect 205026 135922 205094 135978
rect 205150 135922 205218 135978
rect 205274 135922 205342 135978
rect 205398 135922 384970 135978
rect 385026 135922 385094 135978
rect 385150 135922 385218 135978
rect 385274 135922 385342 135978
rect 385398 135922 402970 135978
rect 403026 135922 403094 135978
rect 403150 135922 403218 135978
rect 403274 135922 403342 135978
rect 403398 135922 420970 135978
rect 421026 135922 421094 135978
rect 421150 135922 421218 135978
rect 421274 135922 421342 135978
rect 421398 135922 438970 135978
rect 439026 135922 439094 135978
rect 439150 135922 439218 135978
rect 439274 135922 439342 135978
rect 439398 135922 456970 135978
rect 457026 135922 457094 135978
rect 457150 135922 457218 135978
rect 457274 135922 457342 135978
rect 457398 135922 474970 135978
rect 475026 135922 475094 135978
rect 475150 135922 475218 135978
rect 475274 135922 475342 135978
rect 475398 135922 492970 135978
rect 493026 135922 493094 135978
rect 493150 135922 493218 135978
rect 493274 135922 493342 135978
rect 493398 135922 510970 135978
rect 511026 135922 511094 135978
rect 511150 135922 511218 135978
rect 511274 135922 511342 135978
rect 511398 135922 528970 135978
rect 529026 135922 529094 135978
rect 529150 135922 529218 135978
rect 529274 135922 529342 135978
rect 529398 135922 546970 135978
rect 547026 135922 547094 135978
rect 547150 135922 547218 135978
rect 547274 135922 547342 135978
rect 547398 135922 564970 135978
rect 565026 135922 565094 135978
rect 565150 135922 565218 135978
rect 565274 135922 565342 135978
rect 565398 135922 582970 135978
rect 583026 135922 583094 135978
rect 583150 135922 583218 135978
rect 583274 135922 583342 135978
rect 583398 135922 597456 135978
rect 597512 135922 597580 135978
rect 597636 135922 597704 135978
rect 597760 135922 597828 135978
rect 597884 135922 597980 135978
rect -1916 135826 597980 135922
rect -1916 130350 597980 130446
rect -1916 130294 -860 130350
rect -804 130294 -736 130350
rect -680 130294 -612 130350
rect -556 130294 -488 130350
rect -432 130294 3250 130350
rect 3306 130294 3374 130350
rect 3430 130294 3498 130350
rect 3554 130294 3622 130350
rect 3678 130294 21250 130350
rect 21306 130294 21374 130350
rect 21430 130294 21498 130350
rect 21554 130294 21622 130350
rect 21678 130294 39250 130350
rect 39306 130294 39374 130350
rect 39430 130294 39498 130350
rect 39554 130294 39622 130350
rect 39678 130294 57250 130350
rect 57306 130294 57374 130350
rect 57430 130294 57498 130350
rect 57554 130294 57622 130350
rect 57678 130294 75250 130350
rect 75306 130294 75374 130350
rect 75430 130294 75498 130350
rect 75554 130294 75622 130350
rect 75678 130294 93250 130350
rect 93306 130294 93374 130350
rect 93430 130294 93498 130350
rect 93554 130294 93622 130350
rect 93678 130294 111250 130350
rect 111306 130294 111374 130350
rect 111430 130294 111498 130350
rect 111554 130294 111622 130350
rect 111678 130294 129250 130350
rect 129306 130294 129374 130350
rect 129430 130294 129498 130350
rect 129554 130294 129622 130350
rect 129678 130294 147250 130350
rect 147306 130294 147374 130350
rect 147430 130294 147498 130350
rect 147554 130294 147622 130350
rect 147678 130294 165250 130350
rect 165306 130294 165374 130350
rect 165430 130294 165498 130350
rect 165554 130294 165622 130350
rect 165678 130294 183250 130350
rect 183306 130294 183374 130350
rect 183430 130294 183498 130350
rect 183554 130294 183622 130350
rect 183678 130294 201250 130350
rect 201306 130294 201374 130350
rect 201430 130294 201498 130350
rect 201554 130294 201622 130350
rect 201678 130294 381250 130350
rect 381306 130294 381374 130350
rect 381430 130294 381498 130350
rect 381554 130294 381622 130350
rect 381678 130294 399250 130350
rect 399306 130294 399374 130350
rect 399430 130294 399498 130350
rect 399554 130294 399622 130350
rect 399678 130294 417250 130350
rect 417306 130294 417374 130350
rect 417430 130294 417498 130350
rect 417554 130294 417622 130350
rect 417678 130294 435250 130350
rect 435306 130294 435374 130350
rect 435430 130294 435498 130350
rect 435554 130294 435622 130350
rect 435678 130294 453250 130350
rect 453306 130294 453374 130350
rect 453430 130294 453498 130350
rect 453554 130294 453622 130350
rect 453678 130294 471250 130350
rect 471306 130294 471374 130350
rect 471430 130294 471498 130350
rect 471554 130294 471622 130350
rect 471678 130294 489250 130350
rect 489306 130294 489374 130350
rect 489430 130294 489498 130350
rect 489554 130294 489622 130350
rect 489678 130294 507250 130350
rect 507306 130294 507374 130350
rect 507430 130294 507498 130350
rect 507554 130294 507622 130350
rect 507678 130294 525250 130350
rect 525306 130294 525374 130350
rect 525430 130294 525498 130350
rect 525554 130294 525622 130350
rect 525678 130294 543250 130350
rect 543306 130294 543374 130350
rect 543430 130294 543498 130350
rect 543554 130294 543622 130350
rect 543678 130294 561250 130350
rect 561306 130294 561374 130350
rect 561430 130294 561498 130350
rect 561554 130294 561622 130350
rect 561678 130294 579250 130350
rect 579306 130294 579374 130350
rect 579430 130294 579498 130350
rect 579554 130294 579622 130350
rect 579678 130294 596496 130350
rect 596552 130294 596620 130350
rect 596676 130294 596744 130350
rect 596800 130294 596868 130350
rect 596924 130294 597980 130350
rect -1916 130226 597980 130294
rect -1916 130170 -860 130226
rect -804 130170 -736 130226
rect -680 130170 -612 130226
rect -556 130170 -488 130226
rect -432 130170 3250 130226
rect 3306 130170 3374 130226
rect 3430 130170 3498 130226
rect 3554 130170 3622 130226
rect 3678 130170 21250 130226
rect 21306 130170 21374 130226
rect 21430 130170 21498 130226
rect 21554 130170 21622 130226
rect 21678 130170 39250 130226
rect 39306 130170 39374 130226
rect 39430 130170 39498 130226
rect 39554 130170 39622 130226
rect 39678 130170 57250 130226
rect 57306 130170 57374 130226
rect 57430 130170 57498 130226
rect 57554 130170 57622 130226
rect 57678 130170 75250 130226
rect 75306 130170 75374 130226
rect 75430 130170 75498 130226
rect 75554 130170 75622 130226
rect 75678 130170 93250 130226
rect 93306 130170 93374 130226
rect 93430 130170 93498 130226
rect 93554 130170 93622 130226
rect 93678 130170 111250 130226
rect 111306 130170 111374 130226
rect 111430 130170 111498 130226
rect 111554 130170 111622 130226
rect 111678 130170 129250 130226
rect 129306 130170 129374 130226
rect 129430 130170 129498 130226
rect 129554 130170 129622 130226
rect 129678 130170 147250 130226
rect 147306 130170 147374 130226
rect 147430 130170 147498 130226
rect 147554 130170 147622 130226
rect 147678 130170 165250 130226
rect 165306 130170 165374 130226
rect 165430 130170 165498 130226
rect 165554 130170 165622 130226
rect 165678 130170 183250 130226
rect 183306 130170 183374 130226
rect 183430 130170 183498 130226
rect 183554 130170 183622 130226
rect 183678 130170 201250 130226
rect 201306 130170 201374 130226
rect 201430 130170 201498 130226
rect 201554 130170 201622 130226
rect 201678 130170 381250 130226
rect 381306 130170 381374 130226
rect 381430 130170 381498 130226
rect 381554 130170 381622 130226
rect 381678 130170 399250 130226
rect 399306 130170 399374 130226
rect 399430 130170 399498 130226
rect 399554 130170 399622 130226
rect 399678 130170 417250 130226
rect 417306 130170 417374 130226
rect 417430 130170 417498 130226
rect 417554 130170 417622 130226
rect 417678 130170 435250 130226
rect 435306 130170 435374 130226
rect 435430 130170 435498 130226
rect 435554 130170 435622 130226
rect 435678 130170 453250 130226
rect 453306 130170 453374 130226
rect 453430 130170 453498 130226
rect 453554 130170 453622 130226
rect 453678 130170 471250 130226
rect 471306 130170 471374 130226
rect 471430 130170 471498 130226
rect 471554 130170 471622 130226
rect 471678 130170 489250 130226
rect 489306 130170 489374 130226
rect 489430 130170 489498 130226
rect 489554 130170 489622 130226
rect 489678 130170 507250 130226
rect 507306 130170 507374 130226
rect 507430 130170 507498 130226
rect 507554 130170 507622 130226
rect 507678 130170 525250 130226
rect 525306 130170 525374 130226
rect 525430 130170 525498 130226
rect 525554 130170 525622 130226
rect 525678 130170 543250 130226
rect 543306 130170 543374 130226
rect 543430 130170 543498 130226
rect 543554 130170 543622 130226
rect 543678 130170 561250 130226
rect 561306 130170 561374 130226
rect 561430 130170 561498 130226
rect 561554 130170 561622 130226
rect 561678 130170 579250 130226
rect 579306 130170 579374 130226
rect 579430 130170 579498 130226
rect 579554 130170 579622 130226
rect 579678 130170 596496 130226
rect 596552 130170 596620 130226
rect 596676 130170 596744 130226
rect 596800 130170 596868 130226
rect 596924 130170 597980 130226
rect -1916 130102 597980 130170
rect -1916 130046 -860 130102
rect -804 130046 -736 130102
rect -680 130046 -612 130102
rect -556 130046 -488 130102
rect -432 130046 3250 130102
rect 3306 130046 3374 130102
rect 3430 130046 3498 130102
rect 3554 130046 3622 130102
rect 3678 130046 21250 130102
rect 21306 130046 21374 130102
rect 21430 130046 21498 130102
rect 21554 130046 21622 130102
rect 21678 130046 39250 130102
rect 39306 130046 39374 130102
rect 39430 130046 39498 130102
rect 39554 130046 39622 130102
rect 39678 130046 57250 130102
rect 57306 130046 57374 130102
rect 57430 130046 57498 130102
rect 57554 130046 57622 130102
rect 57678 130046 75250 130102
rect 75306 130046 75374 130102
rect 75430 130046 75498 130102
rect 75554 130046 75622 130102
rect 75678 130046 93250 130102
rect 93306 130046 93374 130102
rect 93430 130046 93498 130102
rect 93554 130046 93622 130102
rect 93678 130046 111250 130102
rect 111306 130046 111374 130102
rect 111430 130046 111498 130102
rect 111554 130046 111622 130102
rect 111678 130046 129250 130102
rect 129306 130046 129374 130102
rect 129430 130046 129498 130102
rect 129554 130046 129622 130102
rect 129678 130046 147250 130102
rect 147306 130046 147374 130102
rect 147430 130046 147498 130102
rect 147554 130046 147622 130102
rect 147678 130046 165250 130102
rect 165306 130046 165374 130102
rect 165430 130046 165498 130102
rect 165554 130046 165622 130102
rect 165678 130046 183250 130102
rect 183306 130046 183374 130102
rect 183430 130046 183498 130102
rect 183554 130046 183622 130102
rect 183678 130046 201250 130102
rect 201306 130046 201374 130102
rect 201430 130046 201498 130102
rect 201554 130046 201622 130102
rect 201678 130046 381250 130102
rect 381306 130046 381374 130102
rect 381430 130046 381498 130102
rect 381554 130046 381622 130102
rect 381678 130046 399250 130102
rect 399306 130046 399374 130102
rect 399430 130046 399498 130102
rect 399554 130046 399622 130102
rect 399678 130046 417250 130102
rect 417306 130046 417374 130102
rect 417430 130046 417498 130102
rect 417554 130046 417622 130102
rect 417678 130046 435250 130102
rect 435306 130046 435374 130102
rect 435430 130046 435498 130102
rect 435554 130046 435622 130102
rect 435678 130046 453250 130102
rect 453306 130046 453374 130102
rect 453430 130046 453498 130102
rect 453554 130046 453622 130102
rect 453678 130046 471250 130102
rect 471306 130046 471374 130102
rect 471430 130046 471498 130102
rect 471554 130046 471622 130102
rect 471678 130046 489250 130102
rect 489306 130046 489374 130102
rect 489430 130046 489498 130102
rect 489554 130046 489622 130102
rect 489678 130046 507250 130102
rect 507306 130046 507374 130102
rect 507430 130046 507498 130102
rect 507554 130046 507622 130102
rect 507678 130046 525250 130102
rect 525306 130046 525374 130102
rect 525430 130046 525498 130102
rect 525554 130046 525622 130102
rect 525678 130046 543250 130102
rect 543306 130046 543374 130102
rect 543430 130046 543498 130102
rect 543554 130046 543622 130102
rect 543678 130046 561250 130102
rect 561306 130046 561374 130102
rect 561430 130046 561498 130102
rect 561554 130046 561622 130102
rect 561678 130046 579250 130102
rect 579306 130046 579374 130102
rect 579430 130046 579498 130102
rect 579554 130046 579622 130102
rect 579678 130046 596496 130102
rect 596552 130046 596620 130102
rect 596676 130046 596744 130102
rect 596800 130046 596868 130102
rect 596924 130046 597980 130102
rect -1916 129978 597980 130046
rect -1916 129922 -860 129978
rect -804 129922 -736 129978
rect -680 129922 -612 129978
rect -556 129922 -488 129978
rect -432 129922 3250 129978
rect 3306 129922 3374 129978
rect 3430 129922 3498 129978
rect 3554 129922 3622 129978
rect 3678 129922 21250 129978
rect 21306 129922 21374 129978
rect 21430 129922 21498 129978
rect 21554 129922 21622 129978
rect 21678 129922 39250 129978
rect 39306 129922 39374 129978
rect 39430 129922 39498 129978
rect 39554 129922 39622 129978
rect 39678 129922 57250 129978
rect 57306 129922 57374 129978
rect 57430 129922 57498 129978
rect 57554 129922 57622 129978
rect 57678 129922 75250 129978
rect 75306 129922 75374 129978
rect 75430 129922 75498 129978
rect 75554 129922 75622 129978
rect 75678 129922 93250 129978
rect 93306 129922 93374 129978
rect 93430 129922 93498 129978
rect 93554 129922 93622 129978
rect 93678 129922 111250 129978
rect 111306 129922 111374 129978
rect 111430 129922 111498 129978
rect 111554 129922 111622 129978
rect 111678 129922 129250 129978
rect 129306 129922 129374 129978
rect 129430 129922 129498 129978
rect 129554 129922 129622 129978
rect 129678 129922 147250 129978
rect 147306 129922 147374 129978
rect 147430 129922 147498 129978
rect 147554 129922 147622 129978
rect 147678 129922 165250 129978
rect 165306 129922 165374 129978
rect 165430 129922 165498 129978
rect 165554 129922 165622 129978
rect 165678 129922 183250 129978
rect 183306 129922 183374 129978
rect 183430 129922 183498 129978
rect 183554 129922 183622 129978
rect 183678 129922 201250 129978
rect 201306 129922 201374 129978
rect 201430 129922 201498 129978
rect 201554 129922 201622 129978
rect 201678 129922 381250 129978
rect 381306 129922 381374 129978
rect 381430 129922 381498 129978
rect 381554 129922 381622 129978
rect 381678 129922 399250 129978
rect 399306 129922 399374 129978
rect 399430 129922 399498 129978
rect 399554 129922 399622 129978
rect 399678 129922 417250 129978
rect 417306 129922 417374 129978
rect 417430 129922 417498 129978
rect 417554 129922 417622 129978
rect 417678 129922 435250 129978
rect 435306 129922 435374 129978
rect 435430 129922 435498 129978
rect 435554 129922 435622 129978
rect 435678 129922 453250 129978
rect 453306 129922 453374 129978
rect 453430 129922 453498 129978
rect 453554 129922 453622 129978
rect 453678 129922 471250 129978
rect 471306 129922 471374 129978
rect 471430 129922 471498 129978
rect 471554 129922 471622 129978
rect 471678 129922 489250 129978
rect 489306 129922 489374 129978
rect 489430 129922 489498 129978
rect 489554 129922 489622 129978
rect 489678 129922 507250 129978
rect 507306 129922 507374 129978
rect 507430 129922 507498 129978
rect 507554 129922 507622 129978
rect 507678 129922 525250 129978
rect 525306 129922 525374 129978
rect 525430 129922 525498 129978
rect 525554 129922 525622 129978
rect 525678 129922 543250 129978
rect 543306 129922 543374 129978
rect 543430 129922 543498 129978
rect 543554 129922 543622 129978
rect 543678 129922 561250 129978
rect 561306 129922 561374 129978
rect 561430 129922 561498 129978
rect 561554 129922 561622 129978
rect 561678 129922 579250 129978
rect 579306 129922 579374 129978
rect 579430 129922 579498 129978
rect 579554 129922 579622 129978
rect 579678 129922 596496 129978
rect 596552 129922 596620 129978
rect 596676 129922 596744 129978
rect 596800 129922 596868 129978
rect 596924 129922 597980 129978
rect -1916 129826 597980 129922
rect -1916 118350 597980 118446
rect -1916 118294 -1820 118350
rect -1764 118294 -1696 118350
rect -1640 118294 -1572 118350
rect -1516 118294 -1448 118350
rect -1392 118294 6970 118350
rect 7026 118294 7094 118350
rect 7150 118294 7218 118350
rect 7274 118294 7342 118350
rect 7398 118294 24970 118350
rect 25026 118294 25094 118350
rect 25150 118294 25218 118350
rect 25274 118294 25342 118350
rect 25398 118294 42970 118350
rect 43026 118294 43094 118350
rect 43150 118294 43218 118350
rect 43274 118294 43342 118350
rect 43398 118294 60970 118350
rect 61026 118294 61094 118350
rect 61150 118294 61218 118350
rect 61274 118294 61342 118350
rect 61398 118294 78970 118350
rect 79026 118294 79094 118350
rect 79150 118294 79218 118350
rect 79274 118294 79342 118350
rect 79398 118294 96970 118350
rect 97026 118294 97094 118350
rect 97150 118294 97218 118350
rect 97274 118294 97342 118350
rect 97398 118294 114970 118350
rect 115026 118294 115094 118350
rect 115150 118294 115218 118350
rect 115274 118294 115342 118350
rect 115398 118294 132970 118350
rect 133026 118294 133094 118350
rect 133150 118294 133218 118350
rect 133274 118294 133342 118350
rect 133398 118294 150970 118350
rect 151026 118294 151094 118350
rect 151150 118294 151218 118350
rect 151274 118294 151342 118350
rect 151398 118294 168970 118350
rect 169026 118294 169094 118350
rect 169150 118294 169218 118350
rect 169274 118294 169342 118350
rect 169398 118294 186970 118350
rect 187026 118294 187094 118350
rect 187150 118294 187218 118350
rect 187274 118294 187342 118350
rect 187398 118294 204970 118350
rect 205026 118294 205094 118350
rect 205150 118294 205218 118350
rect 205274 118294 205342 118350
rect 205398 118294 384970 118350
rect 385026 118294 385094 118350
rect 385150 118294 385218 118350
rect 385274 118294 385342 118350
rect 385398 118294 402970 118350
rect 403026 118294 403094 118350
rect 403150 118294 403218 118350
rect 403274 118294 403342 118350
rect 403398 118294 420970 118350
rect 421026 118294 421094 118350
rect 421150 118294 421218 118350
rect 421274 118294 421342 118350
rect 421398 118294 438970 118350
rect 439026 118294 439094 118350
rect 439150 118294 439218 118350
rect 439274 118294 439342 118350
rect 439398 118294 456970 118350
rect 457026 118294 457094 118350
rect 457150 118294 457218 118350
rect 457274 118294 457342 118350
rect 457398 118294 474970 118350
rect 475026 118294 475094 118350
rect 475150 118294 475218 118350
rect 475274 118294 475342 118350
rect 475398 118294 492970 118350
rect 493026 118294 493094 118350
rect 493150 118294 493218 118350
rect 493274 118294 493342 118350
rect 493398 118294 510970 118350
rect 511026 118294 511094 118350
rect 511150 118294 511218 118350
rect 511274 118294 511342 118350
rect 511398 118294 528970 118350
rect 529026 118294 529094 118350
rect 529150 118294 529218 118350
rect 529274 118294 529342 118350
rect 529398 118294 546970 118350
rect 547026 118294 547094 118350
rect 547150 118294 547218 118350
rect 547274 118294 547342 118350
rect 547398 118294 564970 118350
rect 565026 118294 565094 118350
rect 565150 118294 565218 118350
rect 565274 118294 565342 118350
rect 565398 118294 582970 118350
rect 583026 118294 583094 118350
rect 583150 118294 583218 118350
rect 583274 118294 583342 118350
rect 583398 118294 597456 118350
rect 597512 118294 597580 118350
rect 597636 118294 597704 118350
rect 597760 118294 597828 118350
rect 597884 118294 597980 118350
rect -1916 118226 597980 118294
rect -1916 118170 -1820 118226
rect -1764 118170 -1696 118226
rect -1640 118170 -1572 118226
rect -1516 118170 -1448 118226
rect -1392 118170 6970 118226
rect 7026 118170 7094 118226
rect 7150 118170 7218 118226
rect 7274 118170 7342 118226
rect 7398 118170 24970 118226
rect 25026 118170 25094 118226
rect 25150 118170 25218 118226
rect 25274 118170 25342 118226
rect 25398 118170 42970 118226
rect 43026 118170 43094 118226
rect 43150 118170 43218 118226
rect 43274 118170 43342 118226
rect 43398 118170 60970 118226
rect 61026 118170 61094 118226
rect 61150 118170 61218 118226
rect 61274 118170 61342 118226
rect 61398 118170 78970 118226
rect 79026 118170 79094 118226
rect 79150 118170 79218 118226
rect 79274 118170 79342 118226
rect 79398 118170 96970 118226
rect 97026 118170 97094 118226
rect 97150 118170 97218 118226
rect 97274 118170 97342 118226
rect 97398 118170 114970 118226
rect 115026 118170 115094 118226
rect 115150 118170 115218 118226
rect 115274 118170 115342 118226
rect 115398 118170 132970 118226
rect 133026 118170 133094 118226
rect 133150 118170 133218 118226
rect 133274 118170 133342 118226
rect 133398 118170 150970 118226
rect 151026 118170 151094 118226
rect 151150 118170 151218 118226
rect 151274 118170 151342 118226
rect 151398 118170 168970 118226
rect 169026 118170 169094 118226
rect 169150 118170 169218 118226
rect 169274 118170 169342 118226
rect 169398 118170 186970 118226
rect 187026 118170 187094 118226
rect 187150 118170 187218 118226
rect 187274 118170 187342 118226
rect 187398 118170 204970 118226
rect 205026 118170 205094 118226
rect 205150 118170 205218 118226
rect 205274 118170 205342 118226
rect 205398 118170 384970 118226
rect 385026 118170 385094 118226
rect 385150 118170 385218 118226
rect 385274 118170 385342 118226
rect 385398 118170 402970 118226
rect 403026 118170 403094 118226
rect 403150 118170 403218 118226
rect 403274 118170 403342 118226
rect 403398 118170 420970 118226
rect 421026 118170 421094 118226
rect 421150 118170 421218 118226
rect 421274 118170 421342 118226
rect 421398 118170 438970 118226
rect 439026 118170 439094 118226
rect 439150 118170 439218 118226
rect 439274 118170 439342 118226
rect 439398 118170 456970 118226
rect 457026 118170 457094 118226
rect 457150 118170 457218 118226
rect 457274 118170 457342 118226
rect 457398 118170 474970 118226
rect 475026 118170 475094 118226
rect 475150 118170 475218 118226
rect 475274 118170 475342 118226
rect 475398 118170 492970 118226
rect 493026 118170 493094 118226
rect 493150 118170 493218 118226
rect 493274 118170 493342 118226
rect 493398 118170 510970 118226
rect 511026 118170 511094 118226
rect 511150 118170 511218 118226
rect 511274 118170 511342 118226
rect 511398 118170 528970 118226
rect 529026 118170 529094 118226
rect 529150 118170 529218 118226
rect 529274 118170 529342 118226
rect 529398 118170 546970 118226
rect 547026 118170 547094 118226
rect 547150 118170 547218 118226
rect 547274 118170 547342 118226
rect 547398 118170 564970 118226
rect 565026 118170 565094 118226
rect 565150 118170 565218 118226
rect 565274 118170 565342 118226
rect 565398 118170 582970 118226
rect 583026 118170 583094 118226
rect 583150 118170 583218 118226
rect 583274 118170 583342 118226
rect 583398 118170 597456 118226
rect 597512 118170 597580 118226
rect 597636 118170 597704 118226
rect 597760 118170 597828 118226
rect 597884 118170 597980 118226
rect -1916 118102 597980 118170
rect -1916 118046 -1820 118102
rect -1764 118046 -1696 118102
rect -1640 118046 -1572 118102
rect -1516 118046 -1448 118102
rect -1392 118046 6970 118102
rect 7026 118046 7094 118102
rect 7150 118046 7218 118102
rect 7274 118046 7342 118102
rect 7398 118046 24970 118102
rect 25026 118046 25094 118102
rect 25150 118046 25218 118102
rect 25274 118046 25342 118102
rect 25398 118046 42970 118102
rect 43026 118046 43094 118102
rect 43150 118046 43218 118102
rect 43274 118046 43342 118102
rect 43398 118046 60970 118102
rect 61026 118046 61094 118102
rect 61150 118046 61218 118102
rect 61274 118046 61342 118102
rect 61398 118046 78970 118102
rect 79026 118046 79094 118102
rect 79150 118046 79218 118102
rect 79274 118046 79342 118102
rect 79398 118046 96970 118102
rect 97026 118046 97094 118102
rect 97150 118046 97218 118102
rect 97274 118046 97342 118102
rect 97398 118046 114970 118102
rect 115026 118046 115094 118102
rect 115150 118046 115218 118102
rect 115274 118046 115342 118102
rect 115398 118046 132970 118102
rect 133026 118046 133094 118102
rect 133150 118046 133218 118102
rect 133274 118046 133342 118102
rect 133398 118046 150970 118102
rect 151026 118046 151094 118102
rect 151150 118046 151218 118102
rect 151274 118046 151342 118102
rect 151398 118046 168970 118102
rect 169026 118046 169094 118102
rect 169150 118046 169218 118102
rect 169274 118046 169342 118102
rect 169398 118046 186970 118102
rect 187026 118046 187094 118102
rect 187150 118046 187218 118102
rect 187274 118046 187342 118102
rect 187398 118046 204970 118102
rect 205026 118046 205094 118102
rect 205150 118046 205218 118102
rect 205274 118046 205342 118102
rect 205398 118046 384970 118102
rect 385026 118046 385094 118102
rect 385150 118046 385218 118102
rect 385274 118046 385342 118102
rect 385398 118046 402970 118102
rect 403026 118046 403094 118102
rect 403150 118046 403218 118102
rect 403274 118046 403342 118102
rect 403398 118046 420970 118102
rect 421026 118046 421094 118102
rect 421150 118046 421218 118102
rect 421274 118046 421342 118102
rect 421398 118046 438970 118102
rect 439026 118046 439094 118102
rect 439150 118046 439218 118102
rect 439274 118046 439342 118102
rect 439398 118046 456970 118102
rect 457026 118046 457094 118102
rect 457150 118046 457218 118102
rect 457274 118046 457342 118102
rect 457398 118046 474970 118102
rect 475026 118046 475094 118102
rect 475150 118046 475218 118102
rect 475274 118046 475342 118102
rect 475398 118046 492970 118102
rect 493026 118046 493094 118102
rect 493150 118046 493218 118102
rect 493274 118046 493342 118102
rect 493398 118046 510970 118102
rect 511026 118046 511094 118102
rect 511150 118046 511218 118102
rect 511274 118046 511342 118102
rect 511398 118046 528970 118102
rect 529026 118046 529094 118102
rect 529150 118046 529218 118102
rect 529274 118046 529342 118102
rect 529398 118046 546970 118102
rect 547026 118046 547094 118102
rect 547150 118046 547218 118102
rect 547274 118046 547342 118102
rect 547398 118046 564970 118102
rect 565026 118046 565094 118102
rect 565150 118046 565218 118102
rect 565274 118046 565342 118102
rect 565398 118046 582970 118102
rect 583026 118046 583094 118102
rect 583150 118046 583218 118102
rect 583274 118046 583342 118102
rect 583398 118046 597456 118102
rect 597512 118046 597580 118102
rect 597636 118046 597704 118102
rect 597760 118046 597828 118102
rect 597884 118046 597980 118102
rect -1916 117978 597980 118046
rect -1916 117922 -1820 117978
rect -1764 117922 -1696 117978
rect -1640 117922 -1572 117978
rect -1516 117922 -1448 117978
rect -1392 117922 6970 117978
rect 7026 117922 7094 117978
rect 7150 117922 7218 117978
rect 7274 117922 7342 117978
rect 7398 117922 24970 117978
rect 25026 117922 25094 117978
rect 25150 117922 25218 117978
rect 25274 117922 25342 117978
rect 25398 117922 42970 117978
rect 43026 117922 43094 117978
rect 43150 117922 43218 117978
rect 43274 117922 43342 117978
rect 43398 117922 60970 117978
rect 61026 117922 61094 117978
rect 61150 117922 61218 117978
rect 61274 117922 61342 117978
rect 61398 117922 78970 117978
rect 79026 117922 79094 117978
rect 79150 117922 79218 117978
rect 79274 117922 79342 117978
rect 79398 117922 96970 117978
rect 97026 117922 97094 117978
rect 97150 117922 97218 117978
rect 97274 117922 97342 117978
rect 97398 117922 114970 117978
rect 115026 117922 115094 117978
rect 115150 117922 115218 117978
rect 115274 117922 115342 117978
rect 115398 117922 132970 117978
rect 133026 117922 133094 117978
rect 133150 117922 133218 117978
rect 133274 117922 133342 117978
rect 133398 117922 150970 117978
rect 151026 117922 151094 117978
rect 151150 117922 151218 117978
rect 151274 117922 151342 117978
rect 151398 117922 168970 117978
rect 169026 117922 169094 117978
rect 169150 117922 169218 117978
rect 169274 117922 169342 117978
rect 169398 117922 186970 117978
rect 187026 117922 187094 117978
rect 187150 117922 187218 117978
rect 187274 117922 187342 117978
rect 187398 117922 204970 117978
rect 205026 117922 205094 117978
rect 205150 117922 205218 117978
rect 205274 117922 205342 117978
rect 205398 117922 384970 117978
rect 385026 117922 385094 117978
rect 385150 117922 385218 117978
rect 385274 117922 385342 117978
rect 385398 117922 402970 117978
rect 403026 117922 403094 117978
rect 403150 117922 403218 117978
rect 403274 117922 403342 117978
rect 403398 117922 420970 117978
rect 421026 117922 421094 117978
rect 421150 117922 421218 117978
rect 421274 117922 421342 117978
rect 421398 117922 438970 117978
rect 439026 117922 439094 117978
rect 439150 117922 439218 117978
rect 439274 117922 439342 117978
rect 439398 117922 456970 117978
rect 457026 117922 457094 117978
rect 457150 117922 457218 117978
rect 457274 117922 457342 117978
rect 457398 117922 474970 117978
rect 475026 117922 475094 117978
rect 475150 117922 475218 117978
rect 475274 117922 475342 117978
rect 475398 117922 492970 117978
rect 493026 117922 493094 117978
rect 493150 117922 493218 117978
rect 493274 117922 493342 117978
rect 493398 117922 510970 117978
rect 511026 117922 511094 117978
rect 511150 117922 511218 117978
rect 511274 117922 511342 117978
rect 511398 117922 528970 117978
rect 529026 117922 529094 117978
rect 529150 117922 529218 117978
rect 529274 117922 529342 117978
rect 529398 117922 546970 117978
rect 547026 117922 547094 117978
rect 547150 117922 547218 117978
rect 547274 117922 547342 117978
rect 547398 117922 564970 117978
rect 565026 117922 565094 117978
rect 565150 117922 565218 117978
rect 565274 117922 565342 117978
rect 565398 117922 582970 117978
rect 583026 117922 583094 117978
rect 583150 117922 583218 117978
rect 583274 117922 583342 117978
rect 583398 117922 597456 117978
rect 597512 117922 597580 117978
rect 597636 117922 597704 117978
rect 597760 117922 597828 117978
rect 597884 117922 597980 117978
rect -1916 117826 597980 117922
rect -1916 112350 597980 112446
rect -1916 112294 -860 112350
rect -804 112294 -736 112350
rect -680 112294 -612 112350
rect -556 112294 -488 112350
rect -432 112294 3250 112350
rect 3306 112294 3374 112350
rect 3430 112294 3498 112350
rect 3554 112294 3622 112350
rect 3678 112294 21250 112350
rect 21306 112294 21374 112350
rect 21430 112294 21498 112350
rect 21554 112294 21622 112350
rect 21678 112294 39250 112350
rect 39306 112294 39374 112350
rect 39430 112294 39498 112350
rect 39554 112294 39622 112350
rect 39678 112294 57250 112350
rect 57306 112294 57374 112350
rect 57430 112294 57498 112350
rect 57554 112294 57622 112350
rect 57678 112294 75250 112350
rect 75306 112294 75374 112350
rect 75430 112294 75498 112350
rect 75554 112294 75622 112350
rect 75678 112294 93250 112350
rect 93306 112294 93374 112350
rect 93430 112294 93498 112350
rect 93554 112294 93622 112350
rect 93678 112294 111250 112350
rect 111306 112294 111374 112350
rect 111430 112294 111498 112350
rect 111554 112294 111622 112350
rect 111678 112294 129250 112350
rect 129306 112294 129374 112350
rect 129430 112294 129498 112350
rect 129554 112294 129622 112350
rect 129678 112294 147250 112350
rect 147306 112294 147374 112350
rect 147430 112294 147498 112350
rect 147554 112294 147622 112350
rect 147678 112294 165250 112350
rect 165306 112294 165374 112350
rect 165430 112294 165498 112350
rect 165554 112294 165622 112350
rect 165678 112294 183250 112350
rect 183306 112294 183374 112350
rect 183430 112294 183498 112350
rect 183554 112294 183622 112350
rect 183678 112294 201250 112350
rect 201306 112294 201374 112350
rect 201430 112294 201498 112350
rect 201554 112294 201622 112350
rect 201678 112294 381250 112350
rect 381306 112294 381374 112350
rect 381430 112294 381498 112350
rect 381554 112294 381622 112350
rect 381678 112294 399250 112350
rect 399306 112294 399374 112350
rect 399430 112294 399498 112350
rect 399554 112294 399622 112350
rect 399678 112294 417250 112350
rect 417306 112294 417374 112350
rect 417430 112294 417498 112350
rect 417554 112294 417622 112350
rect 417678 112294 435250 112350
rect 435306 112294 435374 112350
rect 435430 112294 435498 112350
rect 435554 112294 435622 112350
rect 435678 112294 453250 112350
rect 453306 112294 453374 112350
rect 453430 112294 453498 112350
rect 453554 112294 453622 112350
rect 453678 112294 471250 112350
rect 471306 112294 471374 112350
rect 471430 112294 471498 112350
rect 471554 112294 471622 112350
rect 471678 112294 489250 112350
rect 489306 112294 489374 112350
rect 489430 112294 489498 112350
rect 489554 112294 489622 112350
rect 489678 112294 507250 112350
rect 507306 112294 507374 112350
rect 507430 112294 507498 112350
rect 507554 112294 507622 112350
rect 507678 112294 525250 112350
rect 525306 112294 525374 112350
rect 525430 112294 525498 112350
rect 525554 112294 525622 112350
rect 525678 112294 543250 112350
rect 543306 112294 543374 112350
rect 543430 112294 543498 112350
rect 543554 112294 543622 112350
rect 543678 112294 561250 112350
rect 561306 112294 561374 112350
rect 561430 112294 561498 112350
rect 561554 112294 561622 112350
rect 561678 112294 579250 112350
rect 579306 112294 579374 112350
rect 579430 112294 579498 112350
rect 579554 112294 579622 112350
rect 579678 112294 596496 112350
rect 596552 112294 596620 112350
rect 596676 112294 596744 112350
rect 596800 112294 596868 112350
rect 596924 112294 597980 112350
rect -1916 112226 597980 112294
rect -1916 112170 -860 112226
rect -804 112170 -736 112226
rect -680 112170 -612 112226
rect -556 112170 -488 112226
rect -432 112170 3250 112226
rect 3306 112170 3374 112226
rect 3430 112170 3498 112226
rect 3554 112170 3622 112226
rect 3678 112170 21250 112226
rect 21306 112170 21374 112226
rect 21430 112170 21498 112226
rect 21554 112170 21622 112226
rect 21678 112170 39250 112226
rect 39306 112170 39374 112226
rect 39430 112170 39498 112226
rect 39554 112170 39622 112226
rect 39678 112170 57250 112226
rect 57306 112170 57374 112226
rect 57430 112170 57498 112226
rect 57554 112170 57622 112226
rect 57678 112170 75250 112226
rect 75306 112170 75374 112226
rect 75430 112170 75498 112226
rect 75554 112170 75622 112226
rect 75678 112170 93250 112226
rect 93306 112170 93374 112226
rect 93430 112170 93498 112226
rect 93554 112170 93622 112226
rect 93678 112170 111250 112226
rect 111306 112170 111374 112226
rect 111430 112170 111498 112226
rect 111554 112170 111622 112226
rect 111678 112170 129250 112226
rect 129306 112170 129374 112226
rect 129430 112170 129498 112226
rect 129554 112170 129622 112226
rect 129678 112170 147250 112226
rect 147306 112170 147374 112226
rect 147430 112170 147498 112226
rect 147554 112170 147622 112226
rect 147678 112170 165250 112226
rect 165306 112170 165374 112226
rect 165430 112170 165498 112226
rect 165554 112170 165622 112226
rect 165678 112170 183250 112226
rect 183306 112170 183374 112226
rect 183430 112170 183498 112226
rect 183554 112170 183622 112226
rect 183678 112170 201250 112226
rect 201306 112170 201374 112226
rect 201430 112170 201498 112226
rect 201554 112170 201622 112226
rect 201678 112170 381250 112226
rect 381306 112170 381374 112226
rect 381430 112170 381498 112226
rect 381554 112170 381622 112226
rect 381678 112170 399250 112226
rect 399306 112170 399374 112226
rect 399430 112170 399498 112226
rect 399554 112170 399622 112226
rect 399678 112170 417250 112226
rect 417306 112170 417374 112226
rect 417430 112170 417498 112226
rect 417554 112170 417622 112226
rect 417678 112170 435250 112226
rect 435306 112170 435374 112226
rect 435430 112170 435498 112226
rect 435554 112170 435622 112226
rect 435678 112170 453250 112226
rect 453306 112170 453374 112226
rect 453430 112170 453498 112226
rect 453554 112170 453622 112226
rect 453678 112170 471250 112226
rect 471306 112170 471374 112226
rect 471430 112170 471498 112226
rect 471554 112170 471622 112226
rect 471678 112170 489250 112226
rect 489306 112170 489374 112226
rect 489430 112170 489498 112226
rect 489554 112170 489622 112226
rect 489678 112170 507250 112226
rect 507306 112170 507374 112226
rect 507430 112170 507498 112226
rect 507554 112170 507622 112226
rect 507678 112170 525250 112226
rect 525306 112170 525374 112226
rect 525430 112170 525498 112226
rect 525554 112170 525622 112226
rect 525678 112170 543250 112226
rect 543306 112170 543374 112226
rect 543430 112170 543498 112226
rect 543554 112170 543622 112226
rect 543678 112170 561250 112226
rect 561306 112170 561374 112226
rect 561430 112170 561498 112226
rect 561554 112170 561622 112226
rect 561678 112170 579250 112226
rect 579306 112170 579374 112226
rect 579430 112170 579498 112226
rect 579554 112170 579622 112226
rect 579678 112170 596496 112226
rect 596552 112170 596620 112226
rect 596676 112170 596744 112226
rect 596800 112170 596868 112226
rect 596924 112170 597980 112226
rect -1916 112102 597980 112170
rect -1916 112046 -860 112102
rect -804 112046 -736 112102
rect -680 112046 -612 112102
rect -556 112046 -488 112102
rect -432 112046 3250 112102
rect 3306 112046 3374 112102
rect 3430 112046 3498 112102
rect 3554 112046 3622 112102
rect 3678 112046 21250 112102
rect 21306 112046 21374 112102
rect 21430 112046 21498 112102
rect 21554 112046 21622 112102
rect 21678 112046 39250 112102
rect 39306 112046 39374 112102
rect 39430 112046 39498 112102
rect 39554 112046 39622 112102
rect 39678 112046 57250 112102
rect 57306 112046 57374 112102
rect 57430 112046 57498 112102
rect 57554 112046 57622 112102
rect 57678 112046 75250 112102
rect 75306 112046 75374 112102
rect 75430 112046 75498 112102
rect 75554 112046 75622 112102
rect 75678 112046 93250 112102
rect 93306 112046 93374 112102
rect 93430 112046 93498 112102
rect 93554 112046 93622 112102
rect 93678 112046 111250 112102
rect 111306 112046 111374 112102
rect 111430 112046 111498 112102
rect 111554 112046 111622 112102
rect 111678 112046 129250 112102
rect 129306 112046 129374 112102
rect 129430 112046 129498 112102
rect 129554 112046 129622 112102
rect 129678 112046 147250 112102
rect 147306 112046 147374 112102
rect 147430 112046 147498 112102
rect 147554 112046 147622 112102
rect 147678 112046 165250 112102
rect 165306 112046 165374 112102
rect 165430 112046 165498 112102
rect 165554 112046 165622 112102
rect 165678 112046 183250 112102
rect 183306 112046 183374 112102
rect 183430 112046 183498 112102
rect 183554 112046 183622 112102
rect 183678 112046 201250 112102
rect 201306 112046 201374 112102
rect 201430 112046 201498 112102
rect 201554 112046 201622 112102
rect 201678 112046 381250 112102
rect 381306 112046 381374 112102
rect 381430 112046 381498 112102
rect 381554 112046 381622 112102
rect 381678 112046 399250 112102
rect 399306 112046 399374 112102
rect 399430 112046 399498 112102
rect 399554 112046 399622 112102
rect 399678 112046 417250 112102
rect 417306 112046 417374 112102
rect 417430 112046 417498 112102
rect 417554 112046 417622 112102
rect 417678 112046 435250 112102
rect 435306 112046 435374 112102
rect 435430 112046 435498 112102
rect 435554 112046 435622 112102
rect 435678 112046 453250 112102
rect 453306 112046 453374 112102
rect 453430 112046 453498 112102
rect 453554 112046 453622 112102
rect 453678 112046 471250 112102
rect 471306 112046 471374 112102
rect 471430 112046 471498 112102
rect 471554 112046 471622 112102
rect 471678 112046 489250 112102
rect 489306 112046 489374 112102
rect 489430 112046 489498 112102
rect 489554 112046 489622 112102
rect 489678 112046 507250 112102
rect 507306 112046 507374 112102
rect 507430 112046 507498 112102
rect 507554 112046 507622 112102
rect 507678 112046 525250 112102
rect 525306 112046 525374 112102
rect 525430 112046 525498 112102
rect 525554 112046 525622 112102
rect 525678 112046 543250 112102
rect 543306 112046 543374 112102
rect 543430 112046 543498 112102
rect 543554 112046 543622 112102
rect 543678 112046 561250 112102
rect 561306 112046 561374 112102
rect 561430 112046 561498 112102
rect 561554 112046 561622 112102
rect 561678 112046 579250 112102
rect 579306 112046 579374 112102
rect 579430 112046 579498 112102
rect 579554 112046 579622 112102
rect 579678 112046 596496 112102
rect 596552 112046 596620 112102
rect 596676 112046 596744 112102
rect 596800 112046 596868 112102
rect 596924 112046 597980 112102
rect -1916 111978 597980 112046
rect -1916 111922 -860 111978
rect -804 111922 -736 111978
rect -680 111922 -612 111978
rect -556 111922 -488 111978
rect -432 111922 3250 111978
rect 3306 111922 3374 111978
rect 3430 111922 3498 111978
rect 3554 111922 3622 111978
rect 3678 111922 21250 111978
rect 21306 111922 21374 111978
rect 21430 111922 21498 111978
rect 21554 111922 21622 111978
rect 21678 111922 39250 111978
rect 39306 111922 39374 111978
rect 39430 111922 39498 111978
rect 39554 111922 39622 111978
rect 39678 111922 57250 111978
rect 57306 111922 57374 111978
rect 57430 111922 57498 111978
rect 57554 111922 57622 111978
rect 57678 111922 75250 111978
rect 75306 111922 75374 111978
rect 75430 111922 75498 111978
rect 75554 111922 75622 111978
rect 75678 111922 93250 111978
rect 93306 111922 93374 111978
rect 93430 111922 93498 111978
rect 93554 111922 93622 111978
rect 93678 111922 111250 111978
rect 111306 111922 111374 111978
rect 111430 111922 111498 111978
rect 111554 111922 111622 111978
rect 111678 111922 129250 111978
rect 129306 111922 129374 111978
rect 129430 111922 129498 111978
rect 129554 111922 129622 111978
rect 129678 111922 147250 111978
rect 147306 111922 147374 111978
rect 147430 111922 147498 111978
rect 147554 111922 147622 111978
rect 147678 111922 165250 111978
rect 165306 111922 165374 111978
rect 165430 111922 165498 111978
rect 165554 111922 165622 111978
rect 165678 111922 183250 111978
rect 183306 111922 183374 111978
rect 183430 111922 183498 111978
rect 183554 111922 183622 111978
rect 183678 111922 201250 111978
rect 201306 111922 201374 111978
rect 201430 111922 201498 111978
rect 201554 111922 201622 111978
rect 201678 111922 381250 111978
rect 381306 111922 381374 111978
rect 381430 111922 381498 111978
rect 381554 111922 381622 111978
rect 381678 111922 399250 111978
rect 399306 111922 399374 111978
rect 399430 111922 399498 111978
rect 399554 111922 399622 111978
rect 399678 111922 417250 111978
rect 417306 111922 417374 111978
rect 417430 111922 417498 111978
rect 417554 111922 417622 111978
rect 417678 111922 435250 111978
rect 435306 111922 435374 111978
rect 435430 111922 435498 111978
rect 435554 111922 435622 111978
rect 435678 111922 453250 111978
rect 453306 111922 453374 111978
rect 453430 111922 453498 111978
rect 453554 111922 453622 111978
rect 453678 111922 471250 111978
rect 471306 111922 471374 111978
rect 471430 111922 471498 111978
rect 471554 111922 471622 111978
rect 471678 111922 489250 111978
rect 489306 111922 489374 111978
rect 489430 111922 489498 111978
rect 489554 111922 489622 111978
rect 489678 111922 507250 111978
rect 507306 111922 507374 111978
rect 507430 111922 507498 111978
rect 507554 111922 507622 111978
rect 507678 111922 525250 111978
rect 525306 111922 525374 111978
rect 525430 111922 525498 111978
rect 525554 111922 525622 111978
rect 525678 111922 543250 111978
rect 543306 111922 543374 111978
rect 543430 111922 543498 111978
rect 543554 111922 543622 111978
rect 543678 111922 561250 111978
rect 561306 111922 561374 111978
rect 561430 111922 561498 111978
rect 561554 111922 561622 111978
rect 561678 111922 579250 111978
rect 579306 111922 579374 111978
rect 579430 111922 579498 111978
rect 579554 111922 579622 111978
rect 579678 111922 596496 111978
rect 596552 111922 596620 111978
rect 596676 111922 596744 111978
rect 596800 111922 596868 111978
rect 596924 111922 597980 111978
rect -1916 111826 597980 111922
rect -1916 100350 597980 100446
rect -1916 100294 -1820 100350
rect -1764 100294 -1696 100350
rect -1640 100294 -1572 100350
rect -1516 100294 -1448 100350
rect -1392 100294 6970 100350
rect 7026 100294 7094 100350
rect 7150 100294 7218 100350
rect 7274 100294 7342 100350
rect 7398 100294 24970 100350
rect 25026 100294 25094 100350
rect 25150 100294 25218 100350
rect 25274 100294 25342 100350
rect 25398 100294 42970 100350
rect 43026 100294 43094 100350
rect 43150 100294 43218 100350
rect 43274 100294 43342 100350
rect 43398 100294 186970 100350
rect 187026 100294 187094 100350
rect 187150 100294 187218 100350
rect 187274 100294 187342 100350
rect 187398 100294 204970 100350
rect 205026 100294 205094 100350
rect 205150 100294 205218 100350
rect 205274 100294 205342 100350
rect 205398 100294 384970 100350
rect 385026 100294 385094 100350
rect 385150 100294 385218 100350
rect 385274 100294 385342 100350
rect 385398 100294 402970 100350
rect 403026 100294 403094 100350
rect 403150 100294 403218 100350
rect 403274 100294 403342 100350
rect 403398 100294 420970 100350
rect 421026 100294 421094 100350
rect 421150 100294 421218 100350
rect 421274 100294 421342 100350
rect 421398 100294 438970 100350
rect 439026 100294 439094 100350
rect 439150 100294 439218 100350
rect 439274 100294 439342 100350
rect 439398 100294 456970 100350
rect 457026 100294 457094 100350
rect 457150 100294 457218 100350
rect 457274 100294 457342 100350
rect 457398 100294 474970 100350
rect 475026 100294 475094 100350
rect 475150 100294 475218 100350
rect 475274 100294 475342 100350
rect 475398 100294 492970 100350
rect 493026 100294 493094 100350
rect 493150 100294 493218 100350
rect 493274 100294 493342 100350
rect 493398 100294 510970 100350
rect 511026 100294 511094 100350
rect 511150 100294 511218 100350
rect 511274 100294 511342 100350
rect 511398 100294 528970 100350
rect 529026 100294 529094 100350
rect 529150 100294 529218 100350
rect 529274 100294 529342 100350
rect 529398 100294 539878 100350
rect 539934 100294 540002 100350
rect 540058 100294 546970 100350
rect 547026 100294 547094 100350
rect 547150 100294 547218 100350
rect 547274 100294 547342 100350
rect 547398 100294 564970 100350
rect 565026 100294 565094 100350
rect 565150 100294 565218 100350
rect 565274 100294 565342 100350
rect 565398 100294 582970 100350
rect 583026 100294 583094 100350
rect 583150 100294 583218 100350
rect 583274 100294 583342 100350
rect 583398 100294 597456 100350
rect 597512 100294 597580 100350
rect 597636 100294 597704 100350
rect 597760 100294 597828 100350
rect 597884 100294 597980 100350
rect -1916 100226 597980 100294
rect -1916 100170 -1820 100226
rect -1764 100170 -1696 100226
rect -1640 100170 -1572 100226
rect -1516 100170 -1448 100226
rect -1392 100170 6970 100226
rect 7026 100170 7094 100226
rect 7150 100170 7218 100226
rect 7274 100170 7342 100226
rect 7398 100170 24970 100226
rect 25026 100170 25094 100226
rect 25150 100170 25218 100226
rect 25274 100170 25342 100226
rect 25398 100170 42970 100226
rect 43026 100170 43094 100226
rect 43150 100170 43218 100226
rect 43274 100170 43342 100226
rect 43398 100170 186970 100226
rect 187026 100170 187094 100226
rect 187150 100170 187218 100226
rect 187274 100170 187342 100226
rect 187398 100170 204970 100226
rect 205026 100170 205094 100226
rect 205150 100170 205218 100226
rect 205274 100170 205342 100226
rect 205398 100170 384970 100226
rect 385026 100170 385094 100226
rect 385150 100170 385218 100226
rect 385274 100170 385342 100226
rect 385398 100170 402970 100226
rect 403026 100170 403094 100226
rect 403150 100170 403218 100226
rect 403274 100170 403342 100226
rect 403398 100170 420970 100226
rect 421026 100170 421094 100226
rect 421150 100170 421218 100226
rect 421274 100170 421342 100226
rect 421398 100170 438970 100226
rect 439026 100170 439094 100226
rect 439150 100170 439218 100226
rect 439274 100170 439342 100226
rect 439398 100170 456970 100226
rect 457026 100170 457094 100226
rect 457150 100170 457218 100226
rect 457274 100170 457342 100226
rect 457398 100170 474970 100226
rect 475026 100170 475094 100226
rect 475150 100170 475218 100226
rect 475274 100170 475342 100226
rect 475398 100170 492970 100226
rect 493026 100170 493094 100226
rect 493150 100170 493218 100226
rect 493274 100170 493342 100226
rect 493398 100170 510970 100226
rect 511026 100170 511094 100226
rect 511150 100170 511218 100226
rect 511274 100170 511342 100226
rect 511398 100170 528970 100226
rect 529026 100170 529094 100226
rect 529150 100170 529218 100226
rect 529274 100170 529342 100226
rect 529398 100170 539878 100226
rect 539934 100170 540002 100226
rect 540058 100170 546970 100226
rect 547026 100170 547094 100226
rect 547150 100170 547218 100226
rect 547274 100170 547342 100226
rect 547398 100170 564970 100226
rect 565026 100170 565094 100226
rect 565150 100170 565218 100226
rect 565274 100170 565342 100226
rect 565398 100170 582970 100226
rect 583026 100170 583094 100226
rect 583150 100170 583218 100226
rect 583274 100170 583342 100226
rect 583398 100170 597456 100226
rect 597512 100170 597580 100226
rect 597636 100170 597704 100226
rect 597760 100170 597828 100226
rect 597884 100170 597980 100226
rect -1916 100102 597980 100170
rect -1916 100046 -1820 100102
rect -1764 100046 -1696 100102
rect -1640 100046 -1572 100102
rect -1516 100046 -1448 100102
rect -1392 100046 6970 100102
rect 7026 100046 7094 100102
rect 7150 100046 7218 100102
rect 7274 100046 7342 100102
rect 7398 100046 24970 100102
rect 25026 100046 25094 100102
rect 25150 100046 25218 100102
rect 25274 100046 25342 100102
rect 25398 100046 42970 100102
rect 43026 100046 43094 100102
rect 43150 100046 43218 100102
rect 43274 100046 43342 100102
rect 43398 100046 186970 100102
rect 187026 100046 187094 100102
rect 187150 100046 187218 100102
rect 187274 100046 187342 100102
rect 187398 100046 204970 100102
rect 205026 100046 205094 100102
rect 205150 100046 205218 100102
rect 205274 100046 205342 100102
rect 205398 100046 384970 100102
rect 385026 100046 385094 100102
rect 385150 100046 385218 100102
rect 385274 100046 385342 100102
rect 385398 100046 402970 100102
rect 403026 100046 403094 100102
rect 403150 100046 403218 100102
rect 403274 100046 403342 100102
rect 403398 100046 420970 100102
rect 421026 100046 421094 100102
rect 421150 100046 421218 100102
rect 421274 100046 421342 100102
rect 421398 100046 438970 100102
rect 439026 100046 439094 100102
rect 439150 100046 439218 100102
rect 439274 100046 439342 100102
rect 439398 100046 456970 100102
rect 457026 100046 457094 100102
rect 457150 100046 457218 100102
rect 457274 100046 457342 100102
rect 457398 100046 474970 100102
rect 475026 100046 475094 100102
rect 475150 100046 475218 100102
rect 475274 100046 475342 100102
rect 475398 100046 492970 100102
rect 493026 100046 493094 100102
rect 493150 100046 493218 100102
rect 493274 100046 493342 100102
rect 493398 100046 510970 100102
rect 511026 100046 511094 100102
rect 511150 100046 511218 100102
rect 511274 100046 511342 100102
rect 511398 100046 528970 100102
rect 529026 100046 529094 100102
rect 529150 100046 529218 100102
rect 529274 100046 529342 100102
rect 529398 100046 539878 100102
rect 539934 100046 540002 100102
rect 540058 100046 546970 100102
rect 547026 100046 547094 100102
rect 547150 100046 547218 100102
rect 547274 100046 547342 100102
rect 547398 100046 564970 100102
rect 565026 100046 565094 100102
rect 565150 100046 565218 100102
rect 565274 100046 565342 100102
rect 565398 100046 582970 100102
rect 583026 100046 583094 100102
rect 583150 100046 583218 100102
rect 583274 100046 583342 100102
rect 583398 100046 597456 100102
rect 597512 100046 597580 100102
rect 597636 100046 597704 100102
rect 597760 100046 597828 100102
rect 597884 100046 597980 100102
rect -1916 99978 597980 100046
rect -1916 99922 -1820 99978
rect -1764 99922 -1696 99978
rect -1640 99922 -1572 99978
rect -1516 99922 -1448 99978
rect -1392 99922 6970 99978
rect 7026 99922 7094 99978
rect 7150 99922 7218 99978
rect 7274 99922 7342 99978
rect 7398 99922 24970 99978
rect 25026 99922 25094 99978
rect 25150 99922 25218 99978
rect 25274 99922 25342 99978
rect 25398 99922 42970 99978
rect 43026 99922 43094 99978
rect 43150 99922 43218 99978
rect 43274 99922 43342 99978
rect 43398 99922 186970 99978
rect 187026 99922 187094 99978
rect 187150 99922 187218 99978
rect 187274 99922 187342 99978
rect 187398 99922 204970 99978
rect 205026 99922 205094 99978
rect 205150 99922 205218 99978
rect 205274 99922 205342 99978
rect 205398 99922 384970 99978
rect 385026 99922 385094 99978
rect 385150 99922 385218 99978
rect 385274 99922 385342 99978
rect 385398 99922 402970 99978
rect 403026 99922 403094 99978
rect 403150 99922 403218 99978
rect 403274 99922 403342 99978
rect 403398 99922 420970 99978
rect 421026 99922 421094 99978
rect 421150 99922 421218 99978
rect 421274 99922 421342 99978
rect 421398 99922 438970 99978
rect 439026 99922 439094 99978
rect 439150 99922 439218 99978
rect 439274 99922 439342 99978
rect 439398 99922 456970 99978
rect 457026 99922 457094 99978
rect 457150 99922 457218 99978
rect 457274 99922 457342 99978
rect 457398 99922 474970 99978
rect 475026 99922 475094 99978
rect 475150 99922 475218 99978
rect 475274 99922 475342 99978
rect 475398 99922 492970 99978
rect 493026 99922 493094 99978
rect 493150 99922 493218 99978
rect 493274 99922 493342 99978
rect 493398 99922 510970 99978
rect 511026 99922 511094 99978
rect 511150 99922 511218 99978
rect 511274 99922 511342 99978
rect 511398 99922 528970 99978
rect 529026 99922 529094 99978
rect 529150 99922 529218 99978
rect 529274 99922 529342 99978
rect 529398 99922 539878 99978
rect 539934 99922 540002 99978
rect 540058 99922 546970 99978
rect 547026 99922 547094 99978
rect 547150 99922 547218 99978
rect 547274 99922 547342 99978
rect 547398 99922 564970 99978
rect 565026 99922 565094 99978
rect 565150 99922 565218 99978
rect 565274 99922 565342 99978
rect 565398 99922 582970 99978
rect 583026 99922 583094 99978
rect 583150 99922 583218 99978
rect 583274 99922 583342 99978
rect 583398 99922 597456 99978
rect 597512 99922 597580 99978
rect 597636 99922 597704 99978
rect 597760 99922 597828 99978
rect 597884 99922 597980 99978
rect -1916 99826 597980 99922
rect -1916 94350 597980 94446
rect -1916 94294 -860 94350
rect -804 94294 -736 94350
rect -680 94294 -612 94350
rect -556 94294 -488 94350
rect -432 94294 3250 94350
rect 3306 94294 3374 94350
rect 3430 94294 3498 94350
rect 3554 94294 3622 94350
rect 3678 94294 21250 94350
rect 21306 94294 21374 94350
rect 21430 94294 21498 94350
rect 21554 94294 21622 94350
rect 21678 94294 39250 94350
rect 39306 94294 39374 94350
rect 39430 94294 39498 94350
rect 39554 94294 39622 94350
rect 39678 94294 183250 94350
rect 183306 94294 183374 94350
rect 183430 94294 183498 94350
rect 183554 94294 183622 94350
rect 183678 94294 201250 94350
rect 201306 94294 201374 94350
rect 201430 94294 201498 94350
rect 201554 94294 201622 94350
rect 201678 94294 381250 94350
rect 381306 94294 381374 94350
rect 381430 94294 381498 94350
rect 381554 94294 381622 94350
rect 381678 94294 399250 94350
rect 399306 94294 399374 94350
rect 399430 94294 399498 94350
rect 399554 94294 399622 94350
rect 399678 94294 417250 94350
rect 417306 94294 417374 94350
rect 417430 94294 417498 94350
rect 417554 94294 417622 94350
rect 417678 94294 435250 94350
rect 435306 94294 435374 94350
rect 435430 94294 435498 94350
rect 435554 94294 435622 94350
rect 435678 94294 453250 94350
rect 453306 94294 453374 94350
rect 453430 94294 453498 94350
rect 453554 94294 453622 94350
rect 453678 94294 471250 94350
rect 471306 94294 471374 94350
rect 471430 94294 471498 94350
rect 471554 94294 471622 94350
rect 471678 94294 489250 94350
rect 489306 94294 489374 94350
rect 489430 94294 489498 94350
rect 489554 94294 489622 94350
rect 489678 94294 507250 94350
rect 507306 94294 507374 94350
rect 507430 94294 507498 94350
rect 507554 94294 507622 94350
rect 507678 94294 524518 94350
rect 524574 94294 524642 94350
rect 524698 94294 525250 94350
rect 525306 94294 525374 94350
rect 525430 94294 525498 94350
rect 525554 94294 525622 94350
rect 525678 94294 543250 94350
rect 543306 94294 543374 94350
rect 543430 94294 543498 94350
rect 543554 94294 543622 94350
rect 543678 94294 555238 94350
rect 555294 94294 555362 94350
rect 555418 94294 561250 94350
rect 561306 94294 561374 94350
rect 561430 94294 561498 94350
rect 561554 94294 561622 94350
rect 561678 94294 579250 94350
rect 579306 94294 579374 94350
rect 579430 94294 579498 94350
rect 579554 94294 579622 94350
rect 579678 94294 596496 94350
rect 596552 94294 596620 94350
rect 596676 94294 596744 94350
rect 596800 94294 596868 94350
rect 596924 94294 597980 94350
rect -1916 94226 597980 94294
rect -1916 94170 -860 94226
rect -804 94170 -736 94226
rect -680 94170 -612 94226
rect -556 94170 -488 94226
rect -432 94170 3250 94226
rect 3306 94170 3374 94226
rect 3430 94170 3498 94226
rect 3554 94170 3622 94226
rect 3678 94170 21250 94226
rect 21306 94170 21374 94226
rect 21430 94170 21498 94226
rect 21554 94170 21622 94226
rect 21678 94170 39250 94226
rect 39306 94170 39374 94226
rect 39430 94170 39498 94226
rect 39554 94170 39622 94226
rect 39678 94170 183250 94226
rect 183306 94170 183374 94226
rect 183430 94170 183498 94226
rect 183554 94170 183622 94226
rect 183678 94170 201250 94226
rect 201306 94170 201374 94226
rect 201430 94170 201498 94226
rect 201554 94170 201622 94226
rect 201678 94170 381250 94226
rect 381306 94170 381374 94226
rect 381430 94170 381498 94226
rect 381554 94170 381622 94226
rect 381678 94170 399250 94226
rect 399306 94170 399374 94226
rect 399430 94170 399498 94226
rect 399554 94170 399622 94226
rect 399678 94170 417250 94226
rect 417306 94170 417374 94226
rect 417430 94170 417498 94226
rect 417554 94170 417622 94226
rect 417678 94170 435250 94226
rect 435306 94170 435374 94226
rect 435430 94170 435498 94226
rect 435554 94170 435622 94226
rect 435678 94170 453250 94226
rect 453306 94170 453374 94226
rect 453430 94170 453498 94226
rect 453554 94170 453622 94226
rect 453678 94170 471250 94226
rect 471306 94170 471374 94226
rect 471430 94170 471498 94226
rect 471554 94170 471622 94226
rect 471678 94170 489250 94226
rect 489306 94170 489374 94226
rect 489430 94170 489498 94226
rect 489554 94170 489622 94226
rect 489678 94170 507250 94226
rect 507306 94170 507374 94226
rect 507430 94170 507498 94226
rect 507554 94170 507622 94226
rect 507678 94170 524518 94226
rect 524574 94170 524642 94226
rect 524698 94170 525250 94226
rect 525306 94170 525374 94226
rect 525430 94170 525498 94226
rect 525554 94170 525622 94226
rect 525678 94170 543250 94226
rect 543306 94170 543374 94226
rect 543430 94170 543498 94226
rect 543554 94170 543622 94226
rect 543678 94170 555238 94226
rect 555294 94170 555362 94226
rect 555418 94170 561250 94226
rect 561306 94170 561374 94226
rect 561430 94170 561498 94226
rect 561554 94170 561622 94226
rect 561678 94170 579250 94226
rect 579306 94170 579374 94226
rect 579430 94170 579498 94226
rect 579554 94170 579622 94226
rect 579678 94170 596496 94226
rect 596552 94170 596620 94226
rect 596676 94170 596744 94226
rect 596800 94170 596868 94226
rect 596924 94170 597980 94226
rect -1916 94102 597980 94170
rect -1916 94046 -860 94102
rect -804 94046 -736 94102
rect -680 94046 -612 94102
rect -556 94046 -488 94102
rect -432 94046 3250 94102
rect 3306 94046 3374 94102
rect 3430 94046 3498 94102
rect 3554 94046 3622 94102
rect 3678 94046 21250 94102
rect 21306 94046 21374 94102
rect 21430 94046 21498 94102
rect 21554 94046 21622 94102
rect 21678 94046 39250 94102
rect 39306 94046 39374 94102
rect 39430 94046 39498 94102
rect 39554 94046 39622 94102
rect 39678 94046 183250 94102
rect 183306 94046 183374 94102
rect 183430 94046 183498 94102
rect 183554 94046 183622 94102
rect 183678 94046 201250 94102
rect 201306 94046 201374 94102
rect 201430 94046 201498 94102
rect 201554 94046 201622 94102
rect 201678 94046 381250 94102
rect 381306 94046 381374 94102
rect 381430 94046 381498 94102
rect 381554 94046 381622 94102
rect 381678 94046 399250 94102
rect 399306 94046 399374 94102
rect 399430 94046 399498 94102
rect 399554 94046 399622 94102
rect 399678 94046 417250 94102
rect 417306 94046 417374 94102
rect 417430 94046 417498 94102
rect 417554 94046 417622 94102
rect 417678 94046 435250 94102
rect 435306 94046 435374 94102
rect 435430 94046 435498 94102
rect 435554 94046 435622 94102
rect 435678 94046 453250 94102
rect 453306 94046 453374 94102
rect 453430 94046 453498 94102
rect 453554 94046 453622 94102
rect 453678 94046 471250 94102
rect 471306 94046 471374 94102
rect 471430 94046 471498 94102
rect 471554 94046 471622 94102
rect 471678 94046 489250 94102
rect 489306 94046 489374 94102
rect 489430 94046 489498 94102
rect 489554 94046 489622 94102
rect 489678 94046 507250 94102
rect 507306 94046 507374 94102
rect 507430 94046 507498 94102
rect 507554 94046 507622 94102
rect 507678 94046 524518 94102
rect 524574 94046 524642 94102
rect 524698 94046 525250 94102
rect 525306 94046 525374 94102
rect 525430 94046 525498 94102
rect 525554 94046 525622 94102
rect 525678 94046 543250 94102
rect 543306 94046 543374 94102
rect 543430 94046 543498 94102
rect 543554 94046 543622 94102
rect 543678 94046 555238 94102
rect 555294 94046 555362 94102
rect 555418 94046 561250 94102
rect 561306 94046 561374 94102
rect 561430 94046 561498 94102
rect 561554 94046 561622 94102
rect 561678 94046 579250 94102
rect 579306 94046 579374 94102
rect 579430 94046 579498 94102
rect 579554 94046 579622 94102
rect 579678 94046 596496 94102
rect 596552 94046 596620 94102
rect 596676 94046 596744 94102
rect 596800 94046 596868 94102
rect 596924 94046 597980 94102
rect -1916 93978 597980 94046
rect -1916 93922 -860 93978
rect -804 93922 -736 93978
rect -680 93922 -612 93978
rect -556 93922 -488 93978
rect -432 93922 3250 93978
rect 3306 93922 3374 93978
rect 3430 93922 3498 93978
rect 3554 93922 3622 93978
rect 3678 93922 21250 93978
rect 21306 93922 21374 93978
rect 21430 93922 21498 93978
rect 21554 93922 21622 93978
rect 21678 93922 39250 93978
rect 39306 93922 39374 93978
rect 39430 93922 39498 93978
rect 39554 93922 39622 93978
rect 39678 93922 183250 93978
rect 183306 93922 183374 93978
rect 183430 93922 183498 93978
rect 183554 93922 183622 93978
rect 183678 93922 201250 93978
rect 201306 93922 201374 93978
rect 201430 93922 201498 93978
rect 201554 93922 201622 93978
rect 201678 93922 381250 93978
rect 381306 93922 381374 93978
rect 381430 93922 381498 93978
rect 381554 93922 381622 93978
rect 381678 93922 399250 93978
rect 399306 93922 399374 93978
rect 399430 93922 399498 93978
rect 399554 93922 399622 93978
rect 399678 93922 417250 93978
rect 417306 93922 417374 93978
rect 417430 93922 417498 93978
rect 417554 93922 417622 93978
rect 417678 93922 435250 93978
rect 435306 93922 435374 93978
rect 435430 93922 435498 93978
rect 435554 93922 435622 93978
rect 435678 93922 453250 93978
rect 453306 93922 453374 93978
rect 453430 93922 453498 93978
rect 453554 93922 453622 93978
rect 453678 93922 471250 93978
rect 471306 93922 471374 93978
rect 471430 93922 471498 93978
rect 471554 93922 471622 93978
rect 471678 93922 489250 93978
rect 489306 93922 489374 93978
rect 489430 93922 489498 93978
rect 489554 93922 489622 93978
rect 489678 93922 507250 93978
rect 507306 93922 507374 93978
rect 507430 93922 507498 93978
rect 507554 93922 507622 93978
rect 507678 93922 524518 93978
rect 524574 93922 524642 93978
rect 524698 93922 525250 93978
rect 525306 93922 525374 93978
rect 525430 93922 525498 93978
rect 525554 93922 525622 93978
rect 525678 93922 543250 93978
rect 543306 93922 543374 93978
rect 543430 93922 543498 93978
rect 543554 93922 543622 93978
rect 543678 93922 555238 93978
rect 555294 93922 555362 93978
rect 555418 93922 561250 93978
rect 561306 93922 561374 93978
rect 561430 93922 561498 93978
rect 561554 93922 561622 93978
rect 561678 93922 579250 93978
rect 579306 93922 579374 93978
rect 579430 93922 579498 93978
rect 579554 93922 579622 93978
rect 579678 93922 596496 93978
rect 596552 93922 596620 93978
rect 596676 93922 596744 93978
rect 596800 93922 596868 93978
rect 596924 93922 597980 93978
rect -1916 93826 597980 93922
rect -1916 82350 597980 82446
rect -1916 82294 -1820 82350
rect -1764 82294 -1696 82350
rect -1640 82294 -1572 82350
rect -1516 82294 -1448 82350
rect -1392 82294 6970 82350
rect 7026 82294 7094 82350
rect 7150 82294 7218 82350
rect 7274 82294 7342 82350
rect 7398 82294 24970 82350
rect 25026 82294 25094 82350
rect 25150 82294 25218 82350
rect 25274 82294 25342 82350
rect 25398 82294 42970 82350
rect 43026 82294 43094 82350
rect 43150 82294 43218 82350
rect 43274 82294 43342 82350
rect 43398 82294 186970 82350
rect 187026 82294 187094 82350
rect 187150 82294 187218 82350
rect 187274 82294 187342 82350
rect 187398 82294 204970 82350
rect 205026 82294 205094 82350
rect 205150 82294 205218 82350
rect 205274 82294 205342 82350
rect 205398 82294 384970 82350
rect 385026 82294 385094 82350
rect 385150 82294 385218 82350
rect 385274 82294 385342 82350
rect 385398 82294 402970 82350
rect 403026 82294 403094 82350
rect 403150 82294 403218 82350
rect 403274 82294 403342 82350
rect 403398 82294 420970 82350
rect 421026 82294 421094 82350
rect 421150 82294 421218 82350
rect 421274 82294 421342 82350
rect 421398 82294 438970 82350
rect 439026 82294 439094 82350
rect 439150 82294 439218 82350
rect 439274 82294 439342 82350
rect 439398 82294 456970 82350
rect 457026 82294 457094 82350
rect 457150 82294 457218 82350
rect 457274 82294 457342 82350
rect 457398 82294 474970 82350
rect 475026 82294 475094 82350
rect 475150 82294 475218 82350
rect 475274 82294 475342 82350
rect 475398 82294 492970 82350
rect 493026 82294 493094 82350
rect 493150 82294 493218 82350
rect 493274 82294 493342 82350
rect 493398 82294 510970 82350
rect 511026 82294 511094 82350
rect 511150 82294 511218 82350
rect 511274 82294 511342 82350
rect 511398 82294 528970 82350
rect 529026 82294 529094 82350
rect 529150 82294 529218 82350
rect 529274 82294 529342 82350
rect 529398 82294 539878 82350
rect 539934 82294 540002 82350
rect 540058 82294 546970 82350
rect 547026 82294 547094 82350
rect 547150 82294 547218 82350
rect 547274 82294 547342 82350
rect 547398 82294 564970 82350
rect 565026 82294 565094 82350
rect 565150 82294 565218 82350
rect 565274 82294 565342 82350
rect 565398 82294 582970 82350
rect 583026 82294 583094 82350
rect 583150 82294 583218 82350
rect 583274 82294 583342 82350
rect 583398 82294 597456 82350
rect 597512 82294 597580 82350
rect 597636 82294 597704 82350
rect 597760 82294 597828 82350
rect 597884 82294 597980 82350
rect -1916 82226 597980 82294
rect -1916 82170 -1820 82226
rect -1764 82170 -1696 82226
rect -1640 82170 -1572 82226
rect -1516 82170 -1448 82226
rect -1392 82170 6970 82226
rect 7026 82170 7094 82226
rect 7150 82170 7218 82226
rect 7274 82170 7342 82226
rect 7398 82170 24970 82226
rect 25026 82170 25094 82226
rect 25150 82170 25218 82226
rect 25274 82170 25342 82226
rect 25398 82170 42970 82226
rect 43026 82170 43094 82226
rect 43150 82170 43218 82226
rect 43274 82170 43342 82226
rect 43398 82170 186970 82226
rect 187026 82170 187094 82226
rect 187150 82170 187218 82226
rect 187274 82170 187342 82226
rect 187398 82170 204970 82226
rect 205026 82170 205094 82226
rect 205150 82170 205218 82226
rect 205274 82170 205342 82226
rect 205398 82170 384970 82226
rect 385026 82170 385094 82226
rect 385150 82170 385218 82226
rect 385274 82170 385342 82226
rect 385398 82170 402970 82226
rect 403026 82170 403094 82226
rect 403150 82170 403218 82226
rect 403274 82170 403342 82226
rect 403398 82170 420970 82226
rect 421026 82170 421094 82226
rect 421150 82170 421218 82226
rect 421274 82170 421342 82226
rect 421398 82170 438970 82226
rect 439026 82170 439094 82226
rect 439150 82170 439218 82226
rect 439274 82170 439342 82226
rect 439398 82170 456970 82226
rect 457026 82170 457094 82226
rect 457150 82170 457218 82226
rect 457274 82170 457342 82226
rect 457398 82170 474970 82226
rect 475026 82170 475094 82226
rect 475150 82170 475218 82226
rect 475274 82170 475342 82226
rect 475398 82170 492970 82226
rect 493026 82170 493094 82226
rect 493150 82170 493218 82226
rect 493274 82170 493342 82226
rect 493398 82170 510970 82226
rect 511026 82170 511094 82226
rect 511150 82170 511218 82226
rect 511274 82170 511342 82226
rect 511398 82170 528970 82226
rect 529026 82170 529094 82226
rect 529150 82170 529218 82226
rect 529274 82170 529342 82226
rect 529398 82170 539878 82226
rect 539934 82170 540002 82226
rect 540058 82170 546970 82226
rect 547026 82170 547094 82226
rect 547150 82170 547218 82226
rect 547274 82170 547342 82226
rect 547398 82170 564970 82226
rect 565026 82170 565094 82226
rect 565150 82170 565218 82226
rect 565274 82170 565342 82226
rect 565398 82170 582970 82226
rect 583026 82170 583094 82226
rect 583150 82170 583218 82226
rect 583274 82170 583342 82226
rect 583398 82170 597456 82226
rect 597512 82170 597580 82226
rect 597636 82170 597704 82226
rect 597760 82170 597828 82226
rect 597884 82170 597980 82226
rect -1916 82102 597980 82170
rect -1916 82046 -1820 82102
rect -1764 82046 -1696 82102
rect -1640 82046 -1572 82102
rect -1516 82046 -1448 82102
rect -1392 82046 6970 82102
rect 7026 82046 7094 82102
rect 7150 82046 7218 82102
rect 7274 82046 7342 82102
rect 7398 82046 24970 82102
rect 25026 82046 25094 82102
rect 25150 82046 25218 82102
rect 25274 82046 25342 82102
rect 25398 82046 42970 82102
rect 43026 82046 43094 82102
rect 43150 82046 43218 82102
rect 43274 82046 43342 82102
rect 43398 82046 186970 82102
rect 187026 82046 187094 82102
rect 187150 82046 187218 82102
rect 187274 82046 187342 82102
rect 187398 82046 204970 82102
rect 205026 82046 205094 82102
rect 205150 82046 205218 82102
rect 205274 82046 205342 82102
rect 205398 82046 384970 82102
rect 385026 82046 385094 82102
rect 385150 82046 385218 82102
rect 385274 82046 385342 82102
rect 385398 82046 402970 82102
rect 403026 82046 403094 82102
rect 403150 82046 403218 82102
rect 403274 82046 403342 82102
rect 403398 82046 420970 82102
rect 421026 82046 421094 82102
rect 421150 82046 421218 82102
rect 421274 82046 421342 82102
rect 421398 82046 438970 82102
rect 439026 82046 439094 82102
rect 439150 82046 439218 82102
rect 439274 82046 439342 82102
rect 439398 82046 456970 82102
rect 457026 82046 457094 82102
rect 457150 82046 457218 82102
rect 457274 82046 457342 82102
rect 457398 82046 474970 82102
rect 475026 82046 475094 82102
rect 475150 82046 475218 82102
rect 475274 82046 475342 82102
rect 475398 82046 492970 82102
rect 493026 82046 493094 82102
rect 493150 82046 493218 82102
rect 493274 82046 493342 82102
rect 493398 82046 510970 82102
rect 511026 82046 511094 82102
rect 511150 82046 511218 82102
rect 511274 82046 511342 82102
rect 511398 82046 528970 82102
rect 529026 82046 529094 82102
rect 529150 82046 529218 82102
rect 529274 82046 529342 82102
rect 529398 82046 539878 82102
rect 539934 82046 540002 82102
rect 540058 82046 546970 82102
rect 547026 82046 547094 82102
rect 547150 82046 547218 82102
rect 547274 82046 547342 82102
rect 547398 82046 564970 82102
rect 565026 82046 565094 82102
rect 565150 82046 565218 82102
rect 565274 82046 565342 82102
rect 565398 82046 582970 82102
rect 583026 82046 583094 82102
rect 583150 82046 583218 82102
rect 583274 82046 583342 82102
rect 583398 82046 597456 82102
rect 597512 82046 597580 82102
rect 597636 82046 597704 82102
rect 597760 82046 597828 82102
rect 597884 82046 597980 82102
rect -1916 81978 597980 82046
rect -1916 81922 -1820 81978
rect -1764 81922 -1696 81978
rect -1640 81922 -1572 81978
rect -1516 81922 -1448 81978
rect -1392 81922 6970 81978
rect 7026 81922 7094 81978
rect 7150 81922 7218 81978
rect 7274 81922 7342 81978
rect 7398 81922 24970 81978
rect 25026 81922 25094 81978
rect 25150 81922 25218 81978
rect 25274 81922 25342 81978
rect 25398 81922 42970 81978
rect 43026 81922 43094 81978
rect 43150 81922 43218 81978
rect 43274 81922 43342 81978
rect 43398 81922 186970 81978
rect 187026 81922 187094 81978
rect 187150 81922 187218 81978
rect 187274 81922 187342 81978
rect 187398 81922 204970 81978
rect 205026 81922 205094 81978
rect 205150 81922 205218 81978
rect 205274 81922 205342 81978
rect 205398 81922 384970 81978
rect 385026 81922 385094 81978
rect 385150 81922 385218 81978
rect 385274 81922 385342 81978
rect 385398 81922 402970 81978
rect 403026 81922 403094 81978
rect 403150 81922 403218 81978
rect 403274 81922 403342 81978
rect 403398 81922 420970 81978
rect 421026 81922 421094 81978
rect 421150 81922 421218 81978
rect 421274 81922 421342 81978
rect 421398 81922 438970 81978
rect 439026 81922 439094 81978
rect 439150 81922 439218 81978
rect 439274 81922 439342 81978
rect 439398 81922 456970 81978
rect 457026 81922 457094 81978
rect 457150 81922 457218 81978
rect 457274 81922 457342 81978
rect 457398 81922 474970 81978
rect 475026 81922 475094 81978
rect 475150 81922 475218 81978
rect 475274 81922 475342 81978
rect 475398 81922 492970 81978
rect 493026 81922 493094 81978
rect 493150 81922 493218 81978
rect 493274 81922 493342 81978
rect 493398 81922 510970 81978
rect 511026 81922 511094 81978
rect 511150 81922 511218 81978
rect 511274 81922 511342 81978
rect 511398 81922 528970 81978
rect 529026 81922 529094 81978
rect 529150 81922 529218 81978
rect 529274 81922 529342 81978
rect 529398 81922 539878 81978
rect 539934 81922 540002 81978
rect 540058 81922 546970 81978
rect 547026 81922 547094 81978
rect 547150 81922 547218 81978
rect 547274 81922 547342 81978
rect 547398 81922 564970 81978
rect 565026 81922 565094 81978
rect 565150 81922 565218 81978
rect 565274 81922 565342 81978
rect 565398 81922 582970 81978
rect 583026 81922 583094 81978
rect 583150 81922 583218 81978
rect 583274 81922 583342 81978
rect 583398 81922 597456 81978
rect 597512 81922 597580 81978
rect 597636 81922 597704 81978
rect 597760 81922 597828 81978
rect 597884 81922 597980 81978
rect -1916 81826 597980 81922
rect -1916 76350 597980 76446
rect -1916 76294 -860 76350
rect -804 76294 -736 76350
rect -680 76294 -612 76350
rect -556 76294 -488 76350
rect -432 76294 3250 76350
rect 3306 76294 3374 76350
rect 3430 76294 3498 76350
rect 3554 76294 3622 76350
rect 3678 76294 21250 76350
rect 21306 76294 21374 76350
rect 21430 76294 21498 76350
rect 21554 76294 21622 76350
rect 21678 76294 39250 76350
rect 39306 76294 39374 76350
rect 39430 76294 39498 76350
rect 39554 76294 39622 76350
rect 39678 76294 57250 76350
rect 57306 76294 57374 76350
rect 57430 76294 57498 76350
rect 57554 76294 57622 76350
rect 57678 76294 75250 76350
rect 75306 76294 75374 76350
rect 75430 76294 75498 76350
rect 75554 76294 75622 76350
rect 75678 76294 93250 76350
rect 93306 76294 93374 76350
rect 93430 76294 93498 76350
rect 93554 76294 93622 76350
rect 93678 76294 111250 76350
rect 111306 76294 111374 76350
rect 111430 76294 111498 76350
rect 111554 76294 111622 76350
rect 111678 76294 129250 76350
rect 129306 76294 129374 76350
rect 129430 76294 129498 76350
rect 129554 76294 129622 76350
rect 129678 76294 147250 76350
rect 147306 76294 147374 76350
rect 147430 76294 147498 76350
rect 147554 76294 147622 76350
rect 147678 76294 165250 76350
rect 165306 76294 165374 76350
rect 165430 76294 165498 76350
rect 165554 76294 165622 76350
rect 165678 76294 183250 76350
rect 183306 76294 183374 76350
rect 183430 76294 183498 76350
rect 183554 76294 183622 76350
rect 183678 76294 201250 76350
rect 201306 76294 201374 76350
rect 201430 76294 201498 76350
rect 201554 76294 201622 76350
rect 201678 76294 381250 76350
rect 381306 76294 381374 76350
rect 381430 76294 381498 76350
rect 381554 76294 381622 76350
rect 381678 76294 399250 76350
rect 399306 76294 399374 76350
rect 399430 76294 399498 76350
rect 399554 76294 399622 76350
rect 399678 76294 417250 76350
rect 417306 76294 417374 76350
rect 417430 76294 417498 76350
rect 417554 76294 417622 76350
rect 417678 76294 435250 76350
rect 435306 76294 435374 76350
rect 435430 76294 435498 76350
rect 435554 76294 435622 76350
rect 435678 76294 453250 76350
rect 453306 76294 453374 76350
rect 453430 76294 453498 76350
rect 453554 76294 453622 76350
rect 453678 76294 471250 76350
rect 471306 76294 471374 76350
rect 471430 76294 471498 76350
rect 471554 76294 471622 76350
rect 471678 76294 489250 76350
rect 489306 76294 489374 76350
rect 489430 76294 489498 76350
rect 489554 76294 489622 76350
rect 489678 76294 507250 76350
rect 507306 76294 507374 76350
rect 507430 76294 507498 76350
rect 507554 76294 507622 76350
rect 507678 76294 524518 76350
rect 524574 76294 524642 76350
rect 524698 76294 525250 76350
rect 525306 76294 525374 76350
rect 525430 76294 525498 76350
rect 525554 76294 525622 76350
rect 525678 76294 543250 76350
rect 543306 76294 543374 76350
rect 543430 76294 543498 76350
rect 543554 76294 543622 76350
rect 543678 76294 555238 76350
rect 555294 76294 555362 76350
rect 555418 76294 561250 76350
rect 561306 76294 561374 76350
rect 561430 76294 561498 76350
rect 561554 76294 561622 76350
rect 561678 76294 579250 76350
rect 579306 76294 579374 76350
rect 579430 76294 579498 76350
rect 579554 76294 579622 76350
rect 579678 76294 596496 76350
rect 596552 76294 596620 76350
rect 596676 76294 596744 76350
rect 596800 76294 596868 76350
rect 596924 76294 597980 76350
rect -1916 76226 597980 76294
rect -1916 76170 -860 76226
rect -804 76170 -736 76226
rect -680 76170 -612 76226
rect -556 76170 -488 76226
rect -432 76170 3250 76226
rect 3306 76170 3374 76226
rect 3430 76170 3498 76226
rect 3554 76170 3622 76226
rect 3678 76170 21250 76226
rect 21306 76170 21374 76226
rect 21430 76170 21498 76226
rect 21554 76170 21622 76226
rect 21678 76170 39250 76226
rect 39306 76170 39374 76226
rect 39430 76170 39498 76226
rect 39554 76170 39622 76226
rect 39678 76170 57250 76226
rect 57306 76170 57374 76226
rect 57430 76170 57498 76226
rect 57554 76170 57622 76226
rect 57678 76170 75250 76226
rect 75306 76170 75374 76226
rect 75430 76170 75498 76226
rect 75554 76170 75622 76226
rect 75678 76170 93250 76226
rect 93306 76170 93374 76226
rect 93430 76170 93498 76226
rect 93554 76170 93622 76226
rect 93678 76170 111250 76226
rect 111306 76170 111374 76226
rect 111430 76170 111498 76226
rect 111554 76170 111622 76226
rect 111678 76170 129250 76226
rect 129306 76170 129374 76226
rect 129430 76170 129498 76226
rect 129554 76170 129622 76226
rect 129678 76170 147250 76226
rect 147306 76170 147374 76226
rect 147430 76170 147498 76226
rect 147554 76170 147622 76226
rect 147678 76170 165250 76226
rect 165306 76170 165374 76226
rect 165430 76170 165498 76226
rect 165554 76170 165622 76226
rect 165678 76170 183250 76226
rect 183306 76170 183374 76226
rect 183430 76170 183498 76226
rect 183554 76170 183622 76226
rect 183678 76170 201250 76226
rect 201306 76170 201374 76226
rect 201430 76170 201498 76226
rect 201554 76170 201622 76226
rect 201678 76170 381250 76226
rect 381306 76170 381374 76226
rect 381430 76170 381498 76226
rect 381554 76170 381622 76226
rect 381678 76170 399250 76226
rect 399306 76170 399374 76226
rect 399430 76170 399498 76226
rect 399554 76170 399622 76226
rect 399678 76170 417250 76226
rect 417306 76170 417374 76226
rect 417430 76170 417498 76226
rect 417554 76170 417622 76226
rect 417678 76170 435250 76226
rect 435306 76170 435374 76226
rect 435430 76170 435498 76226
rect 435554 76170 435622 76226
rect 435678 76170 453250 76226
rect 453306 76170 453374 76226
rect 453430 76170 453498 76226
rect 453554 76170 453622 76226
rect 453678 76170 471250 76226
rect 471306 76170 471374 76226
rect 471430 76170 471498 76226
rect 471554 76170 471622 76226
rect 471678 76170 489250 76226
rect 489306 76170 489374 76226
rect 489430 76170 489498 76226
rect 489554 76170 489622 76226
rect 489678 76170 507250 76226
rect 507306 76170 507374 76226
rect 507430 76170 507498 76226
rect 507554 76170 507622 76226
rect 507678 76170 524518 76226
rect 524574 76170 524642 76226
rect 524698 76170 525250 76226
rect 525306 76170 525374 76226
rect 525430 76170 525498 76226
rect 525554 76170 525622 76226
rect 525678 76170 543250 76226
rect 543306 76170 543374 76226
rect 543430 76170 543498 76226
rect 543554 76170 543622 76226
rect 543678 76170 555238 76226
rect 555294 76170 555362 76226
rect 555418 76170 561250 76226
rect 561306 76170 561374 76226
rect 561430 76170 561498 76226
rect 561554 76170 561622 76226
rect 561678 76170 579250 76226
rect 579306 76170 579374 76226
rect 579430 76170 579498 76226
rect 579554 76170 579622 76226
rect 579678 76170 596496 76226
rect 596552 76170 596620 76226
rect 596676 76170 596744 76226
rect 596800 76170 596868 76226
rect 596924 76170 597980 76226
rect -1916 76102 597980 76170
rect -1916 76046 -860 76102
rect -804 76046 -736 76102
rect -680 76046 -612 76102
rect -556 76046 -488 76102
rect -432 76046 3250 76102
rect 3306 76046 3374 76102
rect 3430 76046 3498 76102
rect 3554 76046 3622 76102
rect 3678 76046 21250 76102
rect 21306 76046 21374 76102
rect 21430 76046 21498 76102
rect 21554 76046 21622 76102
rect 21678 76046 39250 76102
rect 39306 76046 39374 76102
rect 39430 76046 39498 76102
rect 39554 76046 39622 76102
rect 39678 76046 57250 76102
rect 57306 76046 57374 76102
rect 57430 76046 57498 76102
rect 57554 76046 57622 76102
rect 57678 76046 75250 76102
rect 75306 76046 75374 76102
rect 75430 76046 75498 76102
rect 75554 76046 75622 76102
rect 75678 76046 93250 76102
rect 93306 76046 93374 76102
rect 93430 76046 93498 76102
rect 93554 76046 93622 76102
rect 93678 76046 111250 76102
rect 111306 76046 111374 76102
rect 111430 76046 111498 76102
rect 111554 76046 111622 76102
rect 111678 76046 129250 76102
rect 129306 76046 129374 76102
rect 129430 76046 129498 76102
rect 129554 76046 129622 76102
rect 129678 76046 147250 76102
rect 147306 76046 147374 76102
rect 147430 76046 147498 76102
rect 147554 76046 147622 76102
rect 147678 76046 165250 76102
rect 165306 76046 165374 76102
rect 165430 76046 165498 76102
rect 165554 76046 165622 76102
rect 165678 76046 183250 76102
rect 183306 76046 183374 76102
rect 183430 76046 183498 76102
rect 183554 76046 183622 76102
rect 183678 76046 201250 76102
rect 201306 76046 201374 76102
rect 201430 76046 201498 76102
rect 201554 76046 201622 76102
rect 201678 76046 381250 76102
rect 381306 76046 381374 76102
rect 381430 76046 381498 76102
rect 381554 76046 381622 76102
rect 381678 76046 399250 76102
rect 399306 76046 399374 76102
rect 399430 76046 399498 76102
rect 399554 76046 399622 76102
rect 399678 76046 417250 76102
rect 417306 76046 417374 76102
rect 417430 76046 417498 76102
rect 417554 76046 417622 76102
rect 417678 76046 435250 76102
rect 435306 76046 435374 76102
rect 435430 76046 435498 76102
rect 435554 76046 435622 76102
rect 435678 76046 453250 76102
rect 453306 76046 453374 76102
rect 453430 76046 453498 76102
rect 453554 76046 453622 76102
rect 453678 76046 471250 76102
rect 471306 76046 471374 76102
rect 471430 76046 471498 76102
rect 471554 76046 471622 76102
rect 471678 76046 489250 76102
rect 489306 76046 489374 76102
rect 489430 76046 489498 76102
rect 489554 76046 489622 76102
rect 489678 76046 507250 76102
rect 507306 76046 507374 76102
rect 507430 76046 507498 76102
rect 507554 76046 507622 76102
rect 507678 76046 524518 76102
rect 524574 76046 524642 76102
rect 524698 76046 525250 76102
rect 525306 76046 525374 76102
rect 525430 76046 525498 76102
rect 525554 76046 525622 76102
rect 525678 76046 543250 76102
rect 543306 76046 543374 76102
rect 543430 76046 543498 76102
rect 543554 76046 543622 76102
rect 543678 76046 555238 76102
rect 555294 76046 555362 76102
rect 555418 76046 561250 76102
rect 561306 76046 561374 76102
rect 561430 76046 561498 76102
rect 561554 76046 561622 76102
rect 561678 76046 579250 76102
rect 579306 76046 579374 76102
rect 579430 76046 579498 76102
rect 579554 76046 579622 76102
rect 579678 76046 596496 76102
rect 596552 76046 596620 76102
rect 596676 76046 596744 76102
rect 596800 76046 596868 76102
rect 596924 76046 597980 76102
rect -1916 75978 597980 76046
rect -1916 75922 -860 75978
rect -804 75922 -736 75978
rect -680 75922 -612 75978
rect -556 75922 -488 75978
rect -432 75922 3250 75978
rect 3306 75922 3374 75978
rect 3430 75922 3498 75978
rect 3554 75922 3622 75978
rect 3678 75922 21250 75978
rect 21306 75922 21374 75978
rect 21430 75922 21498 75978
rect 21554 75922 21622 75978
rect 21678 75922 39250 75978
rect 39306 75922 39374 75978
rect 39430 75922 39498 75978
rect 39554 75922 39622 75978
rect 39678 75922 57250 75978
rect 57306 75922 57374 75978
rect 57430 75922 57498 75978
rect 57554 75922 57622 75978
rect 57678 75922 75250 75978
rect 75306 75922 75374 75978
rect 75430 75922 75498 75978
rect 75554 75922 75622 75978
rect 75678 75922 93250 75978
rect 93306 75922 93374 75978
rect 93430 75922 93498 75978
rect 93554 75922 93622 75978
rect 93678 75922 111250 75978
rect 111306 75922 111374 75978
rect 111430 75922 111498 75978
rect 111554 75922 111622 75978
rect 111678 75922 129250 75978
rect 129306 75922 129374 75978
rect 129430 75922 129498 75978
rect 129554 75922 129622 75978
rect 129678 75922 147250 75978
rect 147306 75922 147374 75978
rect 147430 75922 147498 75978
rect 147554 75922 147622 75978
rect 147678 75922 165250 75978
rect 165306 75922 165374 75978
rect 165430 75922 165498 75978
rect 165554 75922 165622 75978
rect 165678 75922 183250 75978
rect 183306 75922 183374 75978
rect 183430 75922 183498 75978
rect 183554 75922 183622 75978
rect 183678 75922 201250 75978
rect 201306 75922 201374 75978
rect 201430 75922 201498 75978
rect 201554 75922 201622 75978
rect 201678 75922 381250 75978
rect 381306 75922 381374 75978
rect 381430 75922 381498 75978
rect 381554 75922 381622 75978
rect 381678 75922 399250 75978
rect 399306 75922 399374 75978
rect 399430 75922 399498 75978
rect 399554 75922 399622 75978
rect 399678 75922 417250 75978
rect 417306 75922 417374 75978
rect 417430 75922 417498 75978
rect 417554 75922 417622 75978
rect 417678 75922 435250 75978
rect 435306 75922 435374 75978
rect 435430 75922 435498 75978
rect 435554 75922 435622 75978
rect 435678 75922 453250 75978
rect 453306 75922 453374 75978
rect 453430 75922 453498 75978
rect 453554 75922 453622 75978
rect 453678 75922 471250 75978
rect 471306 75922 471374 75978
rect 471430 75922 471498 75978
rect 471554 75922 471622 75978
rect 471678 75922 489250 75978
rect 489306 75922 489374 75978
rect 489430 75922 489498 75978
rect 489554 75922 489622 75978
rect 489678 75922 507250 75978
rect 507306 75922 507374 75978
rect 507430 75922 507498 75978
rect 507554 75922 507622 75978
rect 507678 75922 524518 75978
rect 524574 75922 524642 75978
rect 524698 75922 525250 75978
rect 525306 75922 525374 75978
rect 525430 75922 525498 75978
rect 525554 75922 525622 75978
rect 525678 75922 543250 75978
rect 543306 75922 543374 75978
rect 543430 75922 543498 75978
rect 543554 75922 543622 75978
rect 543678 75922 555238 75978
rect 555294 75922 555362 75978
rect 555418 75922 561250 75978
rect 561306 75922 561374 75978
rect 561430 75922 561498 75978
rect 561554 75922 561622 75978
rect 561678 75922 579250 75978
rect 579306 75922 579374 75978
rect 579430 75922 579498 75978
rect 579554 75922 579622 75978
rect 579678 75922 596496 75978
rect 596552 75922 596620 75978
rect 596676 75922 596744 75978
rect 596800 75922 596868 75978
rect 596924 75922 597980 75978
rect -1916 75826 597980 75922
rect -1916 64350 597980 64446
rect -1916 64294 -1820 64350
rect -1764 64294 -1696 64350
rect -1640 64294 -1572 64350
rect -1516 64294 -1448 64350
rect -1392 64294 6970 64350
rect 7026 64294 7094 64350
rect 7150 64294 7218 64350
rect 7274 64294 7342 64350
rect 7398 64294 24970 64350
rect 25026 64294 25094 64350
rect 25150 64294 25218 64350
rect 25274 64294 25342 64350
rect 25398 64294 42970 64350
rect 43026 64294 43094 64350
rect 43150 64294 43218 64350
rect 43274 64294 43342 64350
rect 43398 64294 60970 64350
rect 61026 64294 61094 64350
rect 61150 64294 61218 64350
rect 61274 64294 61342 64350
rect 61398 64294 78970 64350
rect 79026 64294 79094 64350
rect 79150 64294 79218 64350
rect 79274 64294 79342 64350
rect 79398 64294 96970 64350
rect 97026 64294 97094 64350
rect 97150 64294 97218 64350
rect 97274 64294 97342 64350
rect 97398 64294 114970 64350
rect 115026 64294 115094 64350
rect 115150 64294 115218 64350
rect 115274 64294 115342 64350
rect 115398 64294 132970 64350
rect 133026 64294 133094 64350
rect 133150 64294 133218 64350
rect 133274 64294 133342 64350
rect 133398 64294 150970 64350
rect 151026 64294 151094 64350
rect 151150 64294 151218 64350
rect 151274 64294 151342 64350
rect 151398 64294 168970 64350
rect 169026 64294 169094 64350
rect 169150 64294 169218 64350
rect 169274 64294 169342 64350
rect 169398 64294 186970 64350
rect 187026 64294 187094 64350
rect 187150 64294 187218 64350
rect 187274 64294 187342 64350
rect 187398 64294 204970 64350
rect 205026 64294 205094 64350
rect 205150 64294 205218 64350
rect 205274 64294 205342 64350
rect 205398 64294 384970 64350
rect 385026 64294 385094 64350
rect 385150 64294 385218 64350
rect 385274 64294 385342 64350
rect 385398 64294 402970 64350
rect 403026 64294 403094 64350
rect 403150 64294 403218 64350
rect 403274 64294 403342 64350
rect 403398 64294 420970 64350
rect 421026 64294 421094 64350
rect 421150 64294 421218 64350
rect 421274 64294 421342 64350
rect 421398 64294 438970 64350
rect 439026 64294 439094 64350
rect 439150 64294 439218 64350
rect 439274 64294 439342 64350
rect 439398 64294 456970 64350
rect 457026 64294 457094 64350
rect 457150 64294 457218 64350
rect 457274 64294 457342 64350
rect 457398 64294 474970 64350
rect 475026 64294 475094 64350
rect 475150 64294 475218 64350
rect 475274 64294 475342 64350
rect 475398 64294 492970 64350
rect 493026 64294 493094 64350
rect 493150 64294 493218 64350
rect 493274 64294 493342 64350
rect 493398 64294 510970 64350
rect 511026 64294 511094 64350
rect 511150 64294 511218 64350
rect 511274 64294 511342 64350
rect 511398 64294 528970 64350
rect 529026 64294 529094 64350
rect 529150 64294 529218 64350
rect 529274 64294 529342 64350
rect 529398 64294 539878 64350
rect 539934 64294 540002 64350
rect 540058 64294 546970 64350
rect 547026 64294 547094 64350
rect 547150 64294 547218 64350
rect 547274 64294 547342 64350
rect 547398 64294 564970 64350
rect 565026 64294 565094 64350
rect 565150 64294 565218 64350
rect 565274 64294 565342 64350
rect 565398 64294 582970 64350
rect 583026 64294 583094 64350
rect 583150 64294 583218 64350
rect 583274 64294 583342 64350
rect 583398 64294 597456 64350
rect 597512 64294 597580 64350
rect 597636 64294 597704 64350
rect 597760 64294 597828 64350
rect 597884 64294 597980 64350
rect -1916 64226 597980 64294
rect -1916 64170 -1820 64226
rect -1764 64170 -1696 64226
rect -1640 64170 -1572 64226
rect -1516 64170 -1448 64226
rect -1392 64170 6970 64226
rect 7026 64170 7094 64226
rect 7150 64170 7218 64226
rect 7274 64170 7342 64226
rect 7398 64170 24970 64226
rect 25026 64170 25094 64226
rect 25150 64170 25218 64226
rect 25274 64170 25342 64226
rect 25398 64170 42970 64226
rect 43026 64170 43094 64226
rect 43150 64170 43218 64226
rect 43274 64170 43342 64226
rect 43398 64170 60970 64226
rect 61026 64170 61094 64226
rect 61150 64170 61218 64226
rect 61274 64170 61342 64226
rect 61398 64170 78970 64226
rect 79026 64170 79094 64226
rect 79150 64170 79218 64226
rect 79274 64170 79342 64226
rect 79398 64170 96970 64226
rect 97026 64170 97094 64226
rect 97150 64170 97218 64226
rect 97274 64170 97342 64226
rect 97398 64170 114970 64226
rect 115026 64170 115094 64226
rect 115150 64170 115218 64226
rect 115274 64170 115342 64226
rect 115398 64170 132970 64226
rect 133026 64170 133094 64226
rect 133150 64170 133218 64226
rect 133274 64170 133342 64226
rect 133398 64170 150970 64226
rect 151026 64170 151094 64226
rect 151150 64170 151218 64226
rect 151274 64170 151342 64226
rect 151398 64170 168970 64226
rect 169026 64170 169094 64226
rect 169150 64170 169218 64226
rect 169274 64170 169342 64226
rect 169398 64170 186970 64226
rect 187026 64170 187094 64226
rect 187150 64170 187218 64226
rect 187274 64170 187342 64226
rect 187398 64170 204970 64226
rect 205026 64170 205094 64226
rect 205150 64170 205218 64226
rect 205274 64170 205342 64226
rect 205398 64170 384970 64226
rect 385026 64170 385094 64226
rect 385150 64170 385218 64226
rect 385274 64170 385342 64226
rect 385398 64170 402970 64226
rect 403026 64170 403094 64226
rect 403150 64170 403218 64226
rect 403274 64170 403342 64226
rect 403398 64170 420970 64226
rect 421026 64170 421094 64226
rect 421150 64170 421218 64226
rect 421274 64170 421342 64226
rect 421398 64170 438970 64226
rect 439026 64170 439094 64226
rect 439150 64170 439218 64226
rect 439274 64170 439342 64226
rect 439398 64170 456970 64226
rect 457026 64170 457094 64226
rect 457150 64170 457218 64226
rect 457274 64170 457342 64226
rect 457398 64170 474970 64226
rect 475026 64170 475094 64226
rect 475150 64170 475218 64226
rect 475274 64170 475342 64226
rect 475398 64170 492970 64226
rect 493026 64170 493094 64226
rect 493150 64170 493218 64226
rect 493274 64170 493342 64226
rect 493398 64170 510970 64226
rect 511026 64170 511094 64226
rect 511150 64170 511218 64226
rect 511274 64170 511342 64226
rect 511398 64170 528970 64226
rect 529026 64170 529094 64226
rect 529150 64170 529218 64226
rect 529274 64170 529342 64226
rect 529398 64170 539878 64226
rect 539934 64170 540002 64226
rect 540058 64170 546970 64226
rect 547026 64170 547094 64226
rect 547150 64170 547218 64226
rect 547274 64170 547342 64226
rect 547398 64170 564970 64226
rect 565026 64170 565094 64226
rect 565150 64170 565218 64226
rect 565274 64170 565342 64226
rect 565398 64170 582970 64226
rect 583026 64170 583094 64226
rect 583150 64170 583218 64226
rect 583274 64170 583342 64226
rect 583398 64170 597456 64226
rect 597512 64170 597580 64226
rect 597636 64170 597704 64226
rect 597760 64170 597828 64226
rect 597884 64170 597980 64226
rect -1916 64102 597980 64170
rect -1916 64046 -1820 64102
rect -1764 64046 -1696 64102
rect -1640 64046 -1572 64102
rect -1516 64046 -1448 64102
rect -1392 64046 6970 64102
rect 7026 64046 7094 64102
rect 7150 64046 7218 64102
rect 7274 64046 7342 64102
rect 7398 64046 24970 64102
rect 25026 64046 25094 64102
rect 25150 64046 25218 64102
rect 25274 64046 25342 64102
rect 25398 64046 42970 64102
rect 43026 64046 43094 64102
rect 43150 64046 43218 64102
rect 43274 64046 43342 64102
rect 43398 64046 60970 64102
rect 61026 64046 61094 64102
rect 61150 64046 61218 64102
rect 61274 64046 61342 64102
rect 61398 64046 78970 64102
rect 79026 64046 79094 64102
rect 79150 64046 79218 64102
rect 79274 64046 79342 64102
rect 79398 64046 96970 64102
rect 97026 64046 97094 64102
rect 97150 64046 97218 64102
rect 97274 64046 97342 64102
rect 97398 64046 114970 64102
rect 115026 64046 115094 64102
rect 115150 64046 115218 64102
rect 115274 64046 115342 64102
rect 115398 64046 132970 64102
rect 133026 64046 133094 64102
rect 133150 64046 133218 64102
rect 133274 64046 133342 64102
rect 133398 64046 150970 64102
rect 151026 64046 151094 64102
rect 151150 64046 151218 64102
rect 151274 64046 151342 64102
rect 151398 64046 168970 64102
rect 169026 64046 169094 64102
rect 169150 64046 169218 64102
rect 169274 64046 169342 64102
rect 169398 64046 186970 64102
rect 187026 64046 187094 64102
rect 187150 64046 187218 64102
rect 187274 64046 187342 64102
rect 187398 64046 204970 64102
rect 205026 64046 205094 64102
rect 205150 64046 205218 64102
rect 205274 64046 205342 64102
rect 205398 64046 384970 64102
rect 385026 64046 385094 64102
rect 385150 64046 385218 64102
rect 385274 64046 385342 64102
rect 385398 64046 402970 64102
rect 403026 64046 403094 64102
rect 403150 64046 403218 64102
rect 403274 64046 403342 64102
rect 403398 64046 420970 64102
rect 421026 64046 421094 64102
rect 421150 64046 421218 64102
rect 421274 64046 421342 64102
rect 421398 64046 438970 64102
rect 439026 64046 439094 64102
rect 439150 64046 439218 64102
rect 439274 64046 439342 64102
rect 439398 64046 456970 64102
rect 457026 64046 457094 64102
rect 457150 64046 457218 64102
rect 457274 64046 457342 64102
rect 457398 64046 474970 64102
rect 475026 64046 475094 64102
rect 475150 64046 475218 64102
rect 475274 64046 475342 64102
rect 475398 64046 492970 64102
rect 493026 64046 493094 64102
rect 493150 64046 493218 64102
rect 493274 64046 493342 64102
rect 493398 64046 510970 64102
rect 511026 64046 511094 64102
rect 511150 64046 511218 64102
rect 511274 64046 511342 64102
rect 511398 64046 528970 64102
rect 529026 64046 529094 64102
rect 529150 64046 529218 64102
rect 529274 64046 529342 64102
rect 529398 64046 539878 64102
rect 539934 64046 540002 64102
rect 540058 64046 546970 64102
rect 547026 64046 547094 64102
rect 547150 64046 547218 64102
rect 547274 64046 547342 64102
rect 547398 64046 564970 64102
rect 565026 64046 565094 64102
rect 565150 64046 565218 64102
rect 565274 64046 565342 64102
rect 565398 64046 582970 64102
rect 583026 64046 583094 64102
rect 583150 64046 583218 64102
rect 583274 64046 583342 64102
rect 583398 64046 597456 64102
rect 597512 64046 597580 64102
rect 597636 64046 597704 64102
rect 597760 64046 597828 64102
rect 597884 64046 597980 64102
rect -1916 63978 597980 64046
rect -1916 63922 -1820 63978
rect -1764 63922 -1696 63978
rect -1640 63922 -1572 63978
rect -1516 63922 -1448 63978
rect -1392 63922 6970 63978
rect 7026 63922 7094 63978
rect 7150 63922 7218 63978
rect 7274 63922 7342 63978
rect 7398 63922 24970 63978
rect 25026 63922 25094 63978
rect 25150 63922 25218 63978
rect 25274 63922 25342 63978
rect 25398 63922 42970 63978
rect 43026 63922 43094 63978
rect 43150 63922 43218 63978
rect 43274 63922 43342 63978
rect 43398 63922 60970 63978
rect 61026 63922 61094 63978
rect 61150 63922 61218 63978
rect 61274 63922 61342 63978
rect 61398 63922 78970 63978
rect 79026 63922 79094 63978
rect 79150 63922 79218 63978
rect 79274 63922 79342 63978
rect 79398 63922 96970 63978
rect 97026 63922 97094 63978
rect 97150 63922 97218 63978
rect 97274 63922 97342 63978
rect 97398 63922 114970 63978
rect 115026 63922 115094 63978
rect 115150 63922 115218 63978
rect 115274 63922 115342 63978
rect 115398 63922 132970 63978
rect 133026 63922 133094 63978
rect 133150 63922 133218 63978
rect 133274 63922 133342 63978
rect 133398 63922 150970 63978
rect 151026 63922 151094 63978
rect 151150 63922 151218 63978
rect 151274 63922 151342 63978
rect 151398 63922 168970 63978
rect 169026 63922 169094 63978
rect 169150 63922 169218 63978
rect 169274 63922 169342 63978
rect 169398 63922 186970 63978
rect 187026 63922 187094 63978
rect 187150 63922 187218 63978
rect 187274 63922 187342 63978
rect 187398 63922 204970 63978
rect 205026 63922 205094 63978
rect 205150 63922 205218 63978
rect 205274 63922 205342 63978
rect 205398 63922 384970 63978
rect 385026 63922 385094 63978
rect 385150 63922 385218 63978
rect 385274 63922 385342 63978
rect 385398 63922 402970 63978
rect 403026 63922 403094 63978
rect 403150 63922 403218 63978
rect 403274 63922 403342 63978
rect 403398 63922 420970 63978
rect 421026 63922 421094 63978
rect 421150 63922 421218 63978
rect 421274 63922 421342 63978
rect 421398 63922 438970 63978
rect 439026 63922 439094 63978
rect 439150 63922 439218 63978
rect 439274 63922 439342 63978
rect 439398 63922 456970 63978
rect 457026 63922 457094 63978
rect 457150 63922 457218 63978
rect 457274 63922 457342 63978
rect 457398 63922 474970 63978
rect 475026 63922 475094 63978
rect 475150 63922 475218 63978
rect 475274 63922 475342 63978
rect 475398 63922 492970 63978
rect 493026 63922 493094 63978
rect 493150 63922 493218 63978
rect 493274 63922 493342 63978
rect 493398 63922 510970 63978
rect 511026 63922 511094 63978
rect 511150 63922 511218 63978
rect 511274 63922 511342 63978
rect 511398 63922 528970 63978
rect 529026 63922 529094 63978
rect 529150 63922 529218 63978
rect 529274 63922 529342 63978
rect 529398 63922 539878 63978
rect 539934 63922 540002 63978
rect 540058 63922 546970 63978
rect 547026 63922 547094 63978
rect 547150 63922 547218 63978
rect 547274 63922 547342 63978
rect 547398 63922 564970 63978
rect 565026 63922 565094 63978
rect 565150 63922 565218 63978
rect 565274 63922 565342 63978
rect 565398 63922 582970 63978
rect 583026 63922 583094 63978
rect 583150 63922 583218 63978
rect 583274 63922 583342 63978
rect 583398 63922 597456 63978
rect 597512 63922 597580 63978
rect 597636 63922 597704 63978
rect 597760 63922 597828 63978
rect 597884 63922 597980 63978
rect -1916 63826 597980 63922
rect -1916 58350 597980 58446
rect -1916 58294 -860 58350
rect -804 58294 -736 58350
rect -680 58294 -612 58350
rect -556 58294 -488 58350
rect -432 58294 3250 58350
rect 3306 58294 3374 58350
rect 3430 58294 3498 58350
rect 3554 58294 3622 58350
rect 3678 58294 21250 58350
rect 21306 58294 21374 58350
rect 21430 58294 21498 58350
rect 21554 58294 21622 58350
rect 21678 58294 39250 58350
rect 39306 58294 39374 58350
rect 39430 58294 39498 58350
rect 39554 58294 39622 58350
rect 39678 58294 57250 58350
rect 57306 58294 57374 58350
rect 57430 58294 57498 58350
rect 57554 58294 57622 58350
rect 57678 58294 75250 58350
rect 75306 58294 75374 58350
rect 75430 58294 75498 58350
rect 75554 58294 75622 58350
rect 75678 58294 93250 58350
rect 93306 58294 93374 58350
rect 93430 58294 93498 58350
rect 93554 58294 93622 58350
rect 93678 58294 111250 58350
rect 111306 58294 111374 58350
rect 111430 58294 111498 58350
rect 111554 58294 111622 58350
rect 111678 58294 129250 58350
rect 129306 58294 129374 58350
rect 129430 58294 129498 58350
rect 129554 58294 129622 58350
rect 129678 58294 147250 58350
rect 147306 58294 147374 58350
rect 147430 58294 147498 58350
rect 147554 58294 147622 58350
rect 147678 58294 165250 58350
rect 165306 58294 165374 58350
rect 165430 58294 165498 58350
rect 165554 58294 165622 58350
rect 165678 58294 183250 58350
rect 183306 58294 183374 58350
rect 183430 58294 183498 58350
rect 183554 58294 183622 58350
rect 183678 58294 201250 58350
rect 201306 58294 201374 58350
rect 201430 58294 201498 58350
rect 201554 58294 201622 58350
rect 201678 58294 381250 58350
rect 381306 58294 381374 58350
rect 381430 58294 381498 58350
rect 381554 58294 381622 58350
rect 381678 58294 399250 58350
rect 399306 58294 399374 58350
rect 399430 58294 399498 58350
rect 399554 58294 399622 58350
rect 399678 58294 417250 58350
rect 417306 58294 417374 58350
rect 417430 58294 417498 58350
rect 417554 58294 417622 58350
rect 417678 58294 435250 58350
rect 435306 58294 435374 58350
rect 435430 58294 435498 58350
rect 435554 58294 435622 58350
rect 435678 58294 453250 58350
rect 453306 58294 453374 58350
rect 453430 58294 453498 58350
rect 453554 58294 453622 58350
rect 453678 58294 471250 58350
rect 471306 58294 471374 58350
rect 471430 58294 471498 58350
rect 471554 58294 471622 58350
rect 471678 58294 489250 58350
rect 489306 58294 489374 58350
rect 489430 58294 489498 58350
rect 489554 58294 489622 58350
rect 489678 58294 507250 58350
rect 507306 58294 507374 58350
rect 507430 58294 507498 58350
rect 507554 58294 507622 58350
rect 507678 58294 525250 58350
rect 525306 58294 525374 58350
rect 525430 58294 525498 58350
rect 525554 58294 525622 58350
rect 525678 58294 543250 58350
rect 543306 58294 543374 58350
rect 543430 58294 543498 58350
rect 543554 58294 543622 58350
rect 543678 58294 561250 58350
rect 561306 58294 561374 58350
rect 561430 58294 561498 58350
rect 561554 58294 561622 58350
rect 561678 58294 579250 58350
rect 579306 58294 579374 58350
rect 579430 58294 579498 58350
rect 579554 58294 579622 58350
rect 579678 58294 596496 58350
rect 596552 58294 596620 58350
rect 596676 58294 596744 58350
rect 596800 58294 596868 58350
rect 596924 58294 597980 58350
rect -1916 58226 597980 58294
rect -1916 58170 -860 58226
rect -804 58170 -736 58226
rect -680 58170 -612 58226
rect -556 58170 -488 58226
rect -432 58170 3250 58226
rect 3306 58170 3374 58226
rect 3430 58170 3498 58226
rect 3554 58170 3622 58226
rect 3678 58170 21250 58226
rect 21306 58170 21374 58226
rect 21430 58170 21498 58226
rect 21554 58170 21622 58226
rect 21678 58170 39250 58226
rect 39306 58170 39374 58226
rect 39430 58170 39498 58226
rect 39554 58170 39622 58226
rect 39678 58170 57250 58226
rect 57306 58170 57374 58226
rect 57430 58170 57498 58226
rect 57554 58170 57622 58226
rect 57678 58170 75250 58226
rect 75306 58170 75374 58226
rect 75430 58170 75498 58226
rect 75554 58170 75622 58226
rect 75678 58170 93250 58226
rect 93306 58170 93374 58226
rect 93430 58170 93498 58226
rect 93554 58170 93622 58226
rect 93678 58170 111250 58226
rect 111306 58170 111374 58226
rect 111430 58170 111498 58226
rect 111554 58170 111622 58226
rect 111678 58170 129250 58226
rect 129306 58170 129374 58226
rect 129430 58170 129498 58226
rect 129554 58170 129622 58226
rect 129678 58170 147250 58226
rect 147306 58170 147374 58226
rect 147430 58170 147498 58226
rect 147554 58170 147622 58226
rect 147678 58170 165250 58226
rect 165306 58170 165374 58226
rect 165430 58170 165498 58226
rect 165554 58170 165622 58226
rect 165678 58170 183250 58226
rect 183306 58170 183374 58226
rect 183430 58170 183498 58226
rect 183554 58170 183622 58226
rect 183678 58170 201250 58226
rect 201306 58170 201374 58226
rect 201430 58170 201498 58226
rect 201554 58170 201622 58226
rect 201678 58170 381250 58226
rect 381306 58170 381374 58226
rect 381430 58170 381498 58226
rect 381554 58170 381622 58226
rect 381678 58170 399250 58226
rect 399306 58170 399374 58226
rect 399430 58170 399498 58226
rect 399554 58170 399622 58226
rect 399678 58170 417250 58226
rect 417306 58170 417374 58226
rect 417430 58170 417498 58226
rect 417554 58170 417622 58226
rect 417678 58170 435250 58226
rect 435306 58170 435374 58226
rect 435430 58170 435498 58226
rect 435554 58170 435622 58226
rect 435678 58170 453250 58226
rect 453306 58170 453374 58226
rect 453430 58170 453498 58226
rect 453554 58170 453622 58226
rect 453678 58170 471250 58226
rect 471306 58170 471374 58226
rect 471430 58170 471498 58226
rect 471554 58170 471622 58226
rect 471678 58170 489250 58226
rect 489306 58170 489374 58226
rect 489430 58170 489498 58226
rect 489554 58170 489622 58226
rect 489678 58170 507250 58226
rect 507306 58170 507374 58226
rect 507430 58170 507498 58226
rect 507554 58170 507622 58226
rect 507678 58170 525250 58226
rect 525306 58170 525374 58226
rect 525430 58170 525498 58226
rect 525554 58170 525622 58226
rect 525678 58170 543250 58226
rect 543306 58170 543374 58226
rect 543430 58170 543498 58226
rect 543554 58170 543622 58226
rect 543678 58170 561250 58226
rect 561306 58170 561374 58226
rect 561430 58170 561498 58226
rect 561554 58170 561622 58226
rect 561678 58170 579250 58226
rect 579306 58170 579374 58226
rect 579430 58170 579498 58226
rect 579554 58170 579622 58226
rect 579678 58170 596496 58226
rect 596552 58170 596620 58226
rect 596676 58170 596744 58226
rect 596800 58170 596868 58226
rect 596924 58170 597980 58226
rect -1916 58102 597980 58170
rect -1916 58046 -860 58102
rect -804 58046 -736 58102
rect -680 58046 -612 58102
rect -556 58046 -488 58102
rect -432 58046 3250 58102
rect 3306 58046 3374 58102
rect 3430 58046 3498 58102
rect 3554 58046 3622 58102
rect 3678 58046 21250 58102
rect 21306 58046 21374 58102
rect 21430 58046 21498 58102
rect 21554 58046 21622 58102
rect 21678 58046 39250 58102
rect 39306 58046 39374 58102
rect 39430 58046 39498 58102
rect 39554 58046 39622 58102
rect 39678 58046 57250 58102
rect 57306 58046 57374 58102
rect 57430 58046 57498 58102
rect 57554 58046 57622 58102
rect 57678 58046 75250 58102
rect 75306 58046 75374 58102
rect 75430 58046 75498 58102
rect 75554 58046 75622 58102
rect 75678 58046 93250 58102
rect 93306 58046 93374 58102
rect 93430 58046 93498 58102
rect 93554 58046 93622 58102
rect 93678 58046 111250 58102
rect 111306 58046 111374 58102
rect 111430 58046 111498 58102
rect 111554 58046 111622 58102
rect 111678 58046 129250 58102
rect 129306 58046 129374 58102
rect 129430 58046 129498 58102
rect 129554 58046 129622 58102
rect 129678 58046 147250 58102
rect 147306 58046 147374 58102
rect 147430 58046 147498 58102
rect 147554 58046 147622 58102
rect 147678 58046 165250 58102
rect 165306 58046 165374 58102
rect 165430 58046 165498 58102
rect 165554 58046 165622 58102
rect 165678 58046 183250 58102
rect 183306 58046 183374 58102
rect 183430 58046 183498 58102
rect 183554 58046 183622 58102
rect 183678 58046 201250 58102
rect 201306 58046 201374 58102
rect 201430 58046 201498 58102
rect 201554 58046 201622 58102
rect 201678 58046 381250 58102
rect 381306 58046 381374 58102
rect 381430 58046 381498 58102
rect 381554 58046 381622 58102
rect 381678 58046 399250 58102
rect 399306 58046 399374 58102
rect 399430 58046 399498 58102
rect 399554 58046 399622 58102
rect 399678 58046 417250 58102
rect 417306 58046 417374 58102
rect 417430 58046 417498 58102
rect 417554 58046 417622 58102
rect 417678 58046 435250 58102
rect 435306 58046 435374 58102
rect 435430 58046 435498 58102
rect 435554 58046 435622 58102
rect 435678 58046 453250 58102
rect 453306 58046 453374 58102
rect 453430 58046 453498 58102
rect 453554 58046 453622 58102
rect 453678 58046 471250 58102
rect 471306 58046 471374 58102
rect 471430 58046 471498 58102
rect 471554 58046 471622 58102
rect 471678 58046 489250 58102
rect 489306 58046 489374 58102
rect 489430 58046 489498 58102
rect 489554 58046 489622 58102
rect 489678 58046 507250 58102
rect 507306 58046 507374 58102
rect 507430 58046 507498 58102
rect 507554 58046 507622 58102
rect 507678 58046 525250 58102
rect 525306 58046 525374 58102
rect 525430 58046 525498 58102
rect 525554 58046 525622 58102
rect 525678 58046 543250 58102
rect 543306 58046 543374 58102
rect 543430 58046 543498 58102
rect 543554 58046 543622 58102
rect 543678 58046 561250 58102
rect 561306 58046 561374 58102
rect 561430 58046 561498 58102
rect 561554 58046 561622 58102
rect 561678 58046 579250 58102
rect 579306 58046 579374 58102
rect 579430 58046 579498 58102
rect 579554 58046 579622 58102
rect 579678 58046 596496 58102
rect 596552 58046 596620 58102
rect 596676 58046 596744 58102
rect 596800 58046 596868 58102
rect 596924 58046 597980 58102
rect -1916 57978 597980 58046
rect -1916 57922 -860 57978
rect -804 57922 -736 57978
rect -680 57922 -612 57978
rect -556 57922 -488 57978
rect -432 57922 3250 57978
rect 3306 57922 3374 57978
rect 3430 57922 3498 57978
rect 3554 57922 3622 57978
rect 3678 57922 21250 57978
rect 21306 57922 21374 57978
rect 21430 57922 21498 57978
rect 21554 57922 21622 57978
rect 21678 57922 39250 57978
rect 39306 57922 39374 57978
rect 39430 57922 39498 57978
rect 39554 57922 39622 57978
rect 39678 57922 57250 57978
rect 57306 57922 57374 57978
rect 57430 57922 57498 57978
rect 57554 57922 57622 57978
rect 57678 57922 75250 57978
rect 75306 57922 75374 57978
rect 75430 57922 75498 57978
rect 75554 57922 75622 57978
rect 75678 57922 93250 57978
rect 93306 57922 93374 57978
rect 93430 57922 93498 57978
rect 93554 57922 93622 57978
rect 93678 57922 111250 57978
rect 111306 57922 111374 57978
rect 111430 57922 111498 57978
rect 111554 57922 111622 57978
rect 111678 57922 129250 57978
rect 129306 57922 129374 57978
rect 129430 57922 129498 57978
rect 129554 57922 129622 57978
rect 129678 57922 147250 57978
rect 147306 57922 147374 57978
rect 147430 57922 147498 57978
rect 147554 57922 147622 57978
rect 147678 57922 165250 57978
rect 165306 57922 165374 57978
rect 165430 57922 165498 57978
rect 165554 57922 165622 57978
rect 165678 57922 183250 57978
rect 183306 57922 183374 57978
rect 183430 57922 183498 57978
rect 183554 57922 183622 57978
rect 183678 57922 201250 57978
rect 201306 57922 201374 57978
rect 201430 57922 201498 57978
rect 201554 57922 201622 57978
rect 201678 57922 381250 57978
rect 381306 57922 381374 57978
rect 381430 57922 381498 57978
rect 381554 57922 381622 57978
rect 381678 57922 399250 57978
rect 399306 57922 399374 57978
rect 399430 57922 399498 57978
rect 399554 57922 399622 57978
rect 399678 57922 417250 57978
rect 417306 57922 417374 57978
rect 417430 57922 417498 57978
rect 417554 57922 417622 57978
rect 417678 57922 435250 57978
rect 435306 57922 435374 57978
rect 435430 57922 435498 57978
rect 435554 57922 435622 57978
rect 435678 57922 453250 57978
rect 453306 57922 453374 57978
rect 453430 57922 453498 57978
rect 453554 57922 453622 57978
rect 453678 57922 471250 57978
rect 471306 57922 471374 57978
rect 471430 57922 471498 57978
rect 471554 57922 471622 57978
rect 471678 57922 489250 57978
rect 489306 57922 489374 57978
rect 489430 57922 489498 57978
rect 489554 57922 489622 57978
rect 489678 57922 507250 57978
rect 507306 57922 507374 57978
rect 507430 57922 507498 57978
rect 507554 57922 507622 57978
rect 507678 57922 525250 57978
rect 525306 57922 525374 57978
rect 525430 57922 525498 57978
rect 525554 57922 525622 57978
rect 525678 57922 543250 57978
rect 543306 57922 543374 57978
rect 543430 57922 543498 57978
rect 543554 57922 543622 57978
rect 543678 57922 561250 57978
rect 561306 57922 561374 57978
rect 561430 57922 561498 57978
rect 561554 57922 561622 57978
rect 561678 57922 579250 57978
rect 579306 57922 579374 57978
rect 579430 57922 579498 57978
rect 579554 57922 579622 57978
rect 579678 57922 596496 57978
rect 596552 57922 596620 57978
rect 596676 57922 596744 57978
rect 596800 57922 596868 57978
rect 596924 57922 597980 57978
rect -1916 57826 597980 57922
rect -1916 46350 597980 46446
rect -1916 46294 -1820 46350
rect -1764 46294 -1696 46350
rect -1640 46294 -1572 46350
rect -1516 46294 -1448 46350
rect -1392 46294 6970 46350
rect 7026 46294 7094 46350
rect 7150 46294 7218 46350
rect 7274 46294 7342 46350
rect 7398 46294 24970 46350
rect 25026 46294 25094 46350
rect 25150 46294 25218 46350
rect 25274 46294 25342 46350
rect 25398 46294 42970 46350
rect 43026 46294 43094 46350
rect 43150 46294 43218 46350
rect 43274 46294 43342 46350
rect 43398 46294 60970 46350
rect 61026 46294 61094 46350
rect 61150 46294 61218 46350
rect 61274 46294 61342 46350
rect 61398 46294 78970 46350
rect 79026 46294 79094 46350
rect 79150 46294 79218 46350
rect 79274 46294 79342 46350
rect 79398 46294 96970 46350
rect 97026 46294 97094 46350
rect 97150 46294 97218 46350
rect 97274 46294 97342 46350
rect 97398 46294 114970 46350
rect 115026 46294 115094 46350
rect 115150 46294 115218 46350
rect 115274 46294 115342 46350
rect 115398 46294 132970 46350
rect 133026 46294 133094 46350
rect 133150 46294 133218 46350
rect 133274 46294 133342 46350
rect 133398 46294 150970 46350
rect 151026 46294 151094 46350
rect 151150 46294 151218 46350
rect 151274 46294 151342 46350
rect 151398 46294 168970 46350
rect 169026 46294 169094 46350
rect 169150 46294 169218 46350
rect 169274 46294 169342 46350
rect 169398 46294 186970 46350
rect 187026 46294 187094 46350
rect 187150 46294 187218 46350
rect 187274 46294 187342 46350
rect 187398 46294 204970 46350
rect 205026 46294 205094 46350
rect 205150 46294 205218 46350
rect 205274 46294 205342 46350
rect 205398 46294 384970 46350
rect 385026 46294 385094 46350
rect 385150 46294 385218 46350
rect 385274 46294 385342 46350
rect 385398 46294 402970 46350
rect 403026 46294 403094 46350
rect 403150 46294 403218 46350
rect 403274 46294 403342 46350
rect 403398 46294 420970 46350
rect 421026 46294 421094 46350
rect 421150 46294 421218 46350
rect 421274 46294 421342 46350
rect 421398 46294 438970 46350
rect 439026 46294 439094 46350
rect 439150 46294 439218 46350
rect 439274 46294 439342 46350
rect 439398 46294 456970 46350
rect 457026 46294 457094 46350
rect 457150 46294 457218 46350
rect 457274 46294 457342 46350
rect 457398 46294 474970 46350
rect 475026 46294 475094 46350
rect 475150 46294 475218 46350
rect 475274 46294 475342 46350
rect 475398 46294 492970 46350
rect 493026 46294 493094 46350
rect 493150 46294 493218 46350
rect 493274 46294 493342 46350
rect 493398 46294 510970 46350
rect 511026 46294 511094 46350
rect 511150 46294 511218 46350
rect 511274 46294 511342 46350
rect 511398 46294 528970 46350
rect 529026 46294 529094 46350
rect 529150 46294 529218 46350
rect 529274 46294 529342 46350
rect 529398 46294 546970 46350
rect 547026 46294 547094 46350
rect 547150 46294 547218 46350
rect 547274 46294 547342 46350
rect 547398 46294 564970 46350
rect 565026 46294 565094 46350
rect 565150 46294 565218 46350
rect 565274 46294 565342 46350
rect 565398 46294 582970 46350
rect 583026 46294 583094 46350
rect 583150 46294 583218 46350
rect 583274 46294 583342 46350
rect 583398 46294 597456 46350
rect 597512 46294 597580 46350
rect 597636 46294 597704 46350
rect 597760 46294 597828 46350
rect 597884 46294 597980 46350
rect -1916 46226 597980 46294
rect -1916 46170 -1820 46226
rect -1764 46170 -1696 46226
rect -1640 46170 -1572 46226
rect -1516 46170 -1448 46226
rect -1392 46170 6970 46226
rect 7026 46170 7094 46226
rect 7150 46170 7218 46226
rect 7274 46170 7342 46226
rect 7398 46170 24970 46226
rect 25026 46170 25094 46226
rect 25150 46170 25218 46226
rect 25274 46170 25342 46226
rect 25398 46170 42970 46226
rect 43026 46170 43094 46226
rect 43150 46170 43218 46226
rect 43274 46170 43342 46226
rect 43398 46170 60970 46226
rect 61026 46170 61094 46226
rect 61150 46170 61218 46226
rect 61274 46170 61342 46226
rect 61398 46170 78970 46226
rect 79026 46170 79094 46226
rect 79150 46170 79218 46226
rect 79274 46170 79342 46226
rect 79398 46170 96970 46226
rect 97026 46170 97094 46226
rect 97150 46170 97218 46226
rect 97274 46170 97342 46226
rect 97398 46170 114970 46226
rect 115026 46170 115094 46226
rect 115150 46170 115218 46226
rect 115274 46170 115342 46226
rect 115398 46170 132970 46226
rect 133026 46170 133094 46226
rect 133150 46170 133218 46226
rect 133274 46170 133342 46226
rect 133398 46170 150970 46226
rect 151026 46170 151094 46226
rect 151150 46170 151218 46226
rect 151274 46170 151342 46226
rect 151398 46170 168970 46226
rect 169026 46170 169094 46226
rect 169150 46170 169218 46226
rect 169274 46170 169342 46226
rect 169398 46170 186970 46226
rect 187026 46170 187094 46226
rect 187150 46170 187218 46226
rect 187274 46170 187342 46226
rect 187398 46170 204970 46226
rect 205026 46170 205094 46226
rect 205150 46170 205218 46226
rect 205274 46170 205342 46226
rect 205398 46170 384970 46226
rect 385026 46170 385094 46226
rect 385150 46170 385218 46226
rect 385274 46170 385342 46226
rect 385398 46170 402970 46226
rect 403026 46170 403094 46226
rect 403150 46170 403218 46226
rect 403274 46170 403342 46226
rect 403398 46170 420970 46226
rect 421026 46170 421094 46226
rect 421150 46170 421218 46226
rect 421274 46170 421342 46226
rect 421398 46170 438970 46226
rect 439026 46170 439094 46226
rect 439150 46170 439218 46226
rect 439274 46170 439342 46226
rect 439398 46170 456970 46226
rect 457026 46170 457094 46226
rect 457150 46170 457218 46226
rect 457274 46170 457342 46226
rect 457398 46170 474970 46226
rect 475026 46170 475094 46226
rect 475150 46170 475218 46226
rect 475274 46170 475342 46226
rect 475398 46170 492970 46226
rect 493026 46170 493094 46226
rect 493150 46170 493218 46226
rect 493274 46170 493342 46226
rect 493398 46170 510970 46226
rect 511026 46170 511094 46226
rect 511150 46170 511218 46226
rect 511274 46170 511342 46226
rect 511398 46170 528970 46226
rect 529026 46170 529094 46226
rect 529150 46170 529218 46226
rect 529274 46170 529342 46226
rect 529398 46170 546970 46226
rect 547026 46170 547094 46226
rect 547150 46170 547218 46226
rect 547274 46170 547342 46226
rect 547398 46170 564970 46226
rect 565026 46170 565094 46226
rect 565150 46170 565218 46226
rect 565274 46170 565342 46226
rect 565398 46170 582970 46226
rect 583026 46170 583094 46226
rect 583150 46170 583218 46226
rect 583274 46170 583342 46226
rect 583398 46170 597456 46226
rect 597512 46170 597580 46226
rect 597636 46170 597704 46226
rect 597760 46170 597828 46226
rect 597884 46170 597980 46226
rect -1916 46102 597980 46170
rect -1916 46046 -1820 46102
rect -1764 46046 -1696 46102
rect -1640 46046 -1572 46102
rect -1516 46046 -1448 46102
rect -1392 46046 6970 46102
rect 7026 46046 7094 46102
rect 7150 46046 7218 46102
rect 7274 46046 7342 46102
rect 7398 46046 24970 46102
rect 25026 46046 25094 46102
rect 25150 46046 25218 46102
rect 25274 46046 25342 46102
rect 25398 46046 42970 46102
rect 43026 46046 43094 46102
rect 43150 46046 43218 46102
rect 43274 46046 43342 46102
rect 43398 46046 60970 46102
rect 61026 46046 61094 46102
rect 61150 46046 61218 46102
rect 61274 46046 61342 46102
rect 61398 46046 78970 46102
rect 79026 46046 79094 46102
rect 79150 46046 79218 46102
rect 79274 46046 79342 46102
rect 79398 46046 96970 46102
rect 97026 46046 97094 46102
rect 97150 46046 97218 46102
rect 97274 46046 97342 46102
rect 97398 46046 114970 46102
rect 115026 46046 115094 46102
rect 115150 46046 115218 46102
rect 115274 46046 115342 46102
rect 115398 46046 132970 46102
rect 133026 46046 133094 46102
rect 133150 46046 133218 46102
rect 133274 46046 133342 46102
rect 133398 46046 150970 46102
rect 151026 46046 151094 46102
rect 151150 46046 151218 46102
rect 151274 46046 151342 46102
rect 151398 46046 168970 46102
rect 169026 46046 169094 46102
rect 169150 46046 169218 46102
rect 169274 46046 169342 46102
rect 169398 46046 186970 46102
rect 187026 46046 187094 46102
rect 187150 46046 187218 46102
rect 187274 46046 187342 46102
rect 187398 46046 204970 46102
rect 205026 46046 205094 46102
rect 205150 46046 205218 46102
rect 205274 46046 205342 46102
rect 205398 46046 384970 46102
rect 385026 46046 385094 46102
rect 385150 46046 385218 46102
rect 385274 46046 385342 46102
rect 385398 46046 402970 46102
rect 403026 46046 403094 46102
rect 403150 46046 403218 46102
rect 403274 46046 403342 46102
rect 403398 46046 420970 46102
rect 421026 46046 421094 46102
rect 421150 46046 421218 46102
rect 421274 46046 421342 46102
rect 421398 46046 438970 46102
rect 439026 46046 439094 46102
rect 439150 46046 439218 46102
rect 439274 46046 439342 46102
rect 439398 46046 456970 46102
rect 457026 46046 457094 46102
rect 457150 46046 457218 46102
rect 457274 46046 457342 46102
rect 457398 46046 474970 46102
rect 475026 46046 475094 46102
rect 475150 46046 475218 46102
rect 475274 46046 475342 46102
rect 475398 46046 492970 46102
rect 493026 46046 493094 46102
rect 493150 46046 493218 46102
rect 493274 46046 493342 46102
rect 493398 46046 510970 46102
rect 511026 46046 511094 46102
rect 511150 46046 511218 46102
rect 511274 46046 511342 46102
rect 511398 46046 528970 46102
rect 529026 46046 529094 46102
rect 529150 46046 529218 46102
rect 529274 46046 529342 46102
rect 529398 46046 546970 46102
rect 547026 46046 547094 46102
rect 547150 46046 547218 46102
rect 547274 46046 547342 46102
rect 547398 46046 564970 46102
rect 565026 46046 565094 46102
rect 565150 46046 565218 46102
rect 565274 46046 565342 46102
rect 565398 46046 582970 46102
rect 583026 46046 583094 46102
rect 583150 46046 583218 46102
rect 583274 46046 583342 46102
rect 583398 46046 597456 46102
rect 597512 46046 597580 46102
rect 597636 46046 597704 46102
rect 597760 46046 597828 46102
rect 597884 46046 597980 46102
rect -1916 45978 597980 46046
rect -1916 45922 -1820 45978
rect -1764 45922 -1696 45978
rect -1640 45922 -1572 45978
rect -1516 45922 -1448 45978
rect -1392 45922 6970 45978
rect 7026 45922 7094 45978
rect 7150 45922 7218 45978
rect 7274 45922 7342 45978
rect 7398 45922 24970 45978
rect 25026 45922 25094 45978
rect 25150 45922 25218 45978
rect 25274 45922 25342 45978
rect 25398 45922 42970 45978
rect 43026 45922 43094 45978
rect 43150 45922 43218 45978
rect 43274 45922 43342 45978
rect 43398 45922 60970 45978
rect 61026 45922 61094 45978
rect 61150 45922 61218 45978
rect 61274 45922 61342 45978
rect 61398 45922 78970 45978
rect 79026 45922 79094 45978
rect 79150 45922 79218 45978
rect 79274 45922 79342 45978
rect 79398 45922 96970 45978
rect 97026 45922 97094 45978
rect 97150 45922 97218 45978
rect 97274 45922 97342 45978
rect 97398 45922 114970 45978
rect 115026 45922 115094 45978
rect 115150 45922 115218 45978
rect 115274 45922 115342 45978
rect 115398 45922 132970 45978
rect 133026 45922 133094 45978
rect 133150 45922 133218 45978
rect 133274 45922 133342 45978
rect 133398 45922 150970 45978
rect 151026 45922 151094 45978
rect 151150 45922 151218 45978
rect 151274 45922 151342 45978
rect 151398 45922 168970 45978
rect 169026 45922 169094 45978
rect 169150 45922 169218 45978
rect 169274 45922 169342 45978
rect 169398 45922 186970 45978
rect 187026 45922 187094 45978
rect 187150 45922 187218 45978
rect 187274 45922 187342 45978
rect 187398 45922 204970 45978
rect 205026 45922 205094 45978
rect 205150 45922 205218 45978
rect 205274 45922 205342 45978
rect 205398 45922 384970 45978
rect 385026 45922 385094 45978
rect 385150 45922 385218 45978
rect 385274 45922 385342 45978
rect 385398 45922 402970 45978
rect 403026 45922 403094 45978
rect 403150 45922 403218 45978
rect 403274 45922 403342 45978
rect 403398 45922 420970 45978
rect 421026 45922 421094 45978
rect 421150 45922 421218 45978
rect 421274 45922 421342 45978
rect 421398 45922 438970 45978
rect 439026 45922 439094 45978
rect 439150 45922 439218 45978
rect 439274 45922 439342 45978
rect 439398 45922 456970 45978
rect 457026 45922 457094 45978
rect 457150 45922 457218 45978
rect 457274 45922 457342 45978
rect 457398 45922 474970 45978
rect 475026 45922 475094 45978
rect 475150 45922 475218 45978
rect 475274 45922 475342 45978
rect 475398 45922 492970 45978
rect 493026 45922 493094 45978
rect 493150 45922 493218 45978
rect 493274 45922 493342 45978
rect 493398 45922 510970 45978
rect 511026 45922 511094 45978
rect 511150 45922 511218 45978
rect 511274 45922 511342 45978
rect 511398 45922 528970 45978
rect 529026 45922 529094 45978
rect 529150 45922 529218 45978
rect 529274 45922 529342 45978
rect 529398 45922 546970 45978
rect 547026 45922 547094 45978
rect 547150 45922 547218 45978
rect 547274 45922 547342 45978
rect 547398 45922 564970 45978
rect 565026 45922 565094 45978
rect 565150 45922 565218 45978
rect 565274 45922 565342 45978
rect 565398 45922 582970 45978
rect 583026 45922 583094 45978
rect 583150 45922 583218 45978
rect 583274 45922 583342 45978
rect 583398 45922 597456 45978
rect 597512 45922 597580 45978
rect 597636 45922 597704 45978
rect 597760 45922 597828 45978
rect 597884 45922 597980 45978
rect -1916 45826 597980 45922
rect -1916 40350 597980 40446
rect -1916 40294 -860 40350
rect -804 40294 -736 40350
rect -680 40294 -612 40350
rect -556 40294 -488 40350
rect -432 40294 3250 40350
rect 3306 40294 3374 40350
rect 3430 40294 3498 40350
rect 3554 40294 3622 40350
rect 3678 40294 21250 40350
rect 21306 40294 21374 40350
rect 21430 40294 21498 40350
rect 21554 40294 21622 40350
rect 21678 40294 39250 40350
rect 39306 40294 39374 40350
rect 39430 40294 39498 40350
rect 39554 40294 39622 40350
rect 39678 40294 57250 40350
rect 57306 40294 57374 40350
rect 57430 40294 57498 40350
rect 57554 40294 57622 40350
rect 57678 40294 75250 40350
rect 75306 40294 75374 40350
rect 75430 40294 75498 40350
rect 75554 40294 75622 40350
rect 75678 40294 93250 40350
rect 93306 40294 93374 40350
rect 93430 40294 93498 40350
rect 93554 40294 93622 40350
rect 93678 40294 111250 40350
rect 111306 40294 111374 40350
rect 111430 40294 111498 40350
rect 111554 40294 111622 40350
rect 111678 40294 129250 40350
rect 129306 40294 129374 40350
rect 129430 40294 129498 40350
rect 129554 40294 129622 40350
rect 129678 40294 147250 40350
rect 147306 40294 147374 40350
rect 147430 40294 147498 40350
rect 147554 40294 147622 40350
rect 147678 40294 165250 40350
rect 165306 40294 165374 40350
rect 165430 40294 165498 40350
rect 165554 40294 165622 40350
rect 165678 40294 183250 40350
rect 183306 40294 183374 40350
rect 183430 40294 183498 40350
rect 183554 40294 183622 40350
rect 183678 40294 201250 40350
rect 201306 40294 201374 40350
rect 201430 40294 201498 40350
rect 201554 40294 201622 40350
rect 201678 40294 381250 40350
rect 381306 40294 381374 40350
rect 381430 40294 381498 40350
rect 381554 40294 381622 40350
rect 381678 40294 399250 40350
rect 399306 40294 399374 40350
rect 399430 40294 399498 40350
rect 399554 40294 399622 40350
rect 399678 40294 417250 40350
rect 417306 40294 417374 40350
rect 417430 40294 417498 40350
rect 417554 40294 417622 40350
rect 417678 40294 435250 40350
rect 435306 40294 435374 40350
rect 435430 40294 435498 40350
rect 435554 40294 435622 40350
rect 435678 40294 453250 40350
rect 453306 40294 453374 40350
rect 453430 40294 453498 40350
rect 453554 40294 453622 40350
rect 453678 40294 471250 40350
rect 471306 40294 471374 40350
rect 471430 40294 471498 40350
rect 471554 40294 471622 40350
rect 471678 40294 489250 40350
rect 489306 40294 489374 40350
rect 489430 40294 489498 40350
rect 489554 40294 489622 40350
rect 489678 40294 507250 40350
rect 507306 40294 507374 40350
rect 507430 40294 507498 40350
rect 507554 40294 507622 40350
rect 507678 40294 525250 40350
rect 525306 40294 525374 40350
rect 525430 40294 525498 40350
rect 525554 40294 525622 40350
rect 525678 40294 543250 40350
rect 543306 40294 543374 40350
rect 543430 40294 543498 40350
rect 543554 40294 543622 40350
rect 543678 40294 561250 40350
rect 561306 40294 561374 40350
rect 561430 40294 561498 40350
rect 561554 40294 561622 40350
rect 561678 40294 579250 40350
rect 579306 40294 579374 40350
rect 579430 40294 579498 40350
rect 579554 40294 579622 40350
rect 579678 40294 596496 40350
rect 596552 40294 596620 40350
rect 596676 40294 596744 40350
rect 596800 40294 596868 40350
rect 596924 40294 597980 40350
rect -1916 40226 597980 40294
rect -1916 40170 -860 40226
rect -804 40170 -736 40226
rect -680 40170 -612 40226
rect -556 40170 -488 40226
rect -432 40170 3250 40226
rect 3306 40170 3374 40226
rect 3430 40170 3498 40226
rect 3554 40170 3622 40226
rect 3678 40170 21250 40226
rect 21306 40170 21374 40226
rect 21430 40170 21498 40226
rect 21554 40170 21622 40226
rect 21678 40170 39250 40226
rect 39306 40170 39374 40226
rect 39430 40170 39498 40226
rect 39554 40170 39622 40226
rect 39678 40170 57250 40226
rect 57306 40170 57374 40226
rect 57430 40170 57498 40226
rect 57554 40170 57622 40226
rect 57678 40170 75250 40226
rect 75306 40170 75374 40226
rect 75430 40170 75498 40226
rect 75554 40170 75622 40226
rect 75678 40170 93250 40226
rect 93306 40170 93374 40226
rect 93430 40170 93498 40226
rect 93554 40170 93622 40226
rect 93678 40170 111250 40226
rect 111306 40170 111374 40226
rect 111430 40170 111498 40226
rect 111554 40170 111622 40226
rect 111678 40170 129250 40226
rect 129306 40170 129374 40226
rect 129430 40170 129498 40226
rect 129554 40170 129622 40226
rect 129678 40170 147250 40226
rect 147306 40170 147374 40226
rect 147430 40170 147498 40226
rect 147554 40170 147622 40226
rect 147678 40170 165250 40226
rect 165306 40170 165374 40226
rect 165430 40170 165498 40226
rect 165554 40170 165622 40226
rect 165678 40170 183250 40226
rect 183306 40170 183374 40226
rect 183430 40170 183498 40226
rect 183554 40170 183622 40226
rect 183678 40170 201250 40226
rect 201306 40170 201374 40226
rect 201430 40170 201498 40226
rect 201554 40170 201622 40226
rect 201678 40170 381250 40226
rect 381306 40170 381374 40226
rect 381430 40170 381498 40226
rect 381554 40170 381622 40226
rect 381678 40170 399250 40226
rect 399306 40170 399374 40226
rect 399430 40170 399498 40226
rect 399554 40170 399622 40226
rect 399678 40170 417250 40226
rect 417306 40170 417374 40226
rect 417430 40170 417498 40226
rect 417554 40170 417622 40226
rect 417678 40170 435250 40226
rect 435306 40170 435374 40226
rect 435430 40170 435498 40226
rect 435554 40170 435622 40226
rect 435678 40170 453250 40226
rect 453306 40170 453374 40226
rect 453430 40170 453498 40226
rect 453554 40170 453622 40226
rect 453678 40170 471250 40226
rect 471306 40170 471374 40226
rect 471430 40170 471498 40226
rect 471554 40170 471622 40226
rect 471678 40170 489250 40226
rect 489306 40170 489374 40226
rect 489430 40170 489498 40226
rect 489554 40170 489622 40226
rect 489678 40170 507250 40226
rect 507306 40170 507374 40226
rect 507430 40170 507498 40226
rect 507554 40170 507622 40226
rect 507678 40170 525250 40226
rect 525306 40170 525374 40226
rect 525430 40170 525498 40226
rect 525554 40170 525622 40226
rect 525678 40170 543250 40226
rect 543306 40170 543374 40226
rect 543430 40170 543498 40226
rect 543554 40170 543622 40226
rect 543678 40170 561250 40226
rect 561306 40170 561374 40226
rect 561430 40170 561498 40226
rect 561554 40170 561622 40226
rect 561678 40170 579250 40226
rect 579306 40170 579374 40226
rect 579430 40170 579498 40226
rect 579554 40170 579622 40226
rect 579678 40170 596496 40226
rect 596552 40170 596620 40226
rect 596676 40170 596744 40226
rect 596800 40170 596868 40226
rect 596924 40170 597980 40226
rect -1916 40102 597980 40170
rect -1916 40046 -860 40102
rect -804 40046 -736 40102
rect -680 40046 -612 40102
rect -556 40046 -488 40102
rect -432 40046 3250 40102
rect 3306 40046 3374 40102
rect 3430 40046 3498 40102
rect 3554 40046 3622 40102
rect 3678 40046 21250 40102
rect 21306 40046 21374 40102
rect 21430 40046 21498 40102
rect 21554 40046 21622 40102
rect 21678 40046 39250 40102
rect 39306 40046 39374 40102
rect 39430 40046 39498 40102
rect 39554 40046 39622 40102
rect 39678 40046 57250 40102
rect 57306 40046 57374 40102
rect 57430 40046 57498 40102
rect 57554 40046 57622 40102
rect 57678 40046 75250 40102
rect 75306 40046 75374 40102
rect 75430 40046 75498 40102
rect 75554 40046 75622 40102
rect 75678 40046 93250 40102
rect 93306 40046 93374 40102
rect 93430 40046 93498 40102
rect 93554 40046 93622 40102
rect 93678 40046 111250 40102
rect 111306 40046 111374 40102
rect 111430 40046 111498 40102
rect 111554 40046 111622 40102
rect 111678 40046 129250 40102
rect 129306 40046 129374 40102
rect 129430 40046 129498 40102
rect 129554 40046 129622 40102
rect 129678 40046 147250 40102
rect 147306 40046 147374 40102
rect 147430 40046 147498 40102
rect 147554 40046 147622 40102
rect 147678 40046 165250 40102
rect 165306 40046 165374 40102
rect 165430 40046 165498 40102
rect 165554 40046 165622 40102
rect 165678 40046 183250 40102
rect 183306 40046 183374 40102
rect 183430 40046 183498 40102
rect 183554 40046 183622 40102
rect 183678 40046 201250 40102
rect 201306 40046 201374 40102
rect 201430 40046 201498 40102
rect 201554 40046 201622 40102
rect 201678 40046 381250 40102
rect 381306 40046 381374 40102
rect 381430 40046 381498 40102
rect 381554 40046 381622 40102
rect 381678 40046 399250 40102
rect 399306 40046 399374 40102
rect 399430 40046 399498 40102
rect 399554 40046 399622 40102
rect 399678 40046 417250 40102
rect 417306 40046 417374 40102
rect 417430 40046 417498 40102
rect 417554 40046 417622 40102
rect 417678 40046 435250 40102
rect 435306 40046 435374 40102
rect 435430 40046 435498 40102
rect 435554 40046 435622 40102
rect 435678 40046 453250 40102
rect 453306 40046 453374 40102
rect 453430 40046 453498 40102
rect 453554 40046 453622 40102
rect 453678 40046 471250 40102
rect 471306 40046 471374 40102
rect 471430 40046 471498 40102
rect 471554 40046 471622 40102
rect 471678 40046 489250 40102
rect 489306 40046 489374 40102
rect 489430 40046 489498 40102
rect 489554 40046 489622 40102
rect 489678 40046 507250 40102
rect 507306 40046 507374 40102
rect 507430 40046 507498 40102
rect 507554 40046 507622 40102
rect 507678 40046 525250 40102
rect 525306 40046 525374 40102
rect 525430 40046 525498 40102
rect 525554 40046 525622 40102
rect 525678 40046 543250 40102
rect 543306 40046 543374 40102
rect 543430 40046 543498 40102
rect 543554 40046 543622 40102
rect 543678 40046 561250 40102
rect 561306 40046 561374 40102
rect 561430 40046 561498 40102
rect 561554 40046 561622 40102
rect 561678 40046 579250 40102
rect 579306 40046 579374 40102
rect 579430 40046 579498 40102
rect 579554 40046 579622 40102
rect 579678 40046 596496 40102
rect 596552 40046 596620 40102
rect 596676 40046 596744 40102
rect 596800 40046 596868 40102
rect 596924 40046 597980 40102
rect -1916 39978 597980 40046
rect -1916 39922 -860 39978
rect -804 39922 -736 39978
rect -680 39922 -612 39978
rect -556 39922 -488 39978
rect -432 39922 3250 39978
rect 3306 39922 3374 39978
rect 3430 39922 3498 39978
rect 3554 39922 3622 39978
rect 3678 39922 21250 39978
rect 21306 39922 21374 39978
rect 21430 39922 21498 39978
rect 21554 39922 21622 39978
rect 21678 39922 39250 39978
rect 39306 39922 39374 39978
rect 39430 39922 39498 39978
rect 39554 39922 39622 39978
rect 39678 39922 57250 39978
rect 57306 39922 57374 39978
rect 57430 39922 57498 39978
rect 57554 39922 57622 39978
rect 57678 39922 75250 39978
rect 75306 39922 75374 39978
rect 75430 39922 75498 39978
rect 75554 39922 75622 39978
rect 75678 39922 93250 39978
rect 93306 39922 93374 39978
rect 93430 39922 93498 39978
rect 93554 39922 93622 39978
rect 93678 39922 111250 39978
rect 111306 39922 111374 39978
rect 111430 39922 111498 39978
rect 111554 39922 111622 39978
rect 111678 39922 129250 39978
rect 129306 39922 129374 39978
rect 129430 39922 129498 39978
rect 129554 39922 129622 39978
rect 129678 39922 147250 39978
rect 147306 39922 147374 39978
rect 147430 39922 147498 39978
rect 147554 39922 147622 39978
rect 147678 39922 165250 39978
rect 165306 39922 165374 39978
rect 165430 39922 165498 39978
rect 165554 39922 165622 39978
rect 165678 39922 183250 39978
rect 183306 39922 183374 39978
rect 183430 39922 183498 39978
rect 183554 39922 183622 39978
rect 183678 39922 201250 39978
rect 201306 39922 201374 39978
rect 201430 39922 201498 39978
rect 201554 39922 201622 39978
rect 201678 39922 381250 39978
rect 381306 39922 381374 39978
rect 381430 39922 381498 39978
rect 381554 39922 381622 39978
rect 381678 39922 399250 39978
rect 399306 39922 399374 39978
rect 399430 39922 399498 39978
rect 399554 39922 399622 39978
rect 399678 39922 417250 39978
rect 417306 39922 417374 39978
rect 417430 39922 417498 39978
rect 417554 39922 417622 39978
rect 417678 39922 435250 39978
rect 435306 39922 435374 39978
rect 435430 39922 435498 39978
rect 435554 39922 435622 39978
rect 435678 39922 453250 39978
rect 453306 39922 453374 39978
rect 453430 39922 453498 39978
rect 453554 39922 453622 39978
rect 453678 39922 471250 39978
rect 471306 39922 471374 39978
rect 471430 39922 471498 39978
rect 471554 39922 471622 39978
rect 471678 39922 489250 39978
rect 489306 39922 489374 39978
rect 489430 39922 489498 39978
rect 489554 39922 489622 39978
rect 489678 39922 507250 39978
rect 507306 39922 507374 39978
rect 507430 39922 507498 39978
rect 507554 39922 507622 39978
rect 507678 39922 525250 39978
rect 525306 39922 525374 39978
rect 525430 39922 525498 39978
rect 525554 39922 525622 39978
rect 525678 39922 543250 39978
rect 543306 39922 543374 39978
rect 543430 39922 543498 39978
rect 543554 39922 543622 39978
rect 543678 39922 561250 39978
rect 561306 39922 561374 39978
rect 561430 39922 561498 39978
rect 561554 39922 561622 39978
rect 561678 39922 579250 39978
rect 579306 39922 579374 39978
rect 579430 39922 579498 39978
rect 579554 39922 579622 39978
rect 579678 39922 596496 39978
rect 596552 39922 596620 39978
rect 596676 39922 596744 39978
rect 596800 39922 596868 39978
rect 596924 39922 597980 39978
rect -1916 39826 597980 39922
rect -1916 28350 597980 28446
rect -1916 28294 -1820 28350
rect -1764 28294 -1696 28350
rect -1640 28294 -1572 28350
rect -1516 28294 -1448 28350
rect -1392 28294 6970 28350
rect 7026 28294 7094 28350
rect 7150 28294 7218 28350
rect 7274 28294 7342 28350
rect 7398 28294 24970 28350
rect 25026 28294 25094 28350
rect 25150 28294 25218 28350
rect 25274 28294 25342 28350
rect 25398 28294 42970 28350
rect 43026 28294 43094 28350
rect 43150 28294 43218 28350
rect 43274 28294 43342 28350
rect 43398 28294 60970 28350
rect 61026 28294 61094 28350
rect 61150 28294 61218 28350
rect 61274 28294 61342 28350
rect 61398 28294 78970 28350
rect 79026 28294 79094 28350
rect 79150 28294 79218 28350
rect 79274 28294 79342 28350
rect 79398 28294 96970 28350
rect 97026 28294 97094 28350
rect 97150 28294 97218 28350
rect 97274 28294 97342 28350
rect 97398 28294 114970 28350
rect 115026 28294 115094 28350
rect 115150 28294 115218 28350
rect 115274 28294 115342 28350
rect 115398 28294 132970 28350
rect 133026 28294 133094 28350
rect 133150 28294 133218 28350
rect 133274 28294 133342 28350
rect 133398 28294 150970 28350
rect 151026 28294 151094 28350
rect 151150 28294 151218 28350
rect 151274 28294 151342 28350
rect 151398 28294 168970 28350
rect 169026 28294 169094 28350
rect 169150 28294 169218 28350
rect 169274 28294 169342 28350
rect 169398 28294 186970 28350
rect 187026 28294 187094 28350
rect 187150 28294 187218 28350
rect 187274 28294 187342 28350
rect 187398 28294 204970 28350
rect 205026 28294 205094 28350
rect 205150 28294 205218 28350
rect 205274 28294 205342 28350
rect 205398 28294 384970 28350
rect 385026 28294 385094 28350
rect 385150 28294 385218 28350
rect 385274 28294 385342 28350
rect 385398 28294 402970 28350
rect 403026 28294 403094 28350
rect 403150 28294 403218 28350
rect 403274 28294 403342 28350
rect 403398 28294 420970 28350
rect 421026 28294 421094 28350
rect 421150 28294 421218 28350
rect 421274 28294 421342 28350
rect 421398 28294 438970 28350
rect 439026 28294 439094 28350
rect 439150 28294 439218 28350
rect 439274 28294 439342 28350
rect 439398 28294 456970 28350
rect 457026 28294 457094 28350
rect 457150 28294 457218 28350
rect 457274 28294 457342 28350
rect 457398 28294 474970 28350
rect 475026 28294 475094 28350
rect 475150 28294 475218 28350
rect 475274 28294 475342 28350
rect 475398 28294 492970 28350
rect 493026 28294 493094 28350
rect 493150 28294 493218 28350
rect 493274 28294 493342 28350
rect 493398 28294 510970 28350
rect 511026 28294 511094 28350
rect 511150 28294 511218 28350
rect 511274 28294 511342 28350
rect 511398 28294 528970 28350
rect 529026 28294 529094 28350
rect 529150 28294 529218 28350
rect 529274 28294 529342 28350
rect 529398 28294 546970 28350
rect 547026 28294 547094 28350
rect 547150 28294 547218 28350
rect 547274 28294 547342 28350
rect 547398 28294 564970 28350
rect 565026 28294 565094 28350
rect 565150 28294 565218 28350
rect 565274 28294 565342 28350
rect 565398 28294 582970 28350
rect 583026 28294 583094 28350
rect 583150 28294 583218 28350
rect 583274 28294 583342 28350
rect 583398 28294 597456 28350
rect 597512 28294 597580 28350
rect 597636 28294 597704 28350
rect 597760 28294 597828 28350
rect 597884 28294 597980 28350
rect -1916 28226 597980 28294
rect -1916 28170 -1820 28226
rect -1764 28170 -1696 28226
rect -1640 28170 -1572 28226
rect -1516 28170 -1448 28226
rect -1392 28170 6970 28226
rect 7026 28170 7094 28226
rect 7150 28170 7218 28226
rect 7274 28170 7342 28226
rect 7398 28170 24970 28226
rect 25026 28170 25094 28226
rect 25150 28170 25218 28226
rect 25274 28170 25342 28226
rect 25398 28170 42970 28226
rect 43026 28170 43094 28226
rect 43150 28170 43218 28226
rect 43274 28170 43342 28226
rect 43398 28170 60970 28226
rect 61026 28170 61094 28226
rect 61150 28170 61218 28226
rect 61274 28170 61342 28226
rect 61398 28170 78970 28226
rect 79026 28170 79094 28226
rect 79150 28170 79218 28226
rect 79274 28170 79342 28226
rect 79398 28170 96970 28226
rect 97026 28170 97094 28226
rect 97150 28170 97218 28226
rect 97274 28170 97342 28226
rect 97398 28170 114970 28226
rect 115026 28170 115094 28226
rect 115150 28170 115218 28226
rect 115274 28170 115342 28226
rect 115398 28170 132970 28226
rect 133026 28170 133094 28226
rect 133150 28170 133218 28226
rect 133274 28170 133342 28226
rect 133398 28170 150970 28226
rect 151026 28170 151094 28226
rect 151150 28170 151218 28226
rect 151274 28170 151342 28226
rect 151398 28170 168970 28226
rect 169026 28170 169094 28226
rect 169150 28170 169218 28226
rect 169274 28170 169342 28226
rect 169398 28170 186970 28226
rect 187026 28170 187094 28226
rect 187150 28170 187218 28226
rect 187274 28170 187342 28226
rect 187398 28170 204970 28226
rect 205026 28170 205094 28226
rect 205150 28170 205218 28226
rect 205274 28170 205342 28226
rect 205398 28170 384970 28226
rect 385026 28170 385094 28226
rect 385150 28170 385218 28226
rect 385274 28170 385342 28226
rect 385398 28170 402970 28226
rect 403026 28170 403094 28226
rect 403150 28170 403218 28226
rect 403274 28170 403342 28226
rect 403398 28170 420970 28226
rect 421026 28170 421094 28226
rect 421150 28170 421218 28226
rect 421274 28170 421342 28226
rect 421398 28170 438970 28226
rect 439026 28170 439094 28226
rect 439150 28170 439218 28226
rect 439274 28170 439342 28226
rect 439398 28170 456970 28226
rect 457026 28170 457094 28226
rect 457150 28170 457218 28226
rect 457274 28170 457342 28226
rect 457398 28170 474970 28226
rect 475026 28170 475094 28226
rect 475150 28170 475218 28226
rect 475274 28170 475342 28226
rect 475398 28170 492970 28226
rect 493026 28170 493094 28226
rect 493150 28170 493218 28226
rect 493274 28170 493342 28226
rect 493398 28170 510970 28226
rect 511026 28170 511094 28226
rect 511150 28170 511218 28226
rect 511274 28170 511342 28226
rect 511398 28170 528970 28226
rect 529026 28170 529094 28226
rect 529150 28170 529218 28226
rect 529274 28170 529342 28226
rect 529398 28170 546970 28226
rect 547026 28170 547094 28226
rect 547150 28170 547218 28226
rect 547274 28170 547342 28226
rect 547398 28170 564970 28226
rect 565026 28170 565094 28226
rect 565150 28170 565218 28226
rect 565274 28170 565342 28226
rect 565398 28170 582970 28226
rect 583026 28170 583094 28226
rect 583150 28170 583218 28226
rect 583274 28170 583342 28226
rect 583398 28170 597456 28226
rect 597512 28170 597580 28226
rect 597636 28170 597704 28226
rect 597760 28170 597828 28226
rect 597884 28170 597980 28226
rect -1916 28102 597980 28170
rect -1916 28046 -1820 28102
rect -1764 28046 -1696 28102
rect -1640 28046 -1572 28102
rect -1516 28046 -1448 28102
rect -1392 28046 6970 28102
rect 7026 28046 7094 28102
rect 7150 28046 7218 28102
rect 7274 28046 7342 28102
rect 7398 28046 24970 28102
rect 25026 28046 25094 28102
rect 25150 28046 25218 28102
rect 25274 28046 25342 28102
rect 25398 28046 42970 28102
rect 43026 28046 43094 28102
rect 43150 28046 43218 28102
rect 43274 28046 43342 28102
rect 43398 28046 60970 28102
rect 61026 28046 61094 28102
rect 61150 28046 61218 28102
rect 61274 28046 61342 28102
rect 61398 28046 78970 28102
rect 79026 28046 79094 28102
rect 79150 28046 79218 28102
rect 79274 28046 79342 28102
rect 79398 28046 96970 28102
rect 97026 28046 97094 28102
rect 97150 28046 97218 28102
rect 97274 28046 97342 28102
rect 97398 28046 114970 28102
rect 115026 28046 115094 28102
rect 115150 28046 115218 28102
rect 115274 28046 115342 28102
rect 115398 28046 132970 28102
rect 133026 28046 133094 28102
rect 133150 28046 133218 28102
rect 133274 28046 133342 28102
rect 133398 28046 150970 28102
rect 151026 28046 151094 28102
rect 151150 28046 151218 28102
rect 151274 28046 151342 28102
rect 151398 28046 168970 28102
rect 169026 28046 169094 28102
rect 169150 28046 169218 28102
rect 169274 28046 169342 28102
rect 169398 28046 186970 28102
rect 187026 28046 187094 28102
rect 187150 28046 187218 28102
rect 187274 28046 187342 28102
rect 187398 28046 204970 28102
rect 205026 28046 205094 28102
rect 205150 28046 205218 28102
rect 205274 28046 205342 28102
rect 205398 28046 384970 28102
rect 385026 28046 385094 28102
rect 385150 28046 385218 28102
rect 385274 28046 385342 28102
rect 385398 28046 402970 28102
rect 403026 28046 403094 28102
rect 403150 28046 403218 28102
rect 403274 28046 403342 28102
rect 403398 28046 420970 28102
rect 421026 28046 421094 28102
rect 421150 28046 421218 28102
rect 421274 28046 421342 28102
rect 421398 28046 438970 28102
rect 439026 28046 439094 28102
rect 439150 28046 439218 28102
rect 439274 28046 439342 28102
rect 439398 28046 456970 28102
rect 457026 28046 457094 28102
rect 457150 28046 457218 28102
rect 457274 28046 457342 28102
rect 457398 28046 474970 28102
rect 475026 28046 475094 28102
rect 475150 28046 475218 28102
rect 475274 28046 475342 28102
rect 475398 28046 492970 28102
rect 493026 28046 493094 28102
rect 493150 28046 493218 28102
rect 493274 28046 493342 28102
rect 493398 28046 510970 28102
rect 511026 28046 511094 28102
rect 511150 28046 511218 28102
rect 511274 28046 511342 28102
rect 511398 28046 528970 28102
rect 529026 28046 529094 28102
rect 529150 28046 529218 28102
rect 529274 28046 529342 28102
rect 529398 28046 546970 28102
rect 547026 28046 547094 28102
rect 547150 28046 547218 28102
rect 547274 28046 547342 28102
rect 547398 28046 564970 28102
rect 565026 28046 565094 28102
rect 565150 28046 565218 28102
rect 565274 28046 565342 28102
rect 565398 28046 582970 28102
rect 583026 28046 583094 28102
rect 583150 28046 583218 28102
rect 583274 28046 583342 28102
rect 583398 28046 597456 28102
rect 597512 28046 597580 28102
rect 597636 28046 597704 28102
rect 597760 28046 597828 28102
rect 597884 28046 597980 28102
rect -1916 27978 597980 28046
rect -1916 27922 -1820 27978
rect -1764 27922 -1696 27978
rect -1640 27922 -1572 27978
rect -1516 27922 -1448 27978
rect -1392 27922 6970 27978
rect 7026 27922 7094 27978
rect 7150 27922 7218 27978
rect 7274 27922 7342 27978
rect 7398 27922 24970 27978
rect 25026 27922 25094 27978
rect 25150 27922 25218 27978
rect 25274 27922 25342 27978
rect 25398 27922 42970 27978
rect 43026 27922 43094 27978
rect 43150 27922 43218 27978
rect 43274 27922 43342 27978
rect 43398 27922 60970 27978
rect 61026 27922 61094 27978
rect 61150 27922 61218 27978
rect 61274 27922 61342 27978
rect 61398 27922 78970 27978
rect 79026 27922 79094 27978
rect 79150 27922 79218 27978
rect 79274 27922 79342 27978
rect 79398 27922 96970 27978
rect 97026 27922 97094 27978
rect 97150 27922 97218 27978
rect 97274 27922 97342 27978
rect 97398 27922 114970 27978
rect 115026 27922 115094 27978
rect 115150 27922 115218 27978
rect 115274 27922 115342 27978
rect 115398 27922 132970 27978
rect 133026 27922 133094 27978
rect 133150 27922 133218 27978
rect 133274 27922 133342 27978
rect 133398 27922 150970 27978
rect 151026 27922 151094 27978
rect 151150 27922 151218 27978
rect 151274 27922 151342 27978
rect 151398 27922 168970 27978
rect 169026 27922 169094 27978
rect 169150 27922 169218 27978
rect 169274 27922 169342 27978
rect 169398 27922 186970 27978
rect 187026 27922 187094 27978
rect 187150 27922 187218 27978
rect 187274 27922 187342 27978
rect 187398 27922 204970 27978
rect 205026 27922 205094 27978
rect 205150 27922 205218 27978
rect 205274 27922 205342 27978
rect 205398 27922 384970 27978
rect 385026 27922 385094 27978
rect 385150 27922 385218 27978
rect 385274 27922 385342 27978
rect 385398 27922 402970 27978
rect 403026 27922 403094 27978
rect 403150 27922 403218 27978
rect 403274 27922 403342 27978
rect 403398 27922 420970 27978
rect 421026 27922 421094 27978
rect 421150 27922 421218 27978
rect 421274 27922 421342 27978
rect 421398 27922 438970 27978
rect 439026 27922 439094 27978
rect 439150 27922 439218 27978
rect 439274 27922 439342 27978
rect 439398 27922 456970 27978
rect 457026 27922 457094 27978
rect 457150 27922 457218 27978
rect 457274 27922 457342 27978
rect 457398 27922 474970 27978
rect 475026 27922 475094 27978
rect 475150 27922 475218 27978
rect 475274 27922 475342 27978
rect 475398 27922 492970 27978
rect 493026 27922 493094 27978
rect 493150 27922 493218 27978
rect 493274 27922 493342 27978
rect 493398 27922 510970 27978
rect 511026 27922 511094 27978
rect 511150 27922 511218 27978
rect 511274 27922 511342 27978
rect 511398 27922 528970 27978
rect 529026 27922 529094 27978
rect 529150 27922 529218 27978
rect 529274 27922 529342 27978
rect 529398 27922 546970 27978
rect 547026 27922 547094 27978
rect 547150 27922 547218 27978
rect 547274 27922 547342 27978
rect 547398 27922 564970 27978
rect 565026 27922 565094 27978
rect 565150 27922 565218 27978
rect 565274 27922 565342 27978
rect 565398 27922 582970 27978
rect 583026 27922 583094 27978
rect 583150 27922 583218 27978
rect 583274 27922 583342 27978
rect 583398 27922 597456 27978
rect 597512 27922 597580 27978
rect 597636 27922 597704 27978
rect 597760 27922 597828 27978
rect 597884 27922 597980 27978
rect -1916 27826 597980 27922
rect -1916 22350 597980 22446
rect -1916 22294 -860 22350
rect -804 22294 -736 22350
rect -680 22294 -612 22350
rect -556 22294 -488 22350
rect -432 22294 3250 22350
rect 3306 22294 3374 22350
rect 3430 22294 3498 22350
rect 3554 22294 3622 22350
rect 3678 22294 21250 22350
rect 21306 22294 21374 22350
rect 21430 22294 21498 22350
rect 21554 22294 21622 22350
rect 21678 22294 39250 22350
rect 39306 22294 39374 22350
rect 39430 22294 39498 22350
rect 39554 22294 39622 22350
rect 39678 22294 57250 22350
rect 57306 22294 57374 22350
rect 57430 22294 57498 22350
rect 57554 22294 57622 22350
rect 57678 22294 75250 22350
rect 75306 22294 75374 22350
rect 75430 22294 75498 22350
rect 75554 22294 75622 22350
rect 75678 22294 93250 22350
rect 93306 22294 93374 22350
rect 93430 22294 93498 22350
rect 93554 22294 93622 22350
rect 93678 22294 111250 22350
rect 111306 22294 111374 22350
rect 111430 22294 111498 22350
rect 111554 22294 111622 22350
rect 111678 22294 129250 22350
rect 129306 22294 129374 22350
rect 129430 22294 129498 22350
rect 129554 22294 129622 22350
rect 129678 22294 147250 22350
rect 147306 22294 147374 22350
rect 147430 22294 147498 22350
rect 147554 22294 147622 22350
rect 147678 22294 165250 22350
rect 165306 22294 165374 22350
rect 165430 22294 165498 22350
rect 165554 22294 165622 22350
rect 165678 22294 183250 22350
rect 183306 22294 183374 22350
rect 183430 22294 183498 22350
rect 183554 22294 183622 22350
rect 183678 22294 201250 22350
rect 201306 22294 201374 22350
rect 201430 22294 201498 22350
rect 201554 22294 201622 22350
rect 201678 22294 381250 22350
rect 381306 22294 381374 22350
rect 381430 22294 381498 22350
rect 381554 22294 381622 22350
rect 381678 22294 399250 22350
rect 399306 22294 399374 22350
rect 399430 22294 399498 22350
rect 399554 22294 399622 22350
rect 399678 22294 417250 22350
rect 417306 22294 417374 22350
rect 417430 22294 417498 22350
rect 417554 22294 417622 22350
rect 417678 22294 435250 22350
rect 435306 22294 435374 22350
rect 435430 22294 435498 22350
rect 435554 22294 435622 22350
rect 435678 22294 453250 22350
rect 453306 22294 453374 22350
rect 453430 22294 453498 22350
rect 453554 22294 453622 22350
rect 453678 22294 471250 22350
rect 471306 22294 471374 22350
rect 471430 22294 471498 22350
rect 471554 22294 471622 22350
rect 471678 22294 489250 22350
rect 489306 22294 489374 22350
rect 489430 22294 489498 22350
rect 489554 22294 489622 22350
rect 489678 22294 507250 22350
rect 507306 22294 507374 22350
rect 507430 22294 507498 22350
rect 507554 22294 507622 22350
rect 507678 22294 525250 22350
rect 525306 22294 525374 22350
rect 525430 22294 525498 22350
rect 525554 22294 525622 22350
rect 525678 22294 543250 22350
rect 543306 22294 543374 22350
rect 543430 22294 543498 22350
rect 543554 22294 543622 22350
rect 543678 22294 561250 22350
rect 561306 22294 561374 22350
rect 561430 22294 561498 22350
rect 561554 22294 561622 22350
rect 561678 22294 579250 22350
rect 579306 22294 579374 22350
rect 579430 22294 579498 22350
rect 579554 22294 579622 22350
rect 579678 22294 596496 22350
rect 596552 22294 596620 22350
rect 596676 22294 596744 22350
rect 596800 22294 596868 22350
rect 596924 22294 597980 22350
rect -1916 22226 597980 22294
rect -1916 22170 -860 22226
rect -804 22170 -736 22226
rect -680 22170 -612 22226
rect -556 22170 -488 22226
rect -432 22170 3250 22226
rect 3306 22170 3374 22226
rect 3430 22170 3498 22226
rect 3554 22170 3622 22226
rect 3678 22170 21250 22226
rect 21306 22170 21374 22226
rect 21430 22170 21498 22226
rect 21554 22170 21622 22226
rect 21678 22170 39250 22226
rect 39306 22170 39374 22226
rect 39430 22170 39498 22226
rect 39554 22170 39622 22226
rect 39678 22170 57250 22226
rect 57306 22170 57374 22226
rect 57430 22170 57498 22226
rect 57554 22170 57622 22226
rect 57678 22170 75250 22226
rect 75306 22170 75374 22226
rect 75430 22170 75498 22226
rect 75554 22170 75622 22226
rect 75678 22170 93250 22226
rect 93306 22170 93374 22226
rect 93430 22170 93498 22226
rect 93554 22170 93622 22226
rect 93678 22170 111250 22226
rect 111306 22170 111374 22226
rect 111430 22170 111498 22226
rect 111554 22170 111622 22226
rect 111678 22170 129250 22226
rect 129306 22170 129374 22226
rect 129430 22170 129498 22226
rect 129554 22170 129622 22226
rect 129678 22170 147250 22226
rect 147306 22170 147374 22226
rect 147430 22170 147498 22226
rect 147554 22170 147622 22226
rect 147678 22170 165250 22226
rect 165306 22170 165374 22226
rect 165430 22170 165498 22226
rect 165554 22170 165622 22226
rect 165678 22170 183250 22226
rect 183306 22170 183374 22226
rect 183430 22170 183498 22226
rect 183554 22170 183622 22226
rect 183678 22170 201250 22226
rect 201306 22170 201374 22226
rect 201430 22170 201498 22226
rect 201554 22170 201622 22226
rect 201678 22170 381250 22226
rect 381306 22170 381374 22226
rect 381430 22170 381498 22226
rect 381554 22170 381622 22226
rect 381678 22170 399250 22226
rect 399306 22170 399374 22226
rect 399430 22170 399498 22226
rect 399554 22170 399622 22226
rect 399678 22170 417250 22226
rect 417306 22170 417374 22226
rect 417430 22170 417498 22226
rect 417554 22170 417622 22226
rect 417678 22170 435250 22226
rect 435306 22170 435374 22226
rect 435430 22170 435498 22226
rect 435554 22170 435622 22226
rect 435678 22170 453250 22226
rect 453306 22170 453374 22226
rect 453430 22170 453498 22226
rect 453554 22170 453622 22226
rect 453678 22170 471250 22226
rect 471306 22170 471374 22226
rect 471430 22170 471498 22226
rect 471554 22170 471622 22226
rect 471678 22170 489250 22226
rect 489306 22170 489374 22226
rect 489430 22170 489498 22226
rect 489554 22170 489622 22226
rect 489678 22170 507250 22226
rect 507306 22170 507374 22226
rect 507430 22170 507498 22226
rect 507554 22170 507622 22226
rect 507678 22170 525250 22226
rect 525306 22170 525374 22226
rect 525430 22170 525498 22226
rect 525554 22170 525622 22226
rect 525678 22170 543250 22226
rect 543306 22170 543374 22226
rect 543430 22170 543498 22226
rect 543554 22170 543622 22226
rect 543678 22170 561250 22226
rect 561306 22170 561374 22226
rect 561430 22170 561498 22226
rect 561554 22170 561622 22226
rect 561678 22170 579250 22226
rect 579306 22170 579374 22226
rect 579430 22170 579498 22226
rect 579554 22170 579622 22226
rect 579678 22170 596496 22226
rect 596552 22170 596620 22226
rect 596676 22170 596744 22226
rect 596800 22170 596868 22226
rect 596924 22170 597980 22226
rect -1916 22102 597980 22170
rect -1916 22046 -860 22102
rect -804 22046 -736 22102
rect -680 22046 -612 22102
rect -556 22046 -488 22102
rect -432 22046 3250 22102
rect 3306 22046 3374 22102
rect 3430 22046 3498 22102
rect 3554 22046 3622 22102
rect 3678 22046 21250 22102
rect 21306 22046 21374 22102
rect 21430 22046 21498 22102
rect 21554 22046 21622 22102
rect 21678 22046 39250 22102
rect 39306 22046 39374 22102
rect 39430 22046 39498 22102
rect 39554 22046 39622 22102
rect 39678 22046 57250 22102
rect 57306 22046 57374 22102
rect 57430 22046 57498 22102
rect 57554 22046 57622 22102
rect 57678 22046 75250 22102
rect 75306 22046 75374 22102
rect 75430 22046 75498 22102
rect 75554 22046 75622 22102
rect 75678 22046 93250 22102
rect 93306 22046 93374 22102
rect 93430 22046 93498 22102
rect 93554 22046 93622 22102
rect 93678 22046 111250 22102
rect 111306 22046 111374 22102
rect 111430 22046 111498 22102
rect 111554 22046 111622 22102
rect 111678 22046 129250 22102
rect 129306 22046 129374 22102
rect 129430 22046 129498 22102
rect 129554 22046 129622 22102
rect 129678 22046 147250 22102
rect 147306 22046 147374 22102
rect 147430 22046 147498 22102
rect 147554 22046 147622 22102
rect 147678 22046 165250 22102
rect 165306 22046 165374 22102
rect 165430 22046 165498 22102
rect 165554 22046 165622 22102
rect 165678 22046 183250 22102
rect 183306 22046 183374 22102
rect 183430 22046 183498 22102
rect 183554 22046 183622 22102
rect 183678 22046 201250 22102
rect 201306 22046 201374 22102
rect 201430 22046 201498 22102
rect 201554 22046 201622 22102
rect 201678 22046 381250 22102
rect 381306 22046 381374 22102
rect 381430 22046 381498 22102
rect 381554 22046 381622 22102
rect 381678 22046 399250 22102
rect 399306 22046 399374 22102
rect 399430 22046 399498 22102
rect 399554 22046 399622 22102
rect 399678 22046 417250 22102
rect 417306 22046 417374 22102
rect 417430 22046 417498 22102
rect 417554 22046 417622 22102
rect 417678 22046 435250 22102
rect 435306 22046 435374 22102
rect 435430 22046 435498 22102
rect 435554 22046 435622 22102
rect 435678 22046 453250 22102
rect 453306 22046 453374 22102
rect 453430 22046 453498 22102
rect 453554 22046 453622 22102
rect 453678 22046 471250 22102
rect 471306 22046 471374 22102
rect 471430 22046 471498 22102
rect 471554 22046 471622 22102
rect 471678 22046 489250 22102
rect 489306 22046 489374 22102
rect 489430 22046 489498 22102
rect 489554 22046 489622 22102
rect 489678 22046 507250 22102
rect 507306 22046 507374 22102
rect 507430 22046 507498 22102
rect 507554 22046 507622 22102
rect 507678 22046 525250 22102
rect 525306 22046 525374 22102
rect 525430 22046 525498 22102
rect 525554 22046 525622 22102
rect 525678 22046 543250 22102
rect 543306 22046 543374 22102
rect 543430 22046 543498 22102
rect 543554 22046 543622 22102
rect 543678 22046 561250 22102
rect 561306 22046 561374 22102
rect 561430 22046 561498 22102
rect 561554 22046 561622 22102
rect 561678 22046 579250 22102
rect 579306 22046 579374 22102
rect 579430 22046 579498 22102
rect 579554 22046 579622 22102
rect 579678 22046 596496 22102
rect 596552 22046 596620 22102
rect 596676 22046 596744 22102
rect 596800 22046 596868 22102
rect 596924 22046 597980 22102
rect -1916 21978 597980 22046
rect -1916 21922 -860 21978
rect -804 21922 -736 21978
rect -680 21922 -612 21978
rect -556 21922 -488 21978
rect -432 21922 3250 21978
rect 3306 21922 3374 21978
rect 3430 21922 3498 21978
rect 3554 21922 3622 21978
rect 3678 21922 21250 21978
rect 21306 21922 21374 21978
rect 21430 21922 21498 21978
rect 21554 21922 21622 21978
rect 21678 21922 39250 21978
rect 39306 21922 39374 21978
rect 39430 21922 39498 21978
rect 39554 21922 39622 21978
rect 39678 21922 57250 21978
rect 57306 21922 57374 21978
rect 57430 21922 57498 21978
rect 57554 21922 57622 21978
rect 57678 21922 75250 21978
rect 75306 21922 75374 21978
rect 75430 21922 75498 21978
rect 75554 21922 75622 21978
rect 75678 21922 93250 21978
rect 93306 21922 93374 21978
rect 93430 21922 93498 21978
rect 93554 21922 93622 21978
rect 93678 21922 111250 21978
rect 111306 21922 111374 21978
rect 111430 21922 111498 21978
rect 111554 21922 111622 21978
rect 111678 21922 129250 21978
rect 129306 21922 129374 21978
rect 129430 21922 129498 21978
rect 129554 21922 129622 21978
rect 129678 21922 147250 21978
rect 147306 21922 147374 21978
rect 147430 21922 147498 21978
rect 147554 21922 147622 21978
rect 147678 21922 165250 21978
rect 165306 21922 165374 21978
rect 165430 21922 165498 21978
rect 165554 21922 165622 21978
rect 165678 21922 183250 21978
rect 183306 21922 183374 21978
rect 183430 21922 183498 21978
rect 183554 21922 183622 21978
rect 183678 21922 201250 21978
rect 201306 21922 201374 21978
rect 201430 21922 201498 21978
rect 201554 21922 201622 21978
rect 201678 21922 381250 21978
rect 381306 21922 381374 21978
rect 381430 21922 381498 21978
rect 381554 21922 381622 21978
rect 381678 21922 399250 21978
rect 399306 21922 399374 21978
rect 399430 21922 399498 21978
rect 399554 21922 399622 21978
rect 399678 21922 417250 21978
rect 417306 21922 417374 21978
rect 417430 21922 417498 21978
rect 417554 21922 417622 21978
rect 417678 21922 435250 21978
rect 435306 21922 435374 21978
rect 435430 21922 435498 21978
rect 435554 21922 435622 21978
rect 435678 21922 453250 21978
rect 453306 21922 453374 21978
rect 453430 21922 453498 21978
rect 453554 21922 453622 21978
rect 453678 21922 471250 21978
rect 471306 21922 471374 21978
rect 471430 21922 471498 21978
rect 471554 21922 471622 21978
rect 471678 21922 489250 21978
rect 489306 21922 489374 21978
rect 489430 21922 489498 21978
rect 489554 21922 489622 21978
rect 489678 21922 507250 21978
rect 507306 21922 507374 21978
rect 507430 21922 507498 21978
rect 507554 21922 507622 21978
rect 507678 21922 525250 21978
rect 525306 21922 525374 21978
rect 525430 21922 525498 21978
rect 525554 21922 525622 21978
rect 525678 21922 543250 21978
rect 543306 21922 543374 21978
rect 543430 21922 543498 21978
rect 543554 21922 543622 21978
rect 543678 21922 561250 21978
rect 561306 21922 561374 21978
rect 561430 21922 561498 21978
rect 561554 21922 561622 21978
rect 561678 21922 579250 21978
rect 579306 21922 579374 21978
rect 579430 21922 579498 21978
rect 579554 21922 579622 21978
rect 579678 21922 596496 21978
rect 596552 21922 596620 21978
rect 596676 21922 596744 21978
rect 596800 21922 596868 21978
rect 596924 21922 597980 21978
rect -1916 21826 597980 21922
rect -1916 10350 597980 10446
rect -1916 10294 -1820 10350
rect -1764 10294 -1696 10350
rect -1640 10294 -1572 10350
rect -1516 10294 -1448 10350
rect -1392 10294 6970 10350
rect 7026 10294 7094 10350
rect 7150 10294 7218 10350
rect 7274 10294 7342 10350
rect 7398 10294 24970 10350
rect 25026 10294 25094 10350
rect 25150 10294 25218 10350
rect 25274 10294 25342 10350
rect 25398 10294 42970 10350
rect 43026 10294 43094 10350
rect 43150 10294 43218 10350
rect 43274 10294 43342 10350
rect 43398 10294 60970 10350
rect 61026 10294 61094 10350
rect 61150 10294 61218 10350
rect 61274 10294 61342 10350
rect 61398 10294 78970 10350
rect 79026 10294 79094 10350
rect 79150 10294 79218 10350
rect 79274 10294 79342 10350
rect 79398 10294 96970 10350
rect 97026 10294 97094 10350
rect 97150 10294 97218 10350
rect 97274 10294 97342 10350
rect 97398 10294 114970 10350
rect 115026 10294 115094 10350
rect 115150 10294 115218 10350
rect 115274 10294 115342 10350
rect 115398 10294 132970 10350
rect 133026 10294 133094 10350
rect 133150 10294 133218 10350
rect 133274 10294 133342 10350
rect 133398 10294 150970 10350
rect 151026 10294 151094 10350
rect 151150 10294 151218 10350
rect 151274 10294 151342 10350
rect 151398 10294 168970 10350
rect 169026 10294 169094 10350
rect 169150 10294 169218 10350
rect 169274 10294 169342 10350
rect 169398 10294 186970 10350
rect 187026 10294 187094 10350
rect 187150 10294 187218 10350
rect 187274 10294 187342 10350
rect 187398 10294 204970 10350
rect 205026 10294 205094 10350
rect 205150 10294 205218 10350
rect 205274 10294 205342 10350
rect 205398 10294 384970 10350
rect 385026 10294 385094 10350
rect 385150 10294 385218 10350
rect 385274 10294 385342 10350
rect 385398 10294 402970 10350
rect 403026 10294 403094 10350
rect 403150 10294 403218 10350
rect 403274 10294 403342 10350
rect 403398 10294 420970 10350
rect 421026 10294 421094 10350
rect 421150 10294 421218 10350
rect 421274 10294 421342 10350
rect 421398 10294 438970 10350
rect 439026 10294 439094 10350
rect 439150 10294 439218 10350
rect 439274 10294 439342 10350
rect 439398 10294 456970 10350
rect 457026 10294 457094 10350
rect 457150 10294 457218 10350
rect 457274 10294 457342 10350
rect 457398 10294 474970 10350
rect 475026 10294 475094 10350
rect 475150 10294 475218 10350
rect 475274 10294 475342 10350
rect 475398 10294 492970 10350
rect 493026 10294 493094 10350
rect 493150 10294 493218 10350
rect 493274 10294 493342 10350
rect 493398 10294 510970 10350
rect 511026 10294 511094 10350
rect 511150 10294 511218 10350
rect 511274 10294 511342 10350
rect 511398 10294 528970 10350
rect 529026 10294 529094 10350
rect 529150 10294 529218 10350
rect 529274 10294 529342 10350
rect 529398 10294 546970 10350
rect 547026 10294 547094 10350
rect 547150 10294 547218 10350
rect 547274 10294 547342 10350
rect 547398 10294 564970 10350
rect 565026 10294 565094 10350
rect 565150 10294 565218 10350
rect 565274 10294 565342 10350
rect 565398 10294 582970 10350
rect 583026 10294 583094 10350
rect 583150 10294 583218 10350
rect 583274 10294 583342 10350
rect 583398 10294 597456 10350
rect 597512 10294 597580 10350
rect 597636 10294 597704 10350
rect 597760 10294 597828 10350
rect 597884 10294 597980 10350
rect -1916 10226 597980 10294
rect -1916 10170 -1820 10226
rect -1764 10170 -1696 10226
rect -1640 10170 -1572 10226
rect -1516 10170 -1448 10226
rect -1392 10170 6970 10226
rect 7026 10170 7094 10226
rect 7150 10170 7218 10226
rect 7274 10170 7342 10226
rect 7398 10170 24970 10226
rect 25026 10170 25094 10226
rect 25150 10170 25218 10226
rect 25274 10170 25342 10226
rect 25398 10170 42970 10226
rect 43026 10170 43094 10226
rect 43150 10170 43218 10226
rect 43274 10170 43342 10226
rect 43398 10170 60970 10226
rect 61026 10170 61094 10226
rect 61150 10170 61218 10226
rect 61274 10170 61342 10226
rect 61398 10170 78970 10226
rect 79026 10170 79094 10226
rect 79150 10170 79218 10226
rect 79274 10170 79342 10226
rect 79398 10170 96970 10226
rect 97026 10170 97094 10226
rect 97150 10170 97218 10226
rect 97274 10170 97342 10226
rect 97398 10170 114970 10226
rect 115026 10170 115094 10226
rect 115150 10170 115218 10226
rect 115274 10170 115342 10226
rect 115398 10170 132970 10226
rect 133026 10170 133094 10226
rect 133150 10170 133218 10226
rect 133274 10170 133342 10226
rect 133398 10170 150970 10226
rect 151026 10170 151094 10226
rect 151150 10170 151218 10226
rect 151274 10170 151342 10226
rect 151398 10170 168970 10226
rect 169026 10170 169094 10226
rect 169150 10170 169218 10226
rect 169274 10170 169342 10226
rect 169398 10170 186970 10226
rect 187026 10170 187094 10226
rect 187150 10170 187218 10226
rect 187274 10170 187342 10226
rect 187398 10170 204970 10226
rect 205026 10170 205094 10226
rect 205150 10170 205218 10226
rect 205274 10170 205342 10226
rect 205398 10170 384970 10226
rect 385026 10170 385094 10226
rect 385150 10170 385218 10226
rect 385274 10170 385342 10226
rect 385398 10170 402970 10226
rect 403026 10170 403094 10226
rect 403150 10170 403218 10226
rect 403274 10170 403342 10226
rect 403398 10170 420970 10226
rect 421026 10170 421094 10226
rect 421150 10170 421218 10226
rect 421274 10170 421342 10226
rect 421398 10170 438970 10226
rect 439026 10170 439094 10226
rect 439150 10170 439218 10226
rect 439274 10170 439342 10226
rect 439398 10170 456970 10226
rect 457026 10170 457094 10226
rect 457150 10170 457218 10226
rect 457274 10170 457342 10226
rect 457398 10170 474970 10226
rect 475026 10170 475094 10226
rect 475150 10170 475218 10226
rect 475274 10170 475342 10226
rect 475398 10170 492970 10226
rect 493026 10170 493094 10226
rect 493150 10170 493218 10226
rect 493274 10170 493342 10226
rect 493398 10170 510970 10226
rect 511026 10170 511094 10226
rect 511150 10170 511218 10226
rect 511274 10170 511342 10226
rect 511398 10170 528970 10226
rect 529026 10170 529094 10226
rect 529150 10170 529218 10226
rect 529274 10170 529342 10226
rect 529398 10170 546970 10226
rect 547026 10170 547094 10226
rect 547150 10170 547218 10226
rect 547274 10170 547342 10226
rect 547398 10170 564970 10226
rect 565026 10170 565094 10226
rect 565150 10170 565218 10226
rect 565274 10170 565342 10226
rect 565398 10170 582970 10226
rect 583026 10170 583094 10226
rect 583150 10170 583218 10226
rect 583274 10170 583342 10226
rect 583398 10170 597456 10226
rect 597512 10170 597580 10226
rect 597636 10170 597704 10226
rect 597760 10170 597828 10226
rect 597884 10170 597980 10226
rect -1916 10102 597980 10170
rect -1916 10046 -1820 10102
rect -1764 10046 -1696 10102
rect -1640 10046 -1572 10102
rect -1516 10046 -1448 10102
rect -1392 10046 6970 10102
rect 7026 10046 7094 10102
rect 7150 10046 7218 10102
rect 7274 10046 7342 10102
rect 7398 10046 24970 10102
rect 25026 10046 25094 10102
rect 25150 10046 25218 10102
rect 25274 10046 25342 10102
rect 25398 10046 42970 10102
rect 43026 10046 43094 10102
rect 43150 10046 43218 10102
rect 43274 10046 43342 10102
rect 43398 10046 60970 10102
rect 61026 10046 61094 10102
rect 61150 10046 61218 10102
rect 61274 10046 61342 10102
rect 61398 10046 78970 10102
rect 79026 10046 79094 10102
rect 79150 10046 79218 10102
rect 79274 10046 79342 10102
rect 79398 10046 96970 10102
rect 97026 10046 97094 10102
rect 97150 10046 97218 10102
rect 97274 10046 97342 10102
rect 97398 10046 114970 10102
rect 115026 10046 115094 10102
rect 115150 10046 115218 10102
rect 115274 10046 115342 10102
rect 115398 10046 132970 10102
rect 133026 10046 133094 10102
rect 133150 10046 133218 10102
rect 133274 10046 133342 10102
rect 133398 10046 150970 10102
rect 151026 10046 151094 10102
rect 151150 10046 151218 10102
rect 151274 10046 151342 10102
rect 151398 10046 168970 10102
rect 169026 10046 169094 10102
rect 169150 10046 169218 10102
rect 169274 10046 169342 10102
rect 169398 10046 186970 10102
rect 187026 10046 187094 10102
rect 187150 10046 187218 10102
rect 187274 10046 187342 10102
rect 187398 10046 204970 10102
rect 205026 10046 205094 10102
rect 205150 10046 205218 10102
rect 205274 10046 205342 10102
rect 205398 10046 384970 10102
rect 385026 10046 385094 10102
rect 385150 10046 385218 10102
rect 385274 10046 385342 10102
rect 385398 10046 402970 10102
rect 403026 10046 403094 10102
rect 403150 10046 403218 10102
rect 403274 10046 403342 10102
rect 403398 10046 420970 10102
rect 421026 10046 421094 10102
rect 421150 10046 421218 10102
rect 421274 10046 421342 10102
rect 421398 10046 438970 10102
rect 439026 10046 439094 10102
rect 439150 10046 439218 10102
rect 439274 10046 439342 10102
rect 439398 10046 456970 10102
rect 457026 10046 457094 10102
rect 457150 10046 457218 10102
rect 457274 10046 457342 10102
rect 457398 10046 474970 10102
rect 475026 10046 475094 10102
rect 475150 10046 475218 10102
rect 475274 10046 475342 10102
rect 475398 10046 492970 10102
rect 493026 10046 493094 10102
rect 493150 10046 493218 10102
rect 493274 10046 493342 10102
rect 493398 10046 510970 10102
rect 511026 10046 511094 10102
rect 511150 10046 511218 10102
rect 511274 10046 511342 10102
rect 511398 10046 528970 10102
rect 529026 10046 529094 10102
rect 529150 10046 529218 10102
rect 529274 10046 529342 10102
rect 529398 10046 546970 10102
rect 547026 10046 547094 10102
rect 547150 10046 547218 10102
rect 547274 10046 547342 10102
rect 547398 10046 564970 10102
rect 565026 10046 565094 10102
rect 565150 10046 565218 10102
rect 565274 10046 565342 10102
rect 565398 10046 582970 10102
rect 583026 10046 583094 10102
rect 583150 10046 583218 10102
rect 583274 10046 583342 10102
rect 583398 10046 597456 10102
rect 597512 10046 597580 10102
rect 597636 10046 597704 10102
rect 597760 10046 597828 10102
rect 597884 10046 597980 10102
rect -1916 9978 597980 10046
rect -1916 9922 -1820 9978
rect -1764 9922 -1696 9978
rect -1640 9922 -1572 9978
rect -1516 9922 -1448 9978
rect -1392 9922 6970 9978
rect 7026 9922 7094 9978
rect 7150 9922 7218 9978
rect 7274 9922 7342 9978
rect 7398 9922 24970 9978
rect 25026 9922 25094 9978
rect 25150 9922 25218 9978
rect 25274 9922 25342 9978
rect 25398 9922 42970 9978
rect 43026 9922 43094 9978
rect 43150 9922 43218 9978
rect 43274 9922 43342 9978
rect 43398 9922 60970 9978
rect 61026 9922 61094 9978
rect 61150 9922 61218 9978
rect 61274 9922 61342 9978
rect 61398 9922 78970 9978
rect 79026 9922 79094 9978
rect 79150 9922 79218 9978
rect 79274 9922 79342 9978
rect 79398 9922 96970 9978
rect 97026 9922 97094 9978
rect 97150 9922 97218 9978
rect 97274 9922 97342 9978
rect 97398 9922 114970 9978
rect 115026 9922 115094 9978
rect 115150 9922 115218 9978
rect 115274 9922 115342 9978
rect 115398 9922 132970 9978
rect 133026 9922 133094 9978
rect 133150 9922 133218 9978
rect 133274 9922 133342 9978
rect 133398 9922 150970 9978
rect 151026 9922 151094 9978
rect 151150 9922 151218 9978
rect 151274 9922 151342 9978
rect 151398 9922 168970 9978
rect 169026 9922 169094 9978
rect 169150 9922 169218 9978
rect 169274 9922 169342 9978
rect 169398 9922 186970 9978
rect 187026 9922 187094 9978
rect 187150 9922 187218 9978
rect 187274 9922 187342 9978
rect 187398 9922 204970 9978
rect 205026 9922 205094 9978
rect 205150 9922 205218 9978
rect 205274 9922 205342 9978
rect 205398 9922 384970 9978
rect 385026 9922 385094 9978
rect 385150 9922 385218 9978
rect 385274 9922 385342 9978
rect 385398 9922 402970 9978
rect 403026 9922 403094 9978
rect 403150 9922 403218 9978
rect 403274 9922 403342 9978
rect 403398 9922 420970 9978
rect 421026 9922 421094 9978
rect 421150 9922 421218 9978
rect 421274 9922 421342 9978
rect 421398 9922 438970 9978
rect 439026 9922 439094 9978
rect 439150 9922 439218 9978
rect 439274 9922 439342 9978
rect 439398 9922 456970 9978
rect 457026 9922 457094 9978
rect 457150 9922 457218 9978
rect 457274 9922 457342 9978
rect 457398 9922 474970 9978
rect 475026 9922 475094 9978
rect 475150 9922 475218 9978
rect 475274 9922 475342 9978
rect 475398 9922 492970 9978
rect 493026 9922 493094 9978
rect 493150 9922 493218 9978
rect 493274 9922 493342 9978
rect 493398 9922 510970 9978
rect 511026 9922 511094 9978
rect 511150 9922 511218 9978
rect 511274 9922 511342 9978
rect 511398 9922 528970 9978
rect 529026 9922 529094 9978
rect 529150 9922 529218 9978
rect 529274 9922 529342 9978
rect 529398 9922 546970 9978
rect 547026 9922 547094 9978
rect 547150 9922 547218 9978
rect 547274 9922 547342 9978
rect 547398 9922 564970 9978
rect 565026 9922 565094 9978
rect 565150 9922 565218 9978
rect 565274 9922 565342 9978
rect 565398 9922 582970 9978
rect 583026 9922 583094 9978
rect 583150 9922 583218 9978
rect 583274 9922 583342 9978
rect 583398 9922 597456 9978
rect 597512 9922 597580 9978
rect 597636 9922 597704 9978
rect 597760 9922 597828 9978
rect 597884 9922 597980 9978
rect -1916 9826 597980 9922
rect -1916 4350 597980 4446
rect -1916 4294 -860 4350
rect -804 4294 -736 4350
rect -680 4294 -612 4350
rect -556 4294 -488 4350
rect -432 4294 3250 4350
rect 3306 4294 3374 4350
rect 3430 4294 3498 4350
rect 3554 4294 3622 4350
rect 3678 4294 21250 4350
rect 21306 4294 21374 4350
rect 21430 4294 21498 4350
rect 21554 4294 21622 4350
rect 21678 4294 39250 4350
rect 39306 4294 39374 4350
rect 39430 4294 39498 4350
rect 39554 4294 39622 4350
rect 39678 4294 57250 4350
rect 57306 4294 57374 4350
rect 57430 4294 57498 4350
rect 57554 4294 57622 4350
rect 57678 4294 75250 4350
rect 75306 4294 75374 4350
rect 75430 4294 75498 4350
rect 75554 4294 75622 4350
rect 75678 4294 93250 4350
rect 93306 4294 93374 4350
rect 93430 4294 93498 4350
rect 93554 4294 93622 4350
rect 93678 4294 111250 4350
rect 111306 4294 111374 4350
rect 111430 4294 111498 4350
rect 111554 4294 111622 4350
rect 111678 4294 129250 4350
rect 129306 4294 129374 4350
rect 129430 4294 129498 4350
rect 129554 4294 129622 4350
rect 129678 4294 147250 4350
rect 147306 4294 147374 4350
rect 147430 4294 147498 4350
rect 147554 4294 147622 4350
rect 147678 4294 165250 4350
rect 165306 4294 165374 4350
rect 165430 4294 165498 4350
rect 165554 4294 165622 4350
rect 165678 4294 183250 4350
rect 183306 4294 183374 4350
rect 183430 4294 183498 4350
rect 183554 4294 183622 4350
rect 183678 4294 201250 4350
rect 201306 4294 201374 4350
rect 201430 4294 201498 4350
rect 201554 4294 201622 4350
rect 201678 4294 219250 4350
rect 219306 4294 219374 4350
rect 219430 4294 219498 4350
rect 219554 4294 219622 4350
rect 219678 4294 237250 4350
rect 237306 4294 237374 4350
rect 237430 4294 237498 4350
rect 237554 4294 237622 4350
rect 237678 4294 255250 4350
rect 255306 4294 255374 4350
rect 255430 4294 255498 4350
rect 255554 4294 255622 4350
rect 255678 4294 273250 4350
rect 273306 4294 273374 4350
rect 273430 4294 273498 4350
rect 273554 4294 273622 4350
rect 273678 4294 291250 4350
rect 291306 4294 291374 4350
rect 291430 4294 291498 4350
rect 291554 4294 291622 4350
rect 291678 4294 309250 4350
rect 309306 4294 309374 4350
rect 309430 4294 309498 4350
rect 309554 4294 309622 4350
rect 309678 4294 327250 4350
rect 327306 4294 327374 4350
rect 327430 4294 327498 4350
rect 327554 4294 327622 4350
rect 327678 4294 345250 4350
rect 345306 4294 345374 4350
rect 345430 4294 345498 4350
rect 345554 4294 345622 4350
rect 345678 4294 363250 4350
rect 363306 4294 363374 4350
rect 363430 4294 363498 4350
rect 363554 4294 363622 4350
rect 363678 4294 381250 4350
rect 381306 4294 381374 4350
rect 381430 4294 381498 4350
rect 381554 4294 381622 4350
rect 381678 4294 399250 4350
rect 399306 4294 399374 4350
rect 399430 4294 399498 4350
rect 399554 4294 399622 4350
rect 399678 4294 417250 4350
rect 417306 4294 417374 4350
rect 417430 4294 417498 4350
rect 417554 4294 417622 4350
rect 417678 4294 435250 4350
rect 435306 4294 435374 4350
rect 435430 4294 435498 4350
rect 435554 4294 435622 4350
rect 435678 4294 453250 4350
rect 453306 4294 453374 4350
rect 453430 4294 453498 4350
rect 453554 4294 453622 4350
rect 453678 4294 471250 4350
rect 471306 4294 471374 4350
rect 471430 4294 471498 4350
rect 471554 4294 471622 4350
rect 471678 4294 489250 4350
rect 489306 4294 489374 4350
rect 489430 4294 489498 4350
rect 489554 4294 489622 4350
rect 489678 4294 507250 4350
rect 507306 4294 507374 4350
rect 507430 4294 507498 4350
rect 507554 4294 507622 4350
rect 507678 4294 525250 4350
rect 525306 4294 525374 4350
rect 525430 4294 525498 4350
rect 525554 4294 525622 4350
rect 525678 4294 543250 4350
rect 543306 4294 543374 4350
rect 543430 4294 543498 4350
rect 543554 4294 543622 4350
rect 543678 4294 561250 4350
rect 561306 4294 561374 4350
rect 561430 4294 561498 4350
rect 561554 4294 561622 4350
rect 561678 4294 579250 4350
rect 579306 4294 579374 4350
rect 579430 4294 579498 4350
rect 579554 4294 579622 4350
rect 579678 4294 596496 4350
rect 596552 4294 596620 4350
rect 596676 4294 596744 4350
rect 596800 4294 596868 4350
rect 596924 4294 597980 4350
rect -1916 4226 597980 4294
rect -1916 4170 -860 4226
rect -804 4170 -736 4226
rect -680 4170 -612 4226
rect -556 4170 -488 4226
rect -432 4170 3250 4226
rect 3306 4170 3374 4226
rect 3430 4170 3498 4226
rect 3554 4170 3622 4226
rect 3678 4170 21250 4226
rect 21306 4170 21374 4226
rect 21430 4170 21498 4226
rect 21554 4170 21622 4226
rect 21678 4170 39250 4226
rect 39306 4170 39374 4226
rect 39430 4170 39498 4226
rect 39554 4170 39622 4226
rect 39678 4170 57250 4226
rect 57306 4170 57374 4226
rect 57430 4170 57498 4226
rect 57554 4170 57622 4226
rect 57678 4170 75250 4226
rect 75306 4170 75374 4226
rect 75430 4170 75498 4226
rect 75554 4170 75622 4226
rect 75678 4170 93250 4226
rect 93306 4170 93374 4226
rect 93430 4170 93498 4226
rect 93554 4170 93622 4226
rect 93678 4170 111250 4226
rect 111306 4170 111374 4226
rect 111430 4170 111498 4226
rect 111554 4170 111622 4226
rect 111678 4170 129250 4226
rect 129306 4170 129374 4226
rect 129430 4170 129498 4226
rect 129554 4170 129622 4226
rect 129678 4170 147250 4226
rect 147306 4170 147374 4226
rect 147430 4170 147498 4226
rect 147554 4170 147622 4226
rect 147678 4170 165250 4226
rect 165306 4170 165374 4226
rect 165430 4170 165498 4226
rect 165554 4170 165622 4226
rect 165678 4170 183250 4226
rect 183306 4170 183374 4226
rect 183430 4170 183498 4226
rect 183554 4170 183622 4226
rect 183678 4170 201250 4226
rect 201306 4170 201374 4226
rect 201430 4170 201498 4226
rect 201554 4170 201622 4226
rect 201678 4170 219250 4226
rect 219306 4170 219374 4226
rect 219430 4170 219498 4226
rect 219554 4170 219622 4226
rect 219678 4170 237250 4226
rect 237306 4170 237374 4226
rect 237430 4170 237498 4226
rect 237554 4170 237622 4226
rect 237678 4170 255250 4226
rect 255306 4170 255374 4226
rect 255430 4170 255498 4226
rect 255554 4170 255622 4226
rect 255678 4170 273250 4226
rect 273306 4170 273374 4226
rect 273430 4170 273498 4226
rect 273554 4170 273622 4226
rect 273678 4170 291250 4226
rect 291306 4170 291374 4226
rect 291430 4170 291498 4226
rect 291554 4170 291622 4226
rect 291678 4170 309250 4226
rect 309306 4170 309374 4226
rect 309430 4170 309498 4226
rect 309554 4170 309622 4226
rect 309678 4170 327250 4226
rect 327306 4170 327374 4226
rect 327430 4170 327498 4226
rect 327554 4170 327622 4226
rect 327678 4170 345250 4226
rect 345306 4170 345374 4226
rect 345430 4170 345498 4226
rect 345554 4170 345622 4226
rect 345678 4170 363250 4226
rect 363306 4170 363374 4226
rect 363430 4170 363498 4226
rect 363554 4170 363622 4226
rect 363678 4170 381250 4226
rect 381306 4170 381374 4226
rect 381430 4170 381498 4226
rect 381554 4170 381622 4226
rect 381678 4170 399250 4226
rect 399306 4170 399374 4226
rect 399430 4170 399498 4226
rect 399554 4170 399622 4226
rect 399678 4170 417250 4226
rect 417306 4170 417374 4226
rect 417430 4170 417498 4226
rect 417554 4170 417622 4226
rect 417678 4170 435250 4226
rect 435306 4170 435374 4226
rect 435430 4170 435498 4226
rect 435554 4170 435622 4226
rect 435678 4170 453250 4226
rect 453306 4170 453374 4226
rect 453430 4170 453498 4226
rect 453554 4170 453622 4226
rect 453678 4170 471250 4226
rect 471306 4170 471374 4226
rect 471430 4170 471498 4226
rect 471554 4170 471622 4226
rect 471678 4170 489250 4226
rect 489306 4170 489374 4226
rect 489430 4170 489498 4226
rect 489554 4170 489622 4226
rect 489678 4170 507250 4226
rect 507306 4170 507374 4226
rect 507430 4170 507498 4226
rect 507554 4170 507622 4226
rect 507678 4170 525250 4226
rect 525306 4170 525374 4226
rect 525430 4170 525498 4226
rect 525554 4170 525622 4226
rect 525678 4170 543250 4226
rect 543306 4170 543374 4226
rect 543430 4170 543498 4226
rect 543554 4170 543622 4226
rect 543678 4170 561250 4226
rect 561306 4170 561374 4226
rect 561430 4170 561498 4226
rect 561554 4170 561622 4226
rect 561678 4170 579250 4226
rect 579306 4170 579374 4226
rect 579430 4170 579498 4226
rect 579554 4170 579622 4226
rect 579678 4170 596496 4226
rect 596552 4170 596620 4226
rect 596676 4170 596744 4226
rect 596800 4170 596868 4226
rect 596924 4170 597980 4226
rect -1916 4102 597980 4170
rect -1916 4046 -860 4102
rect -804 4046 -736 4102
rect -680 4046 -612 4102
rect -556 4046 -488 4102
rect -432 4046 3250 4102
rect 3306 4046 3374 4102
rect 3430 4046 3498 4102
rect 3554 4046 3622 4102
rect 3678 4046 21250 4102
rect 21306 4046 21374 4102
rect 21430 4046 21498 4102
rect 21554 4046 21622 4102
rect 21678 4046 39250 4102
rect 39306 4046 39374 4102
rect 39430 4046 39498 4102
rect 39554 4046 39622 4102
rect 39678 4046 57250 4102
rect 57306 4046 57374 4102
rect 57430 4046 57498 4102
rect 57554 4046 57622 4102
rect 57678 4046 75250 4102
rect 75306 4046 75374 4102
rect 75430 4046 75498 4102
rect 75554 4046 75622 4102
rect 75678 4046 93250 4102
rect 93306 4046 93374 4102
rect 93430 4046 93498 4102
rect 93554 4046 93622 4102
rect 93678 4046 111250 4102
rect 111306 4046 111374 4102
rect 111430 4046 111498 4102
rect 111554 4046 111622 4102
rect 111678 4046 129250 4102
rect 129306 4046 129374 4102
rect 129430 4046 129498 4102
rect 129554 4046 129622 4102
rect 129678 4046 147250 4102
rect 147306 4046 147374 4102
rect 147430 4046 147498 4102
rect 147554 4046 147622 4102
rect 147678 4046 165250 4102
rect 165306 4046 165374 4102
rect 165430 4046 165498 4102
rect 165554 4046 165622 4102
rect 165678 4046 183250 4102
rect 183306 4046 183374 4102
rect 183430 4046 183498 4102
rect 183554 4046 183622 4102
rect 183678 4046 201250 4102
rect 201306 4046 201374 4102
rect 201430 4046 201498 4102
rect 201554 4046 201622 4102
rect 201678 4046 219250 4102
rect 219306 4046 219374 4102
rect 219430 4046 219498 4102
rect 219554 4046 219622 4102
rect 219678 4046 237250 4102
rect 237306 4046 237374 4102
rect 237430 4046 237498 4102
rect 237554 4046 237622 4102
rect 237678 4046 255250 4102
rect 255306 4046 255374 4102
rect 255430 4046 255498 4102
rect 255554 4046 255622 4102
rect 255678 4046 273250 4102
rect 273306 4046 273374 4102
rect 273430 4046 273498 4102
rect 273554 4046 273622 4102
rect 273678 4046 291250 4102
rect 291306 4046 291374 4102
rect 291430 4046 291498 4102
rect 291554 4046 291622 4102
rect 291678 4046 309250 4102
rect 309306 4046 309374 4102
rect 309430 4046 309498 4102
rect 309554 4046 309622 4102
rect 309678 4046 327250 4102
rect 327306 4046 327374 4102
rect 327430 4046 327498 4102
rect 327554 4046 327622 4102
rect 327678 4046 345250 4102
rect 345306 4046 345374 4102
rect 345430 4046 345498 4102
rect 345554 4046 345622 4102
rect 345678 4046 363250 4102
rect 363306 4046 363374 4102
rect 363430 4046 363498 4102
rect 363554 4046 363622 4102
rect 363678 4046 381250 4102
rect 381306 4046 381374 4102
rect 381430 4046 381498 4102
rect 381554 4046 381622 4102
rect 381678 4046 399250 4102
rect 399306 4046 399374 4102
rect 399430 4046 399498 4102
rect 399554 4046 399622 4102
rect 399678 4046 417250 4102
rect 417306 4046 417374 4102
rect 417430 4046 417498 4102
rect 417554 4046 417622 4102
rect 417678 4046 435250 4102
rect 435306 4046 435374 4102
rect 435430 4046 435498 4102
rect 435554 4046 435622 4102
rect 435678 4046 453250 4102
rect 453306 4046 453374 4102
rect 453430 4046 453498 4102
rect 453554 4046 453622 4102
rect 453678 4046 471250 4102
rect 471306 4046 471374 4102
rect 471430 4046 471498 4102
rect 471554 4046 471622 4102
rect 471678 4046 489250 4102
rect 489306 4046 489374 4102
rect 489430 4046 489498 4102
rect 489554 4046 489622 4102
rect 489678 4046 507250 4102
rect 507306 4046 507374 4102
rect 507430 4046 507498 4102
rect 507554 4046 507622 4102
rect 507678 4046 525250 4102
rect 525306 4046 525374 4102
rect 525430 4046 525498 4102
rect 525554 4046 525622 4102
rect 525678 4046 543250 4102
rect 543306 4046 543374 4102
rect 543430 4046 543498 4102
rect 543554 4046 543622 4102
rect 543678 4046 561250 4102
rect 561306 4046 561374 4102
rect 561430 4046 561498 4102
rect 561554 4046 561622 4102
rect 561678 4046 579250 4102
rect 579306 4046 579374 4102
rect 579430 4046 579498 4102
rect 579554 4046 579622 4102
rect 579678 4046 596496 4102
rect 596552 4046 596620 4102
rect 596676 4046 596744 4102
rect 596800 4046 596868 4102
rect 596924 4046 597980 4102
rect -1916 3978 597980 4046
rect -1916 3922 -860 3978
rect -804 3922 -736 3978
rect -680 3922 -612 3978
rect -556 3922 -488 3978
rect -432 3922 3250 3978
rect 3306 3922 3374 3978
rect 3430 3922 3498 3978
rect 3554 3922 3622 3978
rect 3678 3922 21250 3978
rect 21306 3922 21374 3978
rect 21430 3922 21498 3978
rect 21554 3922 21622 3978
rect 21678 3922 39250 3978
rect 39306 3922 39374 3978
rect 39430 3922 39498 3978
rect 39554 3922 39622 3978
rect 39678 3922 57250 3978
rect 57306 3922 57374 3978
rect 57430 3922 57498 3978
rect 57554 3922 57622 3978
rect 57678 3922 75250 3978
rect 75306 3922 75374 3978
rect 75430 3922 75498 3978
rect 75554 3922 75622 3978
rect 75678 3922 93250 3978
rect 93306 3922 93374 3978
rect 93430 3922 93498 3978
rect 93554 3922 93622 3978
rect 93678 3922 111250 3978
rect 111306 3922 111374 3978
rect 111430 3922 111498 3978
rect 111554 3922 111622 3978
rect 111678 3922 129250 3978
rect 129306 3922 129374 3978
rect 129430 3922 129498 3978
rect 129554 3922 129622 3978
rect 129678 3922 147250 3978
rect 147306 3922 147374 3978
rect 147430 3922 147498 3978
rect 147554 3922 147622 3978
rect 147678 3922 165250 3978
rect 165306 3922 165374 3978
rect 165430 3922 165498 3978
rect 165554 3922 165622 3978
rect 165678 3922 183250 3978
rect 183306 3922 183374 3978
rect 183430 3922 183498 3978
rect 183554 3922 183622 3978
rect 183678 3922 201250 3978
rect 201306 3922 201374 3978
rect 201430 3922 201498 3978
rect 201554 3922 201622 3978
rect 201678 3922 219250 3978
rect 219306 3922 219374 3978
rect 219430 3922 219498 3978
rect 219554 3922 219622 3978
rect 219678 3922 237250 3978
rect 237306 3922 237374 3978
rect 237430 3922 237498 3978
rect 237554 3922 237622 3978
rect 237678 3922 255250 3978
rect 255306 3922 255374 3978
rect 255430 3922 255498 3978
rect 255554 3922 255622 3978
rect 255678 3922 273250 3978
rect 273306 3922 273374 3978
rect 273430 3922 273498 3978
rect 273554 3922 273622 3978
rect 273678 3922 291250 3978
rect 291306 3922 291374 3978
rect 291430 3922 291498 3978
rect 291554 3922 291622 3978
rect 291678 3922 309250 3978
rect 309306 3922 309374 3978
rect 309430 3922 309498 3978
rect 309554 3922 309622 3978
rect 309678 3922 327250 3978
rect 327306 3922 327374 3978
rect 327430 3922 327498 3978
rect 327554 3922 327622 3978
rect 327678 3922 345250 3978
rect 345306 3922 345374 3978
rect 345430 3922 345498 3978
rect 345554 3922 345622 3978
rect 345678 3922 363250 3978
rect 363306 3922 363374 3978
rect 363430 3922 363498 3978
rect 363554 3922 363622 3978
rect 363678 3922 381250 3978
rect 381306 3922 381374 3978
rect 381430 3922 381498 3978
rect 381554 3922 381622 3978
rect 381678 3922 399250 3978
rect 399306 3922 399374 3978
rect 399430 3922 399498 3978
rect 399554 3922 399622 3978
rect 399678 3922 417250 3978
rect 417306 3922 417374 3978
rect 417430 3922 417498 3978
rect 417554 3922 417622 3978
rect 417678 3922 435250 3978
rect 435306 3922 435374 3978
rect 435430 3922 435498 3978
rect 435554 3922 435622 3978
rect 435678 3922 453250 3978
rect 453306 3922 453374 3978
rect 453430 3922 453498 3978
rect 453554 3922 453622 3978
rect 453678 3922 471250 3978
rect 471306 3922 471374 3978
rect 471430 3922 471498 3978
rect 471554 3922 471622 3978
rect 471678 3922 489250 3978
rect 489306 3922 489374 3978
rect 489430 3922 489498 3978
rect 489554 3922 489622 3978
rect 489678 3922 507250 3978
rect 507306 3922 507374 3978
rect 507430 3922 507498 3978
rect 507554 3922 507622 3978
rect 507678 3922 525250 3978
rect 525306 3922 525374 3978
rect 525430 3922 525498 3978
rect 525554 3922 525622 3978
rect 525678 3922 543250 3978
rect 543306 3922 543374 3978
rect 543430 3922 543498 3978
rect 543554 3922 543622 3978
rect 543678 3922 561250 3978
rect 561306 3922 561374 3978
rect 561430 3922 561498 3978
rect 561554 3922 561622 3978
rect 561678 3922 579250 3978
rect 579306 3922 579374 3978
rect 579430 3922 579498 3978
rect 579554 3922 579622 3978
rect 579678 3922 596496 3978
rect 596552 3922 596620 3978
rect 596676 3922 596744 3978
rect 596800 3922 596868 3978
rect 596924 3922 597980 3978
rect -1916 3826 597980 3922
rect -956 -160 597020 -64
rect -956 -216 -860 -160
rect -804 -216 -736 -160
rect -680 -216 -612 -160
rect -556 -216 -488 -160
rect -432 -216 3250 -160
rect 3306 -216 3374 -160
rect 3430 -216 3498 -160
rect 3554 -216 3622 -160
rect 3678 -216 21250 -160
rect 21306 -216 21374 -160
rect 21430 -216 21498 -160
rect 21554 -216 21622 -160
rect 21678 -216 39250 -160
rect 39306 -216 39374 -160
rect 39430 -216 39498 -160
rect 39554 -216 39622 -160
rect 39678 -216 57250 -160
rect 57306 -216 57374 -160
rect 57430 -216 57498 -160
rect 57554 -216 57622 -160
rect 57678 -216 75250 -160
rect 75306 -216 75374 -160
rect 75430 -216 75498 -160
rect 75554 -216 75622 -160
rect 75678 -216 93250 -160
rect 93306 -216 93374 -160
rect 93430 -216 93498 -160
rect 93554 -216 93622 -160
rect 93678 -216 111250 -160
rect 111306 -216 111374 -160
rect 111430 -216 111498 -160
rect 111554 -216 111622 -160
rect 111678 -216 129250 -160
rect 129306 -216 129374 -160
rect 129430 -216 129498 -160
rect 129554 -216 129622 -160
rect 129678 -216 147250 -160
rect 147306 -216 147374 -160
rect 147430 -216 147498 -160
rect 147554 -216 147622 -160
rect 147678 -216 165250 -160
rect 165306 -216 165374 -160
rect 165430 -216 165498 -160
rect 165554 -216 165622 -160
rect 165678 -216 183250 -160
rect 183306 -216 183374 -160
rect 183430 -216 183498 -160
rect 183554 -216 183622 -160
rect 183678 -216 201250 -160
rect 201306 -216 201374 -160
rect 201430 -216 201498 -160
rect 201554 -216 201622 -160
rect 201678 -216 219250 -160
rect 219306 -216 219374 -160
rect 219430 -216 219498 -160
rect 219554 -216 219622 -160
rect 219678 -216 237250 -160
rect 237306 -216 237374 -160
rect 237430 -216 237498 -160
rect 237554 -216 237622 -160
rect 237678 -216 255250 -160
rect 255306 -216 255374 -160
rect 255430 -216 255498 -160
rect 255554 -216 255622 -160
rect 255678 -216 273250 -160
rect 273306 -216 273374 -160
rect 273430 -216 273498 -160
rect 273554 -216 273622 -160
rect 273678 -216 291250 -160
rect 291306 -216 291374 -160
rect 291430 -216 291498 -160
rect 291554 -216 291622 -160
rect 291678 -216 309250 -160
rect 309306 -216 309374 -160
rect 309430 -216 309498 -160
rect 309554 -216 309622 -160
rect 309678 -216 327250 -160
rect 327306 -216 327374 -160
rect 327430 -216 327498 -160
rect 327554 -216 327622 -160
rect 327678 -216 345250 -160
rect 345306 -216 345374 -160
rect 345430 -216 345498 -160
rect 345554 -216 345622 -160
rect 345678 -216 363250 -160
rect 363306 -216 363374 -160
rect 363430 -216 363498 -160
rect 363554 -216 363622 -160
rect 363678 -216 381250 -160
rect 381306 -216 381374 -160
rect 381430 -216 381498 -160
rect 381554 -216 381622 -160
rect 381678 -216 399250 -160
rect 399306 -216 399374 -160
rect 399430 -216 399498 -160
rect 399554 -216 399622 -160
rect 399678 -216 417250 -160
rect 417306 -216 417374 -160
rect 417430 -216 417498 -160
rect 417554 -216 417622 -160
rect 417678 -216 435250 -160
rect 435306 -216 435374 -160
rect 435430 -216 435498 -160
rect 435554 -216 435622 -160
rect 435678 -216 453250 -160
rect 453306 -216 453374 -160
rect 453430 -216 453498 -160
rect 453554 -216 453622 -160
rect 453678 -216 471250 -160
rect 471306 -216 471374 -160
rect 471430 -216 471498 -160
rect 471554 -216 471622 -160
rect 471678 -216 489250 -160
rect 489306 -216 489374 -160
rect 489430 -216 489498 -160
rect 489554 -216 489622 -160
rect 489678 -216 507250 -160
rect 507306 -216 507374 -160
rect 507430 -216 507498 -160
rect 507554 -216 507622 -160
rect 507678 -216 525250 -160
rect 525306 -216 525374 -160
rect 525430 -216 525498 -160
rect 525554 -216 525622 -160
rect 525678 -216 543250 -160
rect 543306 -216 543374 -160
rect 543430 -216 543498 -160
rect 543554 -216 543622 -160
rect 543678 -216 561250 -160
rect 561306 -216 561374 -160
rect 561430 -216 561498 -160
rect 561554 -216 561622 -160
rect 561678 -216 579250 -160
rect 579306 -216 579374 -160
rect 579430 -216 579498 -160
rect 579554 -216 579622 -160
rect 579678 -216 596496 -160
rect 596552 -216 596620 -160
rect 596676 -216 596744 -160
rect 596800 -216 596868 -160
rect 596924 -216 597020 -160
rect -956 -284 597020 -216
rect -956 -340 -860 -284
rect -804 -340 -736 -284
rect -680 -340 -612 -284
rect -556 -340 -488 -284
rect -432 -340 3250 -284
rect 3306 -340 3374 -284
rect 3430 -340 3498 -284
rect 3554 -340 3622 -284
rect 3678 -340 21250 -284
rect 21306 -340 21374 -284
rect 21430 -340 21498 -284
rect 21554 -340 21622 -284
rect 21678 -340 39250 -284
rect 39306 -340 39374 -284
rect 39430 -340 39498 -284
rect 39554 -340 39622 -284
rect 39678 -340 57250 -284
rect 57306 -340 57374 -284
rect 57430 -340 57498 -284
rect 57554 -340 57622 -284
rect 57678 -340 75250 -284
rect 75306 -340 75374 -284
rect 75430 -340 75498 -284
rect 75554 -340 75622 -284
rect 75678 -340 93250 -284
rect 93306 -340 93374 -284
rect 93430 -340 93498 -284
rect 93554 -340 93622 -284
rect 93678 -340 111250 -284
rect 111306 -340 111374 -284
rect 111430 -340 111498 -284
rect 111554 -340 111622 -284
rect 111678 -340 129250 -284
rect 129306 -340 129374 -284
rect 129430 -340 129498 -284
rect 129554 -340 129622 -284
rect 129678 -340 147250 -284
rect 147306 -340 147374 -284
rect 147430 -340 147498 -284
rect 147554 -340 147622 -284
rect 147678 -340 165250 -284
rect 165306 -340 165374 -284
rect 165430 -340 165498 -284
rect 165554 -340 165622 -284
rect 165678 -340 183250 -284
rect 183306 -340 183374 -284
rect 183430 -340 183498 -284
rect 183554 -340 183622 -284
rect 183678 -340 201250 -284
rect 201306 -340 201374 -284
rect 201430 -340 201498 -284
rect 201554 -340 201622 -284
rect 201678 -340 219250 -284
rect 219306 -340 219374 -284
rect 219430 -340 219498 -284
rect 219554 -340 219622 -284
rect 219678 -340 237250 -284
rect 237306 -340 237374 -284
rect 237430 -340 237498 -284
rect 237554 -340 237622 -284
rect 237678 -340 255250 -284
rect 255306 -340 255374 -284
rect 255430 -340 255498 -284
rect 255554 -340 255622 -284
rect 255678 -340 273250 -284
rect 273306 -340 273374 -284
rect 273430 -340 273498 -284
rect 273554 -340 273622 -284
rect 273678 -340 291250 -284
rect 291306 -340 291374 -284
rect 291430 -340 291498 -284
rect 291554 -340 291622 -284
rect 291678 -340 309250 -284
rect 309306 -340 309374 -284
rect 309430 -340 309498 -284
rect 309554 -340 309622 -284
rect 309678 -340 327250 -284
rect 327306 -340 327374 -284
rect 327430 -340 327498 -284
rect 327554 -340 327622 -284
rect 327678 -340 345250 -284
rect 345306 -340 345374 -284
rect 345430 -340 345498 -284
rect 345554 -340 345622 -284
rect 345678 -340 363250 -284
rect 363306 -340 363374 -284
rect 363430 -340 363498 -284
rect 363554 -340 363622 -284
rect 363678 -340 381250 -284
rect 381306 -340 381374 -284
rect 381430 -340 381498 -284
rect 381554 -340 381622 -284
rect 381678 -340 399250 -284
rect 399306 -340 399374 -284
rect 399430 -340 399498 -284
rect 399554 -340 399622 -284
rect 399678 -340 417250 -284
rect 417306 -340 417374 -284
rect 417430 -340 417498 -284
rect 417554 -340 417622 -284
rect 417678 -340 435250 -284
rect 435306 -340 435374 -284
rect 435430 -340 435498 -284
rect 435554 -340 435622 -284
rect 435678 -340 453250 -284
rect 453306 -340 453374 -284
rect 453430 -340 453498 -284
rect 453554 -340 453622 -284
rect 453678 -340 471250 -284
rect 471306 -340 471374 -284
rect 471430 -340 471498 -284
rect 471554 -340 471622 -284
rect 471678 -340 489250 -284
rect 489306 -340 489374 -284
rect 489430 -340 489498 -284
rect 489554 -340 489622 -284
rect 489678 -340 507250 -284
rect 507306 -340 507374 -284
rect 507430 -340 507498 -284
rect 507554 -340 507622 -284
rect 507678 -340 525250 -284
rect 525306 -340 525374 -284
rect 525430 -340 525498 -284
rect 525554 -340 525622 -284
rect 525678 -340 543250 -284
rect 543306 -340 543374 -284
rect 543430 -340 543498 -284
rect 543554 -340 543622 -284
rect 543678 -340 561250 -284
rect 561306 -340 561374 -284
rect 561430 -340 561498 -284
rect 561554 -340 561622 -284
rect 561678 -340 579250 -284
rect 579306 -340 579374 -284
rect 579430 -340 579498 -284
rect 579554 -340 579622 -284
rect 579678 -340 596496 -284
rect 596552 -340 596620 -284
rect 596676 -340 596744 -284
rect 596800 -340 596868 -284
rect 596924 -340 597020 -284
rect -956 -408 597020 -340
rect -956 -464 -860 -408
rect -804 -464 -736 -408
rect -680 -464 -612 -408
rect -556 -464 -488 -408
rect -432 -464 3250 -408
rect 3306 -464 3374 -408
rect 3430 -464 3498 -408
rect 3554 -464 3622 -408
rect 3678 -464 21250 -408
rect 21306 -464 21374 -408
rect 21430 -464 21498 -408
rect 21554 -464 21622 -408
rect 21678 -464 39250 -408
rect 39306 -464 39374 -408
rect 39430 -464 39498 -408
rect 39554 -464 39622 -408
rect 39678 -464 57250 -408
rect 57306 -464 57374 -408
rect 57430 -464 57498 -408
rect 57554 -464 57622 -408
rect 57678 -464 75250 -408
rect 75306 -464 75374 -408
rect 75430 -464 75498 -408
rect 75554 -464 75622 -408
rect 75678 -464 93250 -408
rect 93306 -464 93374 -408
rect 93430 -464 93498 -408
rect 93554 -464 93622 -408
rect 93678 -464 111250 -408
rect 111306 -464 111374 -408
rect 111430 -464 111498 -408
rect 111554 -464 111622 -408
rect 111678 -464 129250 -408
rect 129306 -464 129374 -408
rect 129430 -464 129498 -408
rect 129554 -464 129622 -408
rect 129678 -464 147250 -408
rect 147306 -464 147374 -408
rect 147430 -464 147498 -408
rect 147554 -464 147622 -408
rect 147678 -464 165250 -408
rect 165306 -464 165374 -408
rect 165430 -464 165498 -408
rect 165554 -464 165622 -408
rect 165678 -464 183250 -408
rect 183306 -464 183374 -408
rect 183430 -464 183498 -408
rect 183554 -464 183622 -408
rect 183678 -464 201250 -408
rect 201306 -464 201374 -408
rect 201430 -464 201498 -408
rect 201554 -464 201622 -408
rect 201678 -464 219250 -408
rect 219306 -464 219374 -408
rect 219430 -464 219498 -408
rect 219554 -464 219622 -408
rect 219678 -464 237250 -408
rect 237306 -464 237374 -408
rect 237430 -464 237498 -408
rect 237554 -464 237622 -408
rect 237678 -464 255250 -408
rect 255306 -464 255374 -408
rect 255430 -464 255498 -408
rect 255554 -464 255622 -408
rect 255678 -464 273250 -408
rect 273306 -464 273374 -408
rect 273430 -464 273498 -408
rect 273554 -464 273622 -408
rect 273678 -464 291250 -408
rect 291306 -464 291374 -408
rect 291430 -464 291498 -408
rect 291554 -464 291622 -408
rect 291678 -464 309250 -408
rect 309306 -464 309374 -408
rect 309430 -464 309498 -408
rect 309554 -464 309622 -408
rect 309678 -464 327250 -408
rect 327306 -464 327374 -408
rect 327430 -464 327498 -408
rect 327554 -464 327622 -408
rect 327678 -464 345250 -408
rect 345306 -464 345374 -408
rect 345430 -464 345498 -408
rect 345554 -464 345622 -408
rect 345678 -464 363250 -408
rect 363306 -464 363374 -408
rect 363430 -464 363498 -408
rect 363554 -464 363622 -408
rect 363678 -464 381250 -408
rect 381306 -464 381374 -408
rect 381430 -464 381498 -408
rect 381554 -464 381622 -408
rect 381678 -464 399250 -408
rect 399306 -464 399374 -408
rect 399430 -464 399498 -408
rect 399554 -464 399622 -408
rect 399678 -464 417250 -408
rect 417306 -464 417374 -408
rect 417430 -464 417498 -408
rect 417554 -464 417622 -408
rect 417678 -464 435250 -408
rect 435306 -464 435374 -408
rect 435430 -464 435498 -408
rect 435554 -464 435622 -408
rect 435678 -464 453250 -408
rect 453306 -464 453374 -408
rect 453430 -464 453498 -408
rect 453554 -464 453622 -408
rect 453678 -464 471250 -408
rect 471306 -464 471374 -408
rect 471430 -464 471498 -408
rect 471554 -464 471622 -408
rect 471678 -464 489250 -408
rect 489306 -464 489374 -408
rect 489430 -464 489498 -408
rect 489554 -464 489622 -408
rect 489678 -464 507250 -408
rect 507306 -464 507374 -408
rect 507430 -464 507498 -408
rect 507554 -464 507622 -408
rect 507678 -464 525250 -408
rect 525306 -464 525374 -408
rect 525430 -464 525498 -408
rect 525554 -464 525622 -408
rect 525678 -464 543250 -408
rect 543306 -464 543374 -408
rect 543430 -464 543498 -408
rect 543554 -464 543622 -408
rect 543678 -464 561250 -408
rect 561306 -464 561374 -408
rect 561430 -464 561498 -408
rect 561554 -464 561622 -408
rect 561678 -464 579250 -408
rect 579306 -464 579374 -408
rect 579430 -464 579498 -408
rect 579554 -464 579622 -408
rect 579678 -464 596496 -408
rect 596552 -464 596620 -408
rect 596676 -464 596744 -408
rect 596800 -464 596868 -408
rect 596924 -464 597020 -408
rect -956 -532 597020 -464
rect -956 -588 -860 -532
rect -804 -588 -736 -532
rect -680 -588 -612 -532
rect -556 -588 -488 -532
rect -432 -588 3250 -532
rect 3306 -588 3374 -532
rect 3430 -588 3498 -532
rect 3554 -588 3622 -532
rect 3678 -588 21250 -532
rect 21306 -588 21374 -532
rect 21430 -588 21498 -532
rect 21554 -588 21622 -532
rect 21678 -588 39250 -532
rect 39306 -588 39374 -532
rect 39430 -588 39498 -532
rect 39554 -588 39622 -532
rect 39678 -588 57250 -532
rect 57306 -588 57374 -532
rect 57430 -588 57498 -532
rect 57554 -588 57622 -532
rect 57678 -588 75250 -532
rect 75306 -588 75374 -532
rect 75430 -588 75498 -532
rect 75554 -588 75622 -532
rect 75678 -588 93250 -532
rect 93306 -588 93374 -532
rect 93430 -588 93498 -532
rect 93554 -588 93622 -532
rect 93678 -588 111250 -532
rect 111306 -588 111374 -532
rect 111430 -588 111498 -532
rect 111554 -588 111622 -532
rect 111678 -588 129250 -532
rect 129306 -588 129374 -532
rect 129430 -588 129498 -532
rect 129554 -588 129622 -532
rect 129678 -588 147250 -532
rect 147306 -588 147374 -532
rect 147430 -588 147498 -532
rect 147554 -588 147622 -532
rect 147678 -588 165250 -532
rect 165306 -588 165374 -532
rect 165430 -588 165498 -532
rect 165554 -588 165622 -532
rect 165678 -588 183250 -532
rect 183306 -588 183374 -532
rect 183430 -588 183498 -532
rect 183554 -588 183622 -532
rect 183678 -588 201250 -532
rect 201306 -588 201374 -532
rect 201430 -588 201498 -532
rect 201554 -588 201622 -532
rect 201678 -588 219250 -532
rect 219306 -588 219374 -532
rect 219430 -588 219498 -532
rect 219554 -588 219622 -532
rect 219678 -588 237250 -532
rect 237306 -588 237374 -532
rect 237430 -588 237498 -532
rect 237554 -588 237622 -532
rect 237678 -588 255250 -532
rect 255306 -588 255374 -532
rect 255430 -588 255498 -532
rect 255554 -588 255622 -532
rect 255678 -588 273250 -532
rect 273306 -588 273374 -532
rect 273430 -588 273498 -532
rect 273554 -588 273622 -532
rect 273678 -588 291250 -532
rect 291306 -588 291374 -532
rect 291430 -588 291498 -532
rect 291554 -588 291622 -532
rect 291678 -588 309250 -532
rect 309306 -588 309374 -532
rect 309430 -588 309498 -532
rect 309554 -588 309622 -532
rect 309678 -588 327250 -532
rect 327306 -588 327374 -532
rect 327430 -588 327498 -532
rect 327554 -588 327622 -532
rect 327678 -588 345250 -532
rect 345306 -588 345374 -532
rect 345430 -588 345498 -532
rect 345554 -588 345622 -532
rect 345678 -588 363250 -532
rect 363306 -588 363374 -532
rect 363430 -588 363498 -532
rect 363554 -588 363622 -532
rect 363678 -588 381250 -532
rect 381306 -588 381374 -532
rect 381430 -588 381498 -532
rect 381554 -588 381622 -532
rect 381678 -588 399250 -532
rect 399306 -588 399374 -532
rect 399430 -588 399498 -532
rect 399554 -588 399622 -532
rect 399678 -588 417250 -532
rect 417306 -588 417374 -532
rect 417430 -588 417498 -532
rect 417554 -588 417622 -532
rect 417678 -588 435250 -532
rect 435306 -588 435374 -532
rect 435430 -588 435498 -532
rect 435554 -588 435622 -532
rect 435678 -588 453250 -532
rect 453306 -588 453374 -532
rect 453430 -588 453498 -532
rect 453554 -588 453622 -532
rect 453678 -588 471250 -532
rect 471306 -588 471374 -532
rect 471430 -588 471498 -532
rect 471554 -588 471622 -532
rect 471678 -588 489250 -532
rect 489306 -588 489374 -532
rect 489430 -588 489498 -532
rect 489554 -588 489622 -532
rect 489678 -588 507250 -532
rect 507306 -588 507374 -532
rect 507430 -588 507498 -532
rect 507554 -588 507622 -532
rect 507678 -588 525250 -532
rect 525306 -588 525374 -532
rect 525430 -588 525498 -532
rect 525554 -588 525622 -532
rect 525678 -588 543250 -532
rect 543306 -588 543374 -532
rect 543430 -588 543498 -532
rect 543554 -588 543622 -532
rect 543678 -588 561250 -532
rect 561306 -588 561374 -532
rect 561430 -588 561498 -532
rect 561554 -588 561622 -532
rect 561678 -588 579250 -532
rect 579306 -588 579374 -532
rect 579430 -588 579498 -532
rect 579554 -588 579622 -532
rect 579678 -588 596496 -532
rect 596552 -588 596620 -532
rect 596676 -588 596744 -532
rect 596800 -588 596868 -532
rect 596924 -588 597020 -532
rect -956 -684 597020 -588
rect -1916 -1120 597980 -1024
rect -1916 -1176 -1820 -1120
rect -1764 -1176 -1696 -1120
rect -1640 -1176 -1572 -1120
rect -1516 -1176 -1448 -1120
rect -1392 -1176 6970 -1120
rect 7026 -1176 7094 -1120
rect 7150 -1176 7218 -1120
rect 7274 -1176 7342 -1120
rect 7398 -1176 24970 -1120
rect 25026 -1176 25094 -1120
rect 25150 -1176 25218 -1120
rect 25274 -1176 25342 -1120
rect 25398 -1176 42970 -1120
rect 43026 -1176 43094 -1120
rect 43150 -1176 43218 -1120
rect 43274 -1176 43342 -1120
rect 43398 -1176 60970 -1120
rect 61026 -1176 61094 -1120
rect 61150 -1176 61218 -1120
rect 61274 -1176 61342 -1120
rect 61398 -1176 78970 -1120
rect 79026 -1176 79094 -1120
rect 79150 -1176 79218 -1120
rect 79274 -1176 79342 -1120
rect 79398 -1176 96970 -1120
rect 97026 -1176 97094 -1120
rect 97150 -1176 97218 -1120
rect 97274 -1176 97342 -1120
rect 97398 -1176 114970 -1120
rect 115026 -1176 115094 -1120
rect 115150 -1176 115218 -1120
rect 115274 -1176 115342 -1120
rect 115398 -1176 132970 -1120
rect 133026 -1176 133094 -1120
rect 133150 -1176 133218 -1120
rect 133274 -1176 133342 -1120
rect 133398 -1176 150970 -1120
rect 151026 -1176 151094 -1120
rect 151150 -1176 151218 -1120
rect 151274 -1176 151342 -1120
rect 151398 -1176 168970 -1120
rect 169026 -1176 169094 -1120
rect 169150 -1176 169218 -1120
rect 169274 -1176 169342 -1120
rect 169398 -1176 186970 -1120
rect 187026 -1176 187094 -1120
rect 187150 -1176 187218 -1120
rect 187274 -1176 187342 -1120
rect 187398 -1176 204970 -1120
rect 205026 -1176 205094 -1120
rect 205150 -1176 205218 -1120
rect 205274 -1176 205342 -1120
rect 205398 -1176 384970 -1120
rect 385026 -1176 385094 -1120
rect 385150 -1176 385218 -1120
rect 385274 -1176 385342 -1120
rect 385398 -1176 402970 -1120
rect 403026 -1176 403094 -1120
rect 403150 -1176 403218 -1120
rect 403274 -1176 403342 -1120
rect 403398 -1176 420970 -1120
rect 421026 -1176 421094 -1120
rect 421150 -1176 421218 -1120
rect 421274 -1176 421342 -1120
rect 421398 -1176 438970 -1120
rect 439026 -1176 439094 -1120
rect 439150 -1176 439218 -1120
rect 439274 -1176 439342 -1120
rect 439398 -1176 456970 -1120
rect 457026 -1176 457094 -1120
rect 457150 -1176 457218 -1120
rect 457274 -1176 457342 -1120
rect 457398 -1176 474970 -1120
rect 475026 -1176 475094 -1120
rect 475150 -1176 475218 -1120
rect 475274 -1176 475342 -1120
rect 475398 -1176 492970 -1120
rect 493026 -1176 493094 -1120
rect 493150 -1176 493218 -1120
rect 493274 -1176 493342 -1120
rect 493398 -1176 510970 -1120
rect 511026 -1176 511094 -1120
rect 511150 -1176 511218 -1120
rect 511274 -1176 511342 -1120
rect 511398 -1176 528970 -1120
rect 529026 -1176 529094 -1120
rect 529150 -1176 529218 -1120
rect 529274 -1176 529342 -1120
rect 529398 -1176 546970 -1120
rect 547026 -1176 547094 -1120
rect 547150 -1176 547218 -1120
rect 547274 -1176 547342 -1120
rect 547398 -1176 564970 -1120
rect 565026 -1176 565094 -1120
rect 565150 -1176 565218 -1120
rect 565274 -1176 565342 -1120
rect 565398 -1176 582970 -1120
rect 583026 -1176 583094 -1120
rect 583150 -1176 583218 -1120
rect 583274 -1176 583342 -1120
rect 583398 -1176 597456 -1120
rect 597512 -1176 597580 -1120
rect 597636 -1176 597704 -1120
rect 597760 -1176 597828 -1120
rect 597884 -1176 597980 -1120
rect -1916 -1244 597980 -1176
rect -1916 -1300 -1820 -1244
rect -1764 -1300 -1696 -1244
rect -1640 -1300 -1572 -1244
rect -1516 -1300 -1448 -1244
rect -1392 -1300 6970 -1244
rect 7026 -1300 7094 -1244
rect 7150 -1300 7218 -1244
rect 7274 -1300 7342 -1244
rect 7398 -1300 24970 -1244
rect 25026 -1300 25094 -1244
rect 25150 -1300 25218 -1244
rect 25274 -1300 25342 -1244
rect 25398 -1300 42970 -1244
rect 43026 -1300 43094 -1244
rect 43150 -1300 43218 -1244
rect 43274 -1300 43342 -1244
rect 43398 -1300 60970 -1244
rect 61026 -1300 61094 -1244
rect 61150 -1300 61218 -1244
rect 61274 -1300 61342 -1244
rect 61398 -1300 78970 -1244
rect 79026 -1300 79094 -1244
rect 79150 -1300 79218 -1244
rect 79274 -1300 79342 -1244
rect 79398 -1300 96970 -1244
rect 97026 -1300 97094 -1244
rect 97150 -1300 97218 -1244
rect 97274 -1300 97342 -1244
rect 97398 -1300 114970 -1244
rect 115026 -1300 115094 -1244
rect 115150 -1300 115218 -1244
rect 115274 -1300 115342 -1244
rect 115398 -1300 132970 -1244
rect 133026 -1300 133094 -1244
rect 133150 -1300 133218 -1244
rect 133274 -1300 133342 -1244
rect 133398 -1300 150970 -1244
rect 151026 -1300 151094 -1244
rect 151150 -1300 151218 -1244
rect 151274 -1300 151342 -1244
rect 151398 -1300 168970 -1244
rect 169026 -1300 169094 -1244
rect 169150 -1300 169218 -1244
rect 169274 -1300 169342 -1244
rect 169398 -1300 186970 -1244
rect 187026 -1300 187094 -1244
rect 187150 -1300 187218 -1244
rect 187274 -1300 187342 -1244
rect 187398 -1300 204970 -1244
rect 205026 -1300 205094 -1244
rect 205150 -1300 205218 -1244
rect 205274 -1300 205342 -1244
rect 205398 -1300 384970 -1244
rect 385026 -1300 385094 -1244
rect 385150 -1300 385218 -1244
rect 385274 -1300 385342 -1244
rect 385398 -1300 402970 -1244
rect 403026 -1300 403094 -1244
rect 403150 -1300 403218 -1244
rect 403274 -1300 403342 -1244
rect 403398 -1300 420970 -1244
rect 421026 -1300 421094 -1244
rect 421150 -1300 421218 -1244
rect 421274 -1300 421342 -1244
rect 421398 -1300 438970 -1244
rect 439026 -1300 439094 -1244
rect 439150 -1300 439218 -1244
rect 439274 -1300 439342 -1244
rect 439398 -1300 456970 -1244
rect 457026 -1300 457094 -1244
rect 457150 -1300 457218 -1244
rect 457274 -1300 457342 -1244
rect 457398 -1300 474970 -1244
rect 475026 -1300 475094 -1244
rect 475150 -1300 475218 -1244
rect 475274 -1300 475342 -1244
rect 475398 -1300 492970 -1244
rect 493026 -1300 493094 -1244
rect 493150 -1300 493218 -1244
rect 493274 -1300 493342 -1244
rect 493398 -1300 510970 -1244
rect 511026 -1300 511094 -1244
rect 511150 -1300 511218 -1244
rect 511274 -1300 511342 -1244
rect 511398 -1300 528970 -1244
rect 529026 -1300 529094 -1244
rect 529150 -1300 529218 -1244
rect 529274 -1300 529342 -1244
rect 529398 -1300 546970 -1244
rect 547026 -1300 547094 -1244
rect 547150 -1300 547218 -1244
rect 547274 -1300 547342 -1244
rect 547398 -1300 564970 -1244
rect 565026 -1300 565094 -1244
rect 565150 -1300 565218 -1244
rect 565274 -1300 565342 -1244
rect 565398 -1300 582970 -1244
rect 583026 -1300 583094 -1244
rect 583150 -1300 583218 -1244
rect 583274 -1300 583342 -1244
rect 583398 -1300 597456 -1244
rect 597512 -1300 597580 -1244
rect 597636 -1300 597704 -1244
rect 597760 -1300 597828 -1244
rect 597884 -1300 597980 -1244
rect -1916 -1368 597980 -1300
rect -1916 -1424 -1820 -1368
rect -1764 -1424 -1696 -1368
rect -1640 -1424 -1572 -1368
rect -1516 -1424 -1448 -1368
rect -1392 -1424 6970 -1368
rect 7026 -1424 7094 -1368
rect 7150 -1424 7218 -1368
rect 7274 -1424 7342 -1368
rect 7398 -1424 24970 -1368
rect 25026 -1424 25094 -1368
rect 25150 -1424 25218 -1368
rect 25274 -1424 25342 -1368
rect 25398 -1424 42970 -1368
rect 43026 -1424 43094 -1368
rect 43150 -1424 43218 -1368
rect 43274 -1424 43342 -1368
rect 43398 -1424 60970 -1368
rect 61026 -1424 61094 -1368
rect 61150 -1424 61218 -1368
rect 61274 -1424 61342 -1368
rect 61398 -1424 78970 -1368
rect 79026 -1424 79094 -1368
rect 79150 -1424 79218 -1368
rect 79274 -1424 79342 -1368
rect 79398 -1424 96970 -1368
rect 97026 -1424 97094 -1368
rect 97150 -1424 97218 -1368
rect 97274 -1424 97342 -1368
rect 97398 -1424 114970 -1368
rect 115026 -1424 115094 -1368
rect 115150 -1424 115218 -1368
rect 115274 -1424 115342 -1368
rect 115398 -1424 132970 -1368
rect 133026 -1424 133094 -1368
rect 133150 -1424 133218 -1368
rect 133274 -1424 133342 -1368
rect 133398 -1424 150970 -1368
rect 151026 -1424 151094 -1368
rect 151150 -1424 151218 -1368
rect 151274 -1424 151342 -1368
rect 151398 -1424 168970 -1368
rect 169026 -1424 169094 -1368
rect 169150 -1424 169218 -1368
rect 169274 -1424 169342 -1368
rect 169398 -1424 186970 -1368
rect 187026 -1424 187094 -1368
rect 187150 -1424 187218 -1368
rect 187274 -1424 187342 -1368
rect 187398 -1424 204970 -1368
rect 205026 -1424 205094 -1368
rect 205150 -1424 205218 -1368
rect 205274 -1424 205342 -1368
rect 205398 -1424 384970 -1368
rect 385026 -1424 385094 -1368
rect 385150 -1424 385218 -1368
rect 385274 -1424 385342 -1368
rect 385398 -1424 402970 -1368
rect 403026 -1424 403094 -1368
rect 403150 -1424 403218 -1368
rect 403274 -1424 403342 -1368
rect 403398 -1424 420970 -1368
rect 421026 -1424 421094 -1368
rect 421150 -1424 421218 -1368
rect 421274 -1424 421342 -1368
rect 421398 -1424 438970 -1368
rect 439026 -1424 439094 -1368
rect 439150 -1424 439218 -1368
rect 439274 -1424 439342 -1368
rect 439398 -1424 456970 -1368
rect 457026 -1424 457094 -1368
rect 457150 -1424 457218 -1368
rect 457274 -1424 457342 -1368
rect 457398 -1424 474970 -1368
rect 475026 -1424 475094 -1368
rect 475150 -1424 475218 -1368
rect 475274 -1424 475342 -1368
rect 475398 -1424 492970 -1368
rect 493026 -1424 493094 -1368
rect 493150 -1424 493218 -1368
rect 493274 -1424 493342 -1368
rect 493398 -1424 510970 -1368
rect 511026 -1424 511094 -1368
rect 511150 -1424 511218 -1368
rect 511274 -1424 511342 -1368
rect 511398 -1424 528970 -1368
rect 529026 -1424 529094 -1368
rect 529150 -1424 529218 -1368
rect 529274 -1424 529342 -1368
rect 529398 -1424 546970 -1368
rect 547026 -1424 547094 -1368
rect 547150 -1424 547218 -1368
rect 547274 -1424 547342 -1368
rect 547398 -1424 564970 -1368
rect 565026 -1424 565094 -1368
rect 565150 -1424 565218 -1368
rect 565274 -1424 565342 -1368
rect 565398 -1424 582970 -1368
rect 583026 -1424 583094 -1368
rect 583150 -1424 583218 -1368
rect 583274 -1424 583342 -1368
rect 583398 -1424 597456 -1368
rect 597512 -1424 597580 -1368
rect 597636 -1424 597704 -1368
rect 597760 -1424 597828 -1368
rect 597884 -1424 597980 -1368
rect -1916 -1492 597980 -1424
rect -1916 -1548 -1820 -1492
rect -1764 -1548 -1696 -1492
rect -1640 -1548 -1572 -1492
rect -1516 -1548 -1448 -1492
rect -1392 -1548 6970 -1492
rect 7026 -1548 7094 -1492
rect 7150 -1548 7218 -1492
rect 7274 -1548 7342 -1492
rect 7398 -1548 24970 -1492
rect 25026 -1548 25094 -1492
rect 25150 -1548 25218 -1492
rect 25274 -1548 25342 -1492
rect 25398 -1548 42970 -1492
rect 43026 -1548 43094 -1492
rect 43150 -1548 43218 -1492
rect 43274 -1548 43342 -1492
rect 43398 -1548 60970 -1492
rect 61026 -1548 61094 -1492
rect 61150 -1548 61218 -1492
rect 61274 -1548 61342 -1492
rect 61398 -1548 78970 -1492
rect 79026 -1548 79094 -1492
rect 79150 -1548 79218 -1492
rect 79274 -1548 79342 -1492
rect 79398 -1548 96970 -1492
rect 97026 -1548 97094 -1492
rect 97150 -1548 97218 -1492
rect 97274 -1548 97342 -1492
rect 97398 -1548 114970 -1492
rect 115026 -1548 115094 -1492
rect 115150 -1548 115218 -1492
rect 115274 -1548 115342 -1492
rect 115398 -1548 132970 -1492
rect 133026 -1548 133094 -1492
rect 133150 -1548 133218 -1492
rect 133274 -1548 133342 -1492
rect 133398 -1548 150970 -1492
rect 151026 -1548 151094 -1492
rect 151150 -1548 151218 -1492
rect 151274 -1548 151342 -1492
rect 151398 -1548 168970 -1492
rect 169026 -1548 169094 -1492
rect 169150 -1548 169218 -1492
rect 169274 -1548 169342 -1492
rect 169398 -1548 186970 -1492
rect 187026 -1548 187094 -1492
rect 187150 -1548 187218 -1492
rect 187274 -1548 187342 -1492
rect 187398 -1548 204970 -1492
rect 205026 -1548 205094 -1492
rect 205150 -1548 205218 -1492
rect 205274 -1548 205342 -1492
rect 205398 -1548 384970 -1492
rect 385026 -1548 385094 -1492
rect 385150 -1548 385218 -1492
rect 385274 -1548 385342 -1492
rect 385398 -1548 402970 -1492
rect 403026 -1548 403094 -1492
rect 403150 -1548 403218 -1492
rect 403274 -1548 403342 -1492
rect 403398 -1548 420970 -1492
rect 421026 -1548 421094 -1492
rect 421150 -1548 421218 -1492
rect 421274 -1548 421342 -1492
rect 421398 -1548 438970 -1492
rect 439026 -1548 439094 -1492
rect 439150 -1548 439218 -1492
rect 439274 -1548 439342 -1492
rect 439398 -1548 456970 -1492
rect 457026 -1548 457094 -1492
rect 457150 -1548 457218 -1492
rect 457274 -1548 457342 -1492
rect 457398 -1548 474970 -1492
rect 475026 -1548 475094 -1492
rect 475150 -1548 475218 -1492
rect 475274 -1548 475342 -1492
rect 475398 -1548 492970 -1492
rect 493026 -1548 493094 -1492
rect 493150 -1548 493218 -1492
rect 493274 -1548 493342 -1492
rect 493398 -1548 510970 -1492
rect 511026 -1548 511094 -1492
rect 511150 -1548 511218 -1492
rect 511274 -1548 511342 -1492
rect 511398 -1548 528970 -1492
rect 529026 -1548 529094 -1492
rect 529150 -1548 529218 -1492
rect 529274 -1548 529342 -1492
rect 529398 -1548 546970 -1492
rect 547026 -1548 547094 -1492
rect 547150 -1548 547218 -1492
rect 547274 -1548 547342 -1492
rect 547398 -1548 564970 -1492
rect 565026 -1548 565094 -1492
rect 565150 -1548 565218 -1492
rect 565274 -1548 565342 -1492
rect 565398 -1548 582970 -1492
rect 583026 -1548 583094 -1492
rect 583150 -1548 583218 -1492
rect 583274 -1548 583342 -1492
rect 583398 -1548 597456 -1492
rect 597512 -1548 597580 -1492
rect 597636 -1548 597704 -1492
rect 597760 -1548 597828 -1492
rect 597884 -1548 597980 -1492
rect -1916 -1644 597980 -1548
use clock_mux  clock_mux_mod
timestamp 0
transform 1 0 520000 0 1 60000
box 0 0 50000 46316
use controller_core  controller_core_mod
timestamp 0
transform 1 0 21600 0 1 70000
box 0 0 158798 46000
use driver_core  driver_core_0
timestamp 0
transform 1 0 198000 0 1 10000
box 1344 0 178958 140396
use driver_core  driver_core_1
timestamp 0
transform 1 0 9000 0 1 160000
box 1344 0 178958 140396
use driver_core  driver_core_2
timestamp 0
transform 1 0 198000 0 1 160000
box 1344 0 178958 140396
use driver_core  driver_core_3
timestamp 0
transform 1 0 9000 0 1 320000
box 1344 0 178958 140396
use driver_core  driver_core_4
timestamp 0
transform 1 0 198000 0 1 320000
box 1344 0 178958 140396
use driver_core  driver_core_8
timestamp 0
transform 1 0 399000 0 1 320000
box 1344 0 178958 140396
use driver_core  driver_core_9
timestamp 0
transform 1 0 399000 0 1 160000
box 1344 0 178958 140396
use spi_core  spi_core_mod
timestamp 0
transform 1 0 12000 0 1 20000
box 0 0 50000 48272
<< labels >>
flabel metal3 s 591560 240408 593000 240632 0 FreeSans 896 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 451192 591560 451416 593000 0 FreeSans 896 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 385784 591560 386008 593000 0 FreeSans 896 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 320376 591560 320600 593000 0 FreeSans 896 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 254968 591560 255192 593000 0 FreeSans 896 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 189560 591560 189784 593000 0 FreeSans 896 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 124152 591560 124376 593000 0 FreeSans 896 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 58744 591560 58968 593000 0 FreeSans 896 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 583800 480 584024 0 FreeSans 896 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 540344 480 540568 0 FreeSans 896 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 496888 480 497112 0 FreeSans 896 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 591560 284760 593000 284984 0 FreeSans 896 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 453432 480 453656 0 FreeSans 896 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 409976 480 410200 0 FreeSans 896 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 366520 480 366744 0 FreeSans 896 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 323064 480 323288 0 FreeSans 896 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 279608 480 279832 0 FreeSans 896 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 236152 480 236376 0 FreeSans 896 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 192696 480 192920 0 FreeSans 896 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 149240 480 149464 0 FreeSans 896 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 105784 480 106008 0 FreeSans 896 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 591560 329112 593000 329336 0 FreeSans 896 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 591560 373464 593000 373688 0 FreeSans 896 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 591560 417816 593000 418040 0 FreeSans 896 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 591560 462168 593000 462392 0 FreeSans 896 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 591560 506520 593000 506744 0 FreeSans 896 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 591560 550872 593000 551096 0 FreeSans 896 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 582008 591560 582232 593000 0 FreeSans 896 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 516600 591560 516824 593000 0 FreeSans 896 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 591560 7560 593000 7784 0 FreeSans 896 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 591560 384552 593000 384776 0 FreeSans 896 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 591560 428904 593000 429128 0 FreeSans 896 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 591560 473256 593000 473480 0 FreeSans 896 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 591560 517608 593000 517832 0 FreeSans 896 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 591560 561960 593000 562184 0 FreeSans 896 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 565656 591560 565880 593000 0 FreeSans 896 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 500248 591560 500472 593000 0 FreeSans 896 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 434840 591560 435064 593000 0 FreeSans 896 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 369432 591560 369656 593000 0 FreeSans 896 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 304024 591560 304248 593000 0 FreeSans 896 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 591560 40824 593000 41048 0 FreeSans 896 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 238616 591560 238840 593000 0 FreeSans 896 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 173208 591560 173432 593000 0 FreeSans 896 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 107800 591560 108024 593000 0 FreeSans 896 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 42392 591560 42616 593000 0 FreeSans 896 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 572936 480 573160 0 FreeSans 896 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 529480 480 529704 0 FreeSans 896 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 486024 480 486248 0 FreeSans 896 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 442568 480 442792 0 FreeSans 896 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 399112 480 399336 0 FreeSans 896 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 355656 480 355880 0 FreeSans 896 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 591560 74088 593000 74312 0 FreeSans 896 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 312200 480 312424 0 FreeSans 896 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 268744 480 268968 0 FreeSans 896 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 225288 480 225512 0 FreeSans 896 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 181832 480 182056 0 FreeSans 896 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 138376 480 138600 0 FreeSans 896 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 94920 480 95144 0 FreeSans 896 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 62328 480 62552 0 FreeSans 896 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 29736 480 29960 0 FreeSans 896 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 591560 107352 593000 107576 0 FreeSans 896 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 591560 140616 593000 140840 0 FreeSans 896 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 591560 173880 593000 174104 0 FreeSans 896 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 591560 207144 593000 207368 0 FreeSans 896 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 591560 251496 593000 251720 0 FreeSans 896 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 591560 295848 593000 296072 0 FreeSans 896 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 591560 340200 593000 340424 0 FreeSans 896 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 591560 29736 593000 29960 0 FreeSans 896 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 591560 406728 593000 406952 0 FreeSans 896 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 591560 451080 593000 451304 0 FreeSans 896 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 591560 495432 593000 495656 0 FreeSans 896 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 591560 539784 593000 540008 0 FreeSans 896 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 591560 584136 593000 584360 0 FreeSans 896 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 532952 591560 533176 593000 0 FreeSans 896 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 467544 591560 467768 593000 0 FreeSans 896 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 402136 591560 402360 593000 0 FreeSans 896 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 336728 591560 336952 593000 0 FreeSans 896 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 271320 591560 271544 593000 0 FreeSans 896 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 591560 63000 593000 63224 0 FreeSans 896 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 205912 591560 206136 593000 0 FreeSans 896 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 140504 591560 140728 593000 0 FreeSans 896 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 75096 591560 75320 593000 0 FreeSans 896 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 9688 591560 9912 593000 0 FreeSans 896 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 551208 480 551432 0 FreeSans 896 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 507752 480 507976 0 FreeSans 896 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 464296 480 464520 0 FreeSans 896 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 420840 480 421064 0 FreeSans 896 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 377384 480 377608 0 FreeSans 896 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 333928 480 334152 0 FreeSans 896 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 591560 96264 593000 96488 0 FreeSans 896 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 290472 480 290696 0 FreeSans 896 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 247016 480 247240 0 FreeSans 896 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 203560 480 203784 0 FreeSans 896 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 160104 480 160328 0 FreeSans 896 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 116648 480 116872 0 FreeSans 896 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 73192 480 73416 0 FreeSans 896 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 40600 480 40824 0 FreeSans 896 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 8008 480 8232 0 FreeSans 896 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 591560 129528 593000 129752 0 FreeSans 896 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 591560 162792 593000 163016 0 FreeSans 896 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 591560 196056 593000 196280 0 FreeSans 896 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 591560 229320 593000 229544 0 FreeSans 896 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 591560 273672 593000 273896 0 FreeSans 896 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 591560 318024 593000 318248 0 FreeSans 896 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 591560 362376 593000 362600 0 FreeSans 896 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 591560 18648 593000 18872 0 FreeSans 896 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 591560 395640 593000 395864 0 FreeSans 896 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 591560 439992 593000 440216 0 FreeSans 896 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 591560 484344 593000 484568 0 FreeSans 896 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 591560 528696 593000 528920 0 FreeSans 896 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 591560 573048 593000 573272 0 FreeSans 896 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 549304 591560 549528 593000 0 FreeSans 896 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 483896 591560 484120 593000 0 FreeSans 896 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 418488 591560 418712 593000 0 FreeSans 896 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 353080 591560 353304 593000 0 FreeSans 896 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 287672 591560 287896 593000 0 FreeSans 896 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 591560 51912 593000 52136 0 FreeSans 896 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 222264 591560 222488 593000 0 FreeSans 896 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 156856 591560 157080 593000 0 FreeSans 896 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 91448 591560 91672 593000 0 FreeSans 896 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 26040 591560 26264 593000 0 FreeSans 896 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 562072 480 562296 0 FreeSans 896 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 518616 480 518840 0 FreeSans 896 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 475160 480 475384 0 FreeSans 896 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 431704 480 431928 0 FreeSans 896 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 388248 480 388472 0 FreeSans 896 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 344792 480 345016 0 FreeSans 896 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 591560 85176 593000 85400 0 FreeSans 896 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 301336 480 301560 0 FreeSans 896 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 257880 480 258104 0 FreeSans 896 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 214424 480 214648 0 FreeSans 896 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 170968 480 171192 0 FreeSans 896 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 127512 480 127736 0 FreeSans 896 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 84056 480 84280 0 FreeSans 896 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 51464 480 51688 0 FreeSans 896 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 18872 480 19096 0 FreeSans 896 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 591560 118440 593000 118664 0 FreeSans 896 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 591560 151704 593000 151928 0 FreeSans 896 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 591560 184968 593000 185192 0 FreeSans 896 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 591560 218232 593000 218456 0 FreeSans 896 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 591560 262584 593000 262808 0 FreeSans 896 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 591560 306936 593000 307160 0 FreeSans 896 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 591560 351288 593000 351512 0 FreeSans 896 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 138488 -960 138712 480 0 FreeSans 896 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 474488 -960 474712 480 0 FreeSans 896 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 477848 -960 478072 480 0 FreeSans 896 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 481208 -960 481432 480 0 FreeSans 896 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 484568 -960 484792 480 0 FreeSans 896 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 487928 -960 488152 480 0 FreeSans 896 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 491288 -960 491512 480 0 FreeSans 896 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 494648 -960 494872 480 0 FreeSans 896 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 498008 -960 498232 480 0 FreeSans 896 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 501368 -960 501592 480 0 FreeSans 896 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 504728 -960 504952 480 0 FreeSans 896 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 172088 -960 172312 480 0 FreeSans 896 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 508088 -960 508312 480 0 FreeSans 896 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 511448 -960 511672 480 0 FreeSans 896 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 514808 -960 515032 480 0 FreeSans 896 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 518168 -960 518392 480 0 FreeSans 896 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 521528 -960 521752 480 0 FreeSans 896 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 524888 -960 525112 480 0 FreeSans 896 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 528248 -960 528472 480 0 FreeSans 896 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 531608 -960 531832 480 0 FreeSans 896 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 534968 -960 535192 480 0 FreeSans 896 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 538328 -960 538552 480 0 FreeSans 896 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 175448 -960 175672 480 0 FreeSans 896 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 541688 -960 541912 480 0 FreeSans 896 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 545048 -960 545272 480 0 FreeSans 896 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 548408 -960 548632 480 0 FreeSans 896 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 551768 -960 551992 480 0 FreeSans 896 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 555128 -960 555352 480 0 FreeSans 896 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 558488 -960 558712 480 0 FreeSans 896 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 561848 -960 562072 480 0 FreeSans 896 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 565208 -960 565432 480 0 FreeSans 896 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 178808 -960 179032 480 0 FreeSans 896 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 182168 -960 182392 480 0 FreeSans 896 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 185528 -960 185752 480 0 FreeSans 896 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 188888 -960 189112 480 0 FreeSans 896 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 192248 -960 192472 480 0 FreeSans 896 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 195608 -960 195832 480 0 FreeSans 896 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 198968 -960 199192 480 0 FreeSans 896 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 202328 -960 202552 480 0 FreeSans 896 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 141848 -960 142072 480 0 FreeSans 896 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 205688 -960 205912 480 0 FreeSans 896 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 209048 -960 209272 480 0 FreeSans 896 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 212408 -960 212632 480 0 FreeSans 896 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 215768 -960 215992 480 0 FreeSans 896 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 219128 -960 219352 480 0 FreeSans 896 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 222488 -960 222712 480 0 FreeSans 896 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 225848 -960 226072 480 0 FreeSans 896 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 229208 -960 229432 480 0 FreeSans 896 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 232568 -960 232792 480 0 FreeSans 896 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 235928 -960 236152 480 0 FreeSans 896 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 145208 -960 145432 480 0 FreeSans 896 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 239288 -960 239512 480 0 FreeSans 896 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 242648 -960 242872 480 0 FreeSans 896 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 246008 -960 246232 480 0 FreeSans 896 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 249368 -960 249592 480 0 FreeSans 896 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 252728 -960 252952 480 0 FreeSans 896 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 256088 -960 256312 480 0 FreeSans 896 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 259448 -960 259672 480 0 FreeSans 896 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 262808 -960 263032 480 0 FreeSans 896 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 266168 -960 266392 480 0 FreeSans 896 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 269528 -960 269752 480 0 FreeSans 896 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 148568 -960 148792 480 0 FreeSans 896 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 272888 -960 273112 480 0 FreeSans 896 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 276248 -960 276472 480 0 FreeSans 896 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 279608 -960 279832 480 0 FreeSans 896 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 282968 -960 283192 480 0 FreeSans 896 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 286328 -960 286552 480 0 FreeSans 896 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 289688 -960 289912 480 0 FreeSans 896 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 293048 -960 293272 480 0 FreeSans 896 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 296408 -960 296632 480 0 FreeSans 896 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 299768 -960 299992 480 0 FreeSans 896 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 303128 -960 303352 480 0 FreeSans 896 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 151928 -960 152152 480 0 FreeSans 896 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 306488 -960 306712 480 0 FreeSans 896 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 309848 -960 310072 480 0 FreeSans 896 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 313208 -960 313432 480 0 FreeSans 896 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 316568 -960 316792 480 0 FreeSans 896 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 319928 -960 320152 480 0 FreeSans 896 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 323288 -960 323512 480 0 FreeSans 896 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 326648 -960 326872 480 0 FreeSans 896 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 330008 -960 330232 480 0 FreeSans 896 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 333368 -960 333592 480 0 FreeSans 896 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 336728 -960 336952 480 0 FreeSans 896 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 155288 -960 155512 480 0 FreeSans 896 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 340088 -960 340312 480 0 FreeSans 896 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 343448 -960 343672 480 0 FreeSans 896 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 346808 -960 347032 480 0 FreeSans 896 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 350168 -960 350392 480 0 FreeSans 896 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 353528 -960 353752 480 0 FreeSans 896 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356888 -960 357112 480 0 FreeSans 896 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 360248 -960 360472 480 0 FreeSans 896 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363608 -960 363832 480 0 FreeSans 896 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366968 -960 367192 480 0 FreeSans 896 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370328 -960 370552 480 0 FreeSans 896 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 158648 -960 158872 480 0 FreeSans 896 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 373688 -960 373912 480 0 FreeSans 896 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377048 -960 377272 480 0 FreeSans 896 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 380408 -960 380632 480 0 FreeSans 896 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 383768 -960 383992 480 0 FreeSans 896 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 387128 -960 387352 480 0 FreeSans 896 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 390488 -960 390712 480 0 FreeSans 896 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 393848 -960 394072 480 0 FreeSans 896 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 397208 -960 397432 480 0 FreeSans 896 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 400568 -960 400792 480 0 FreeSans 896 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 403928 -960 404152 480 0 FreeSans 896 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 162008 -960 162232 480 0 FreeSans 896 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 407288 -960 407512 480 0 FreeSans 896 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 410648 -960 410872 480 0 FreeSans 896 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 414008 -960 414232 480 0 FreeSans 896 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 417368 -960 417592 480 0 FreeSans 896 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 420728 -960 420952 480 0 FreeSans 896 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 424088 -960 424312 480 0 FreeSans 896 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 427448 -960 427672 480 0 FreeSans 896 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 430808 -960 431032 480 0 FreeSans 896 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 434168 -960 434392 480 0 FreeSans 896 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 437528 -960 437752 480 0 FreeSans 896 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 165368 -960 165592 480 0 FreeSans 896 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 440888 -960 441112 480 0 FreeSans 896 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 444248 -960 444472 480 0 FreeSans 896 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 447608 -960 447832 480 0 FreeSans 896 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 450968 -960 451192 480 0 FreeSans 896 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 454328 -960 454552 480 0 FreeSans 896 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 457688 -960 457912 480 0 FreeSans 896 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 461048 -960 461272 480 0 FreeSans 896 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 464408 -960 464632 480 0 FreeSans 896 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 467768 -960 467992 480 0 FreeSans 896 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 471128 -960 471352 480 0 FreeSans 896 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 168728 -960 168952 480 0 FreeSans 896 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 139608 -960 139832 480 0 FreeSans 896 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 475608 -960 475832 480 0 FreeSans 896 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 478968 -960 479192 480 0 FreeSans 896 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 482328 -960 482552 480 0 FreeSans 896 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 485688 -960 485912 480 0 FreeSans 896 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 489048 -960 489272 480 0 FreeSans 896 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 492408 -960 492632 480 0 FreeSans 896 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 495768 -960 495992 480 0 FreeSans 896 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 499128 -960 499352 480 0 FreeSans 896 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 502488 -960 502712 480 0 FreeSans 896 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 505848 -960 506072 480 0 FreeSans 896 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 173208 -960 173432 480 0 FreeSans 896 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 509208 -960 509432 480 0 FreeSans 896 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 512568 -960 512792 480 0 FreeSans 896 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 515928 -960 516152 480 0 FreeSans 896 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 519288 -960 519512 480 0 FreeSans 896 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 522648 -960 522872 480 0 FreeSans 896 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 526008 -960 526232 480 0 FreeSans 896 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 529368 -960 529592 480 0 FreeSans 896 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 532728 -960 532952 480 0 FreeSans 896 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 536088 -960 536312 480 0 FreeSans 896 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 539448 -960 539672 480 0 FreeSans 896 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 176568 -960 176792 480 0 FreeSans 896 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 542808 -960 543032 480 0 FreeSans 896 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 546168 -960 546392 480 0 FreeSans 896 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 549528 -960 549752 480 0 FreeSans 896 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 552888 -960 553112 480 0 FreeSans 896 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 556248 -960 556472 480 0 FreeSans 896 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 559608 -960 559832 480 0 FreeSans 896 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 562968 -960 563192 480 0 FreeSans 896 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 566328 -960 566552 480 0 FreeSans 896 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 179928 -960 180152 480 0 FreeSans 896 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 183288 -960 183512 480 0 FreeSans 896 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 186648 -960 186872 480 0 FreeSans 896 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 190008 -960 190232 480 0 FreeSans 896 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 193368 -960 193592 480 0 FreeSans 896 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 196728 -960 196952 480 0 FreeSans 896 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 200088 -960 200312 480 0 FreeSans 896 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 203448 -960 203672 480 0 FreeSans 896 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 142968 -960 143192 480 0 FreeSans 896 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 206808 -960 207032 480 0 FreeSans 896 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 210168 -960 210392 480 0 FreeSans 896 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 213528 -960 213752 480 0 FreeSans 896 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 216888 -960 217112 480 0 FreeSans 896 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 220248 -960 220472 480 0 FreeSans 896 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 223608 -960 223832 480 0 FreeSans 896 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 226968 -960 227192 480 0 FreeSans 896 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 230328 -960 230552 480 0 FreeSans 896 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 233688 -960 233912 480 0 FreeSans 896 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 237048 -960 237272 480 0 FreeSans 896 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 146328 -960 146552 480 0 FreeSans 896 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 240408 -960 240632 480 0 FreeSans 896 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 243768 -960 243992 480 0 FreeSans 896 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 247128 -960 247352 480 0 FreeSans 896 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 250488 -960 250712 480 0 FreeSans 896 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 253848 -960 254072 480 0 FreeSans 896 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 257208 -960 257432 480 0 FreeSans 896 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 260568 -960 260792 480 0 FreeSans 896 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 263928 -960 264152 480 0 FreeSans 896 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 267288 -960 267512 480 0 FreeSans 896 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 270648 -960 270872 480 0 FreeSans 896 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 149688 -960 149912 480 0 FreeSans 896 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 274008 -960 274232 480 0 FreeSans 896 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 277368 -960 277592 480 0 FreeSans 896 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 280728 -960 280952 480 0 FreeSans 896 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 284088 -960 284312 480 0 FreeSans 896 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 287448 -960 287672 480 0 FreeSans 896 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 290808 -960 291032 480 0 FreeSans 896 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 294168 -960 294392 480 0 FreeSans 896 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 297528 -960 297752 480 0 FreeSans 896 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 300888 -960 301112 480 0 FreeSans 896 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 304248 -960 304472 480 0 FreeSans 896 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 153048 -960 153272 480 0 FreeSans 896 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 307608 -960 307832 480 0 FreeSans 896 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 310968 -960 311192 480 0 FreeSans 896 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 314328 -960 314552 480 0 FreeSans 896 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 317688 -960 317912 480 0 FreeSans 896 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 321048 -960 321272 480 0 FreeSans 896 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 324408 -960 324632 480 0 FreeSans 896 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 327768 -960 327992 480 0 FreeSans 896 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 331128 -960 331352 480 0 FreeSans 896 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 334488 -960 334712 480 0 FreeSans 896 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 337848 -960 338072 480 0 FreeSans 896 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 156408 -960 156632 480 0 FreeSans 896 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 341208 -960 341432 480 0 FreeSans 896 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 344568 -960 344792 480 0 FreeSans 896 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 347928 -960 348152 480 0 FreeSans 896 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 351288 -960 351512 480 0 FreeSans 896 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354648 -960 354872 480 0 FreeSans 896 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 358008 -960 358232 480 0 FreeSans 896 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361368 -960 361592 480 0 FreeSans 896 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364728 -960 364952 480 0 FreeSans 896 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368088 -960 368312 480 0 FreeSans 896 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371448 -960 371672 480 0 FreeSans 896 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 159768 -960 159992 480 0 FreeSans 896 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 374808 -960 375032 480 0 FreeSans 896 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378168 -960 378392 480 0 FreeSans 896 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 381528 -960 381752 480 0 FreeSans 896 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 384888 -960 385112 480 0 FreeSans 896 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 388248 -960 388472 480 0 FreeSans 896 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 391608 -960 391832 480 0 FreeSans 896 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 394968 -960 395192 480 0 FreeSans 896 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 398328 -960 398552 480 0 FreeSans 896 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 401688 -960 401912 480 0 FreeSans 896 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 405048 -960 405272 480 0 FreeSans 896 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 163128 -960 163352 480 0 FreeSans 896 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 408408 -960 408632 480 0 FreeSans 896 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 411768 -960 411992 480 0 FreeSans 896 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 415128 -960 415352 480 0 FreeSans 896 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 418488 -960 418712 480 0 FreeSans 896 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 421848 -960 422072 480 0 FreeSans 896 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 425208 -960 425432 480 0 FreeSans 896 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 428568 -960 428792 480 0 FreeSans 896 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 431928 -960 432152 480 0 FreeSans 896 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 435288 -960 435512 480 0 FreeSans 896 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 438648 -960 438872 480 0 FreeSans 896 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 166488 -960 166712 480 0 FreeSans 896 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 442008 -960 442232 480 0 FreeSans 896 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 445368 -960 445592 480 0 FreeSans 896 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 448728 -960 448952 480 0 FreeSans 896 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 452088 -960 452312 480 0 FreeSans 896 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 455448 -960 455672 480 0 FreeSans 896 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 458808 -960 459032 480 0 FreeSans 896 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 462168 -960 462392 480 0 FreeSans 896 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 465528 -960 465752 480 0 FreeSans 896 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 468888 -960 469112 480 0 FreeSans 896 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 472248 -960 472472 480 0 FreeSans 896 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 169848 -960 170072 480 0 FreeSans 896 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 140728 -960 140952 480 0 FreeSans 896 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 476728 -960 476952 480 0 FreeSans 896 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 480088 -960 480312 480 0 FreeSans 896 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 483448 -960 483672 480 0 FreeSans 896 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 486808 -960 487032 480 0 FreeSans 896 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 490168 -960 490392 480 0 FreeSans 896 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 493528 -960 493752 480 0 FreeSans 896 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 496888 -960 497112 480 0 FreeSans 896 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 500248 -960 500472 480 0 FreeSans 896 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 503608 -960 503832 480 0 FreeSans 896 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 506968 -960 507192 480 0 FreeSans 896 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 174328 -960 174552 480 0 FreeSans 896 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 510328 -960 510552 480 0 FreeSans 896 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 513688 -960 513912 480 0 FreeSans 896 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 517048 -960 517272 480 0 FreeSans 896 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 520408 -960 520632 480 0 FreeSans 896 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 523768 -960 523992 480 0 FreeSans 896 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 527128 -960 527352 480 0 FreeSans 896 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 530488 -960 530712 480 0 FreeSans 896 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 533848 -960 534072 480 0 FreeSans 896 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 537208 -960 537432 480 0 FreeSans 896 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 540568 -960 540792 480 0 FreeSans 896 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 177688 -960 177912 480 0 FreeSans 896 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 543928 -960 544152 480 0 FreeSans 896 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 547288 -960 547512 480 0 FreeSans 896 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 550648 -960 550872 480 0 FreeSans 896 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 554008 -960 554232 480 0 FreeSans 896 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 557368 -960 557592 480 0 FreeSans 896 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 560728 -960 560952 480 0 FreeSans 896 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 564088 -960 564312 480 0 FreeSans 896 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 567448 -960 567672 480 0 FreeSans 896 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 181048 -960 181272 480 0 FreeSans 896 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 184408 -960 184632 480 0 FreeSans 896 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 187768 -960 187992 480 0 FreeSans 896 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 191128 -960 191352 480 0 FreeSans 896 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 194488 -960 194712 480 0 FreeSans 896 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 197848 -960 198072 480 0 FreeSans 896 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 201208 -960 201432 480 0 FreeSans 896 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 204568 -960 204792 480 0 FreeSans 896 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 144088 -960 144312 480 0 FreeSans 896 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 207928 -960 208152 480 0 FreeSans 896 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 211288 -960 211512 480 0 FreeSans 896 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 214648 -960 214872 480 0 FreeSans 896 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 218008 -960 218232 480 0 FreeSans 896 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 221368 -960 221592 480 0 FreeSans 896 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 224728 -960 224952 480 0 FreeSans 896 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 228088 -960 228312 480 0 FreeSans 896 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 231448 -960 231672 480 0 FreeSans 896 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 234808 -960 235032 480 0 FreeSans 896 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 238168 -960 238392 480 0 FreeSans 896 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 147448 -960 147672 480 0 FreeSans 896 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 241528 -960 241752 480 0 FreeSans 896 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 244888 -960 245112 480 0 FreeSans 896 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 248248 -960 248472 480 0 FreeSans 896 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 251608 -960 251832 480 0 FreeSans 896 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 254968 -960 255192 480 0 FreeSans 896 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 258328 -960 258552 480 0 FreeSans 896 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 261688 -960 261912 480 0 FreeSans 896 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 265048 -960 265272 480 0 FreeSans 896 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 268408 -960 268632 480 0 FreeSans 896 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 271768 -960 271992 480 0 FreeSans 896 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 150808 -960 151032 480 0 FreeSans 896 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 275128 -960 275352 480 0 FreeSans 896 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 278488 -960 278712 480 0 FreeSans 896 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 281848 -960 282072 480 0 FreeSans 896 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 285208 -960 285432 480 0 FreeSans 896 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 288568 -960 288792 480 0 FreeSans 896 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 291928 -960 292152 480 0 FreeSans 896 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 295288 -960 295512 480 0 FreeSans 896 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 298648 -960 298872 480 0 FreeSans 896 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 302008 -960 302232 480 0 FreeSans 896 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 305368 -960 305592 480 0 FreeSans 896 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 154168 -960 154392 480 0 FreeSans 896 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 308728 -960 308952 480 0 FreeSans 896 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 312088 -960 312312 480 0 FreeSans 896 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 315448 -960 315672 480 0 FreeSans 896 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 318808 -960 319032 480 0 FreeSans 896 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 322168 -960 322392 480 0 FreeSans 896 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 325528 -960 325752 480 0 FreeSans 896 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 328888 -960 329112 480 0 FreeSans 896 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 332248 -960 332472 480 0 FreeSans 896 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 335608 -960 335832 480 0 FreeSans 896 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 338968 -960 339192 480 0 FreeSans 896 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 157528 -960 157752 480 0 FreeSans 896 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 342328 -960 342552 480 0 FreeSans 896 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 345688 -960 345912 480 0 FreeSans 896 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 349048 -960 349272 480 0 FreeSans 896 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 352408 -960 352632 480 0 FreeSans 896 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355768 -960 355992 480 0 FreeSans 896 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 359128 -960 359352 480 0 FreeSans 896 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362488 -960 362712 480 0 FreeSans 896 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365848 -960 366072 480 0 FreeSans 896 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369208 -960 369432 480 0 FreeSans 896 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372568 -960 372792 480 0 FreeSans 896 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 160888 -960 161112 480 0 FreeSans 896 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 375928 -960 376152 480 0 FreeSans 896 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379288 -960 379512 480 0 FreeSans 896 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 382648 -960 382872 480 0 FreeSans 896 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 386008 -960 386232 480 0 FreeSans 896 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 389368 -960 389592 480 0 FreeSans 896 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 392728 -960 392952 480 0 FreeSans 896 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 396088 -960 396312 480 0 FreeSans 896 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 399448 -960 399672 480 0 FreeSans 896 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 402808 -960 403032 480 0 FreeSans 896 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 406168 -960 406392 480 0 FreeSans 896 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 164248 -960 164472 480 0 FreeSans 896 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 409528 -960 409752 480 0 FreeSans 896 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 412888 -960 413112 480 0 FreeSans 896 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 416248 -960 416472 480 0 FreeSans 896 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 419608 -960 419832 480 0 FreeSans 896 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 422968 -960 423192 480 0 FreeSans 896 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 426328 -960 426552 480 0 FreeSans 896 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 429688 -960 429912 480 0 FreeSans 896 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 433048 -960 433272 480 0 FreeSans 896 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 436408 -960 436632 480 0 FreeSans 896 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 439768 -960 439992 480 0 FreeSans 896 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 167608 -960 167832 480 0 FreeSans 896 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 443128 -960 443352 480 0 FreeSans 896 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 446488 -960 446712 480 0 FreeSans 896 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 449848 -960 450072 480 0 FreeSans 896 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 453208 -960 453432 480 0 FreeSans 896 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 456568 -960 456792 480 0 FreeSans 896 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 459928 -960 460152 480 0 FreeSans 896 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 463288 -960 463512 480 0 FreeSans 896 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 466648 -960 466872 480 0 FreeSans 896 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 470008 -960 470232 480 0 FreeSans 896 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 473368 -960 473592 480 0 FreeSans 896 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 170968 -960 171192 480 0 FreeSans 896 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 568568 -960 568792 480 0 FreeSans 896 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 569688 -960 569912 480 0 FreeSans 896 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 570808 -960 571032 480 0 FreeSans 896 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 571928 -960 572152 480 0 FreeSans 896 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -956 -684 -336 597308 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal5 s -956 -684 597020 -64 0 FreeSans 4608 0 0 0 vdd
port 531 nsew power bidirectional
flabel metal5 s -956 596688 597020 597308 0 FreeSans 4608 0 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 596400 -684 597020 597308 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 3154 -1644 3774 598268 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 21154 -1644 21774 158858 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 21154 458342 21774 598268 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 39154 -1644 39774 158858 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 39154 458342 39774 598268 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 57154 -1644 57774 77594 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 57154 111238 57774 158858 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 57154 458342 57774 598268 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 75154 -1644 75774 77594 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 75154 111238 75774 158858 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 75154 458342 75774 598268 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 93154 -1644 93774 77594 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 93154 111238 93774 158858 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 93154 458342 93774 598268 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 111154 -1644 111774 77594 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 111154 111238 111774 158858 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 111154 458342 111774 598268 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 129154 -1644 129774 77594 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 129154 111238 129774 158858 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 129154 458342 129774 598268 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 147154 -1644 147774 77594 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 147154 111238 147774 158858 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 147154 458342 147774 598268 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 165154 -1644 165774 77594 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 165154 111238 165774 158858 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 165154 458342 165774 598268 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 183154 -1644 183774 158858 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 183154 458342 183774 598268 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 201154 -1644 201774 598268 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 219154 -1644 219774 8858 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 219154 148342 219774 158858 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 219154 458342 219774 598268 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 237154 -1644 237774 8858 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 237154 148342 237774 158858 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 237154 458342 237774 598268 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 255154 -1644 255774 8858 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 255154 148342 255774 158858 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 255154 458342 255774 598268 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 273154 -1644 273774 8858 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 273154 148342 273774 158858 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 273154 458342 273774 598268 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 291154 -1644 291774 8858 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 291154 148342 291774 158858 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 291154 458342 291774 598268 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 309154 -1644 309774 8858 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 309154 148342 309774 158858 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 309154 458342 309774 598268 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 327154 -1644 327774 8858 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 327154 148342 327774 158858 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 327154 458342 327774 598268 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 345154 -1644 345774 8858 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 345154 148342 345774 158858 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 345154 458342 345774 598268 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 363154 -1644 363774 8858 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 363154 148342 363774 158858 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 363154 458342 363774 598268 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 381154 -1644 381774 598268 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 399154 -1644 399774 598268 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 417154 -1644 417774 158858 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 417154 458342 417774 598268 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 435154 -1644 435774 158858 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 435154 458342 435774 598268 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 453154 -1644 453774 158858 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 453154 458342 453774 598268 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 471154 -1644 471774 158858 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 471154 458342 471774 598268 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 489154 -1644 489774 158858 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 489154 458342 489774 598268 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 507154 -1644 507774 158858 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 507154 458342 507774 598268 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 525154 -1644 525774 158858 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 525154 458342 525774 598268 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 543154 -1644 543774 158858 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 543154 458342 543774 598268 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 561154 -1644 561774 158858 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 561154 458342 561774 598268 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s 579154 -1644 579774 598268 0 FreeSans 2560 90 0 0 vdd
port 531 nsew power bidirectional
flabel metal5 s -1916 3826 597980 4446 0 FreeSans 4608 0 0 0 vdd
port 531 nsew power bidirectional
flabel metal5 s -1916 21826 597980 22446 0 FreeSans 4608 0 0 0 vdd
port 531 nsew power bidirectional
flabel metal5 s -1916 39826 597980 40446 0 FreeSans 4608 0 0 0 vdd
port 531 nsew power bidirectional
flabel metal5 s -1916 57826 597980 58446 0 FreeSans 4608 0 0 0 vdd
port 531 nsew power bidirectional
flabel metal5 s -1916 75826 597980 76446 0 FreeSans 4608 0 0 0 vdd
port 531 nsew power bidirectional
flabel metal5 s -1916 93826 597980 94446 0 FreeSans 4608 0 0 0 vdd
port 531 nsew power bidirectional
flabel metal5 s -1916 111826 597980 112446 0 FreeSans 4608 0 0 0 vdd
port 531 nsew power bidirectional
flabel metal5 s -1916 129826 597980 130446 0 FreeSans 4608 0 0 0 vdd
port 531 nsew power bidirectional
flabel metal5 s -1916 147826 597980 148446 0 FreeSans 4608 0 0 0 vdd
port 531 nsew power bidirectional
flabel metal5 s -1916 165826 597980 166446 0 FreeSans 4608 0 0 0 vdd
port 531 nsew power bidirectional
flabel metal5 s -1916 183826 597980 184446 0 FreeSans 4608 0 0 0 vdd
port 531 nsew power bidirectional
flabel metal5 s -1916 201826 597980 202446 0 FreeSans 4608 0 0 0 vdd
port 531 nsew power bidirectional
flabel metal5 s -1916 219826 597980 220446 0 FreeSans 4608 0 0 0 vdd
port 531 nsew power bidirectional
flabel metal5 s -1916 237826 597980 238446 0 FreeSans 4608 0 0 0 vdd
port 531 nsew power bidirectional
flabel metal5 s -1916 255826 597980 256446 0 FreeSans 4608 0 0 0 vdd
port 531 nsew power bidirectional
flabel metal5 s -1916 273826 597980 274446 0 FreeSans 4608 0 0 0 vdd
port 531 nsew power bidirectional
flabel metal5 s -1916 291826 597980 292446 0 FreeSans 4608 0 0 0 vdd
port 531 nsew power bidirectional
flabel metal5 s -1916 309826 597980 310446 0 FreeSans 4608 0 0 0 vdd
port 531 nsew power bidirectional
flabel metal5 s -1916 327826 597980 328446 0 FreeSans 4608 0 0 0 vdd
port 531 nsew power bidirectional
flabel metal5 s -1916 345826 597980 346446 0 FreeSans 4608 0 0 0 vdd
port 531 nsew power bidirectional
flabel metal5 s -1916 363826 597980 364446 0 FreeSans 4608 0 0 0 vdd
port 531 nsew power bidirectional
flabel metal5 s -1916 381826 597980 382446 0 FreeSans 4608 0 0 0 vdd
port 531 nsew power bidirectional
flabel metal5 s -1916 399826 597980 400446 0 FreeSans 4608 0 0 0 vdd
port 531 nsew power bidirectional
flabel metal5 s -1916 417826 597980 418446 0 FreeSans 4608 0 0 0 vdd
port 531 nsew power bidirectional
flabel metal5 s -1916 435826 597980 436446 0 FreeSans 4608 0 0 0 vdd
port 531 nsew power bidirectional
flabel metal5 s -1916 453826 597980 454446 0 FreeSans 4608 0 0 0 vdd
port 531 nsew power bidirectional
flabel metal5 s -1916 471826 597980 472446 0 FreeSans 4608 0 0 0 vdd
port 531 nsew power bidirectional
flabel metal5 s -1916 489826 597980 490446 0 FreeSans 4608 0 0 0 vdd
port 531 nsew power bidirectional
flabel metal5 s -1916 507826 597980 508446 0 FreeSans 4608 0 0 0 vdd
port 531 nsew power bidirectional
flabel metal5 s -1916 525826 597980 526446 0 FreeSans 4608 0 0 0 vdd
port 531 nsew power bidirectional
flabel metal5 s -1916 543826 597980 544446 0 FreeSans 4608 0 0 0 vdd
port 531 nsew power bidirectional
flabel metal5 s -1916 561826 597980 562446 0 FreeSans 4608 0 0 0 vdd
port 531 nsew power bidirectional
flabel metal5 s -1916 579826 597980 580446 0 FreeSans 4608 0 0 0 vdd
port 531 nsew power bidirectional
flabel metal4 s -1916 -1644 -1296 598268 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal5 s -1916 -1644 597980 -1024 0 FreeSans 4608 0 0 0 vss
port 532 nsew ground bidirectional
flabel metal5 s -1916 597648 597980 598268 0 FreeSans 4608 0 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 597360 -1644 597980 598268 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 6874 -1644 7494 598268 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 24874 -1644 25494 158858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 24874 298342 25494 318858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 24874 458342 25494 598268 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 42874 -1644 43494 158858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 42874 298342 43494 318858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 42874 458342 43494 598268 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 60874 -1644 61494 77594 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 60874 111238 61494 158858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 60874 298342 61494 318858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 60874 458342 61494 598268 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 78874 -1644 79494 77594 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 78874 111238 79494 158858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 78874 298342 79494 318858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 78874 458342 79494 598268 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 96874 -1644 97494 77594 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 96874 111238 97494 158858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 96874 298342 97494 318858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 96874 458342 97494 598268 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 114874 -1644 115494 77594 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 114874 111238 115494 158858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 114874 298342 115494 318858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 114874 458342 115494 598268 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 132874 -1644 133494 77594 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 132874 111238 133494 158858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 132874 298342 133494 318858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 132874 458342 133494 598268 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 150874 -1644 151494 77594 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 150874 111238 151494 158858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 150874 298342 151494 318858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 150874 458342 151494 598268 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 168874 -1644 169494 77594 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 168874 111238 169494 158858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 168874 298342 169494 318858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 168874 458342 169494 598268 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 186874 -1644 187494 158858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 186874 298342 187494 318858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 186874 458342 187494 598268 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 204874 -1644 205494 598268 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 222874 148342 223494 158858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 222874 298342 223494 318858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 222874 458342 223494 598268 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 240874 148342 241494 158858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 240874 298342 241494 318858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 240874 458342 241494 598268 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 258874 148342 259494 158858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 258874 298342 259494 318858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 258874 458342 259494 598268 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 276874 148342 277494 158858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 276874 298342 277494 318858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 276874 458342 277494 598268 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 294874 148342 295494 158858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 294874 298342 295494 318858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 294874 458342 295494 598268 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 312874 148342 313494 158858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 312874 298342 313494 318858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 312874 458342 313494 598268 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 330874 148342 331494 158858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 330874 298342 331494 318858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 330874 458342 331494 598268 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 348874 148342 349494 158858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 348874 298342 349494 318858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 348874 458342 349494 598268 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 366874 148342 367494 158858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 366874 298342 367494 318858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 366874 458342 367494 598268 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 384874 -1644 385494 598268 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 402874 -1644 403494 598268 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 420874 -1644 421494 158858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 420874 298342 421494 318858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 420874 458342 421494 598268 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 438874 -1644 439494 158858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 438874 298342 439494 318858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 438874 458342 439494 598268 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 456874 -1644 457494 158858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 456874 298342 457494 318858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 456874 458342 457494 598268 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 474874 -1644 475494 158858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 474874 298342 475494 318858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 474874 458342 475494 598268 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 492874 -1644 493494 158858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 492874 298342 493494 318858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 492874 458342 493494 598268 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 510874 -1644 511494 158858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 510874 298342 511494 318858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 510874 458342 511494 598268 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 528874 -1644 529494 158858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 528874 298342 529494 318858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 528874 458342 529494 598268 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 546874 -1644 547494 158858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 546874 298342 547494 318858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 546874 458342 547494 598268 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 564874 -1644 565494 158858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 564874 298342 565494 318858 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 564874 458342 565494 598268 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal4 s 582874 -1644 583494 598268 0 FreeSans 2560 90 0 0 vss
port 532 nsew ground bidirectional
flabel metal5 s -1916 9826 597980 10446 0 FreeSans 4608 0 0 0 vss
port 532 nsew ground bidirectional
flabel metal5 s -1916 27826 597980 28446 0 FreeSans 4608 0 0 0 vss
port 532 nsew ground bidirectional
flabel metal5 s -1916 45826 597980 46446 0 FreeSans 4608 0 0 0 vss
port 532 nsew ground bidirectional
flabel metal5 s -1916 63826 597980 64446 0 FreeSans 4608 0 0 0 vss
port 532 nsew ground bidirectional
flabel metal5 s -1916 81826 597980 82446 0 FreeSans 4608 0 0 0 vss
port 532 nsew ground bidirectional
flabel metal5 s -1916 99826 597980 100446 0 FreeSans 4608 0 0 0 vss
port 532 nsew ground bidirectional
flabel metal5 s -1916 117826 597980 118446 0 FreeSans 4608 0 0 0 vss
port 532 nsew ground bidirectional
flabel metal5 s -1916 135826 597980 136446 0 FreeSans 4608 0 0 0 vss
port 532 nsew ground bidirectional
flabel metal5 s -1916 153826 597980 154446 0 FreeSans 4608 0 0 0 vss
port 532 nsew ground bidirectional
flabel metal5 s -1916 171826 597980 172446 0 FreeSans 4608 0 0 0 vss
port 532 nsew ground bidirectional
flabel metal5 s -1916 189826 597980 190446 0 FreeSans 4608 0 0 0 vss
port 532 nsew ground bidirectional
flabel metal5 s -1916 207826 597980 208446 0 FreeSans 4608 0 0 0 vss
port 532 nsew ground bidirectional
flabel metal5 s -1916 225826 597980 226446 0 FreeSans 4608 0 0 0 vss
port 532 nsew ground bidirectional
flabel metal5 s -1916 243826 597980 244446 0 FreeSans 4608 0 0 0 vss
port 532 nsew ground bidirectional
flabel metal5 s -1916 261826 597980 262446 0 FreeSans 4608 0 0 0 vss
port 532 nsew ground bidirectional
flabel metal5 s -1916 279826 597980 280446 0 FreeSans 4608 0 0 0 vss
port 532 nsew ground bidirectional
flabel metal5 s -1916 297826 597980 298446 0 FreeSans 4608 0 0 0 vss
port 532 nsew ground bidirectional
flabel metal5 s -1916 315826 597980 316446 0 FreeSans 4608 0 0 0 vss
port 532 nsew ground bidirectional
flabel metal5 s -1916 333826 597980 334446 0 FreeSans 4608 0 0 0 vss
port 532 nsew ground bidirectional
flabel metal5 s -1916 351826 597980 352446 0 FreeSans 4608 0 0 0 vss
port 532 nsew ground bidirectional
flabel metal5 s -1916 369826 597980 370446 0 FreeSans 4608 0 0 0 vss
port 532 nsew ground bidirectional
flabel metal5 s -1916 387826 597980 388446 0 FreeSans 4608 0 0 0 vss
port 532 nsew ground bidirectional
flabel metal5 s -1916 405826 597980 406446 0 FreeSans 4608 0 0 0 vss
port 532 nsew ground bidirectional
flabel metal5 s -1916 423826 597980 424446 0 FreeSans 4608 0 0 0 vss
port 532 nsew ground bidirectional
flabel metal5 s -1916 441826 597980 442446 0 FreeSans 4608 0 0 0 vss
port 532 nsew ground bidirectional
flabel metal5 s -1916 459826 597980 460446 0 FreeSans 4608 0 0 0 vss
port 532 nsew ground bidirectional
flabel metal5 s -1916 477826 597980 478446 0 FreeSans 4608 0 0 0 vss
port 532 nsew ground bidirectional
flabel metal5 s -1916 495826 597980 496446 0 FreeSans 4608 0 0 0 vss
port 532 nsew ground bidirectional
flabel metal5 s -1916 513826 597980 514446 0 FreeSans 4608 0 0 0 vss
port 532 nsew ground bidirectional
flabel metal5 s -1916 531826 597980 532446 0 FreeSans 4608 0 0 0 vss
port 532 nsew ground bidirectional
flabel metal5 s -1916 549826 597980 550446 0 FreeSans 4608 0 0 0 vss
port 532 nsew ground bidirectional
flabel metal5 s -1916 567826 597980 568446 0 FreeSans 4608 0 0 0 vss
port 532 nsew ground bidirectional
flabel metal5 s -1916 585826 597980 586446 0 FreeSans 4608 0 0 0 vss
port 532 nsew ground bidirectional
flabel metal2 s 19768 -960 19992 480 0 FreeSans 896 90 0 0 wb_clk_i
port 533 nsew signal input
flabel metal2 s 20888 -960 21112 480 0 FreeSans 896 90 0 0 wb_rst_i
port 534 nsew signal input
flabel metal2 s 22008 -960 22232 480 0 FreeSans 896 90 0 0 wbs_ack_o
port 535 nsew signal tristate
flabel metal2 s 26488 -960 26712 480 0 FreeSans 896 90 0 0 wbs_adr_i[0]
port 536 nsew signal input
flabel metal2 s 64568 -960 64792 480 0 FreeSans 896 90 0 0 wbs_adr_i[10]
port 537 nsew signal input
flabel metal2 s 67928 -960 68152 480 0 FreeSans 896 90 0 0 wbs_adr_i[11]
port 538 nsew signal input
flabel metal2 s 71288 -960 71512 480 0 FreeSans 896 90 0 0 wbs_adr_i[12]
port 539 nsew signal input
flabel metal2 s 74648 -960 74872 480 0 FreeSans 896 90 0 0 wbs_adr_i[13]
port 540 nsew signal input
flabel metal2 s 78008 -960 78232 480 0 FreeSans 896 90 0 0 wbs_adr_i[14]
port 541 nsew signal input
flabel metal2 s 81368 -960 81592 480 0 FreeSans 896 90 0 0 wbs_adr_i[15]
port 542 nsew signal input
flabel metal2 s 84728 -960 84952 480 0 FreeSans 896 90 0 0 wbs_adr_i[16]
port 543 nsew signal input
flabel metal2 s 88088 -960 88312 480 0 FreeSans 896 90 0 0 wbs_adr_i[17]
port 544 nsew signal input
flabel metal2 s 91448 -960 91672 480 0 FreeSans 896 90 0 0 wbs_adr_i[18]
port 545 nsew signal input
flabel metal2 s 94808 -960 95032 480 0 FreeSans 896 90 0 0 wbs_adr_i[19]
port 546 nsew signal input
flabel metal2 s 30968 -960 31192 480 0 FreeSans 896 90 0 0 wbs_adr_i[1]
port 547 nsew signal input
flabel metal2 s 98168 -960 98392 480 0 FreeSans 896 90 0 0 wbs_adr_i[20]
port 548 nsew signal input
flabel metal2 s 101528 -960 101752 480 0 FreeSans 896 90 0 0 wbs_adr_i[21]
port 549 nsew signal input
flabel metal2 s 104888 -960 105112 480 0 FreeSans 896 90 0 0 wbs_adr_i[22]
port 550 nsew signal input
flabel metal2 s 108248 -960 108472 480 0 FreeSans 896 90 0 0 wbs_adr_i[23]
port 551 nsew signal input
flabel metal2 s 111608 -960 111832 480 0 FreeSans 896 90 0 0 wbs_adr_i[24]
port 552 nsew signal input
flabel metal2 s 114968 -960 115192 480 0 FreeSans 896 90 0 0 wbs_adr_i[25]
port 553 nsew signal input
flabel metal2 s 118328 -960 118552 480 0 FreeSans 896 90 0 0 wbs_adr_i[26]
port 554 nsew signal input
flabel metal2 s 121688 -960 121912 480 0 FreeSans 896 90 0 0 wbs_adr_i[27]
port 555 nsew signal input
flabel metal2 s 125048 -960 125272 480 0 FreeSans 896 90 0 0 wbs_adr_i[28]
port 556 nsew signal input
flabel metal2 s 128408 -960 128632 480 0 FreeSans 896 90 0 0 wbs_adr_i[29]
port 557 nsew signal input
flabel metal2 s 35448 -960 35672 480 0 FreeSans 896 90 0 0 wbs_adr_i[2]
port 558 nsew signal input
flabel metal2 s 131768 -960 131992 480 0 FreeSans 896 90 0 0 wbs_adr_i[30]
port 559 nsew signal input
flabel metal2 s 135128 -960 135352 480 0 FreeSans 896 90 0 0 wbs_adr_i[31]
port 560 nsew signal input
flabel metal2 s 39928 -960 40152 480 0 FreeSans 896 90 0 0 wbs_adr_i[3]
port 561 nsew signal input
flabel metal2 s 44408 -960 44632 480 0 FreeSans 896 90 0 0 wbs_adr_i[4]
port 562 nsew signal input
flabel metal2 s 47768 -960 47992 480 0 FreeSans 896 90 0 0 wbs_adr_i[5]
port 563 nsew signal input
flabel metal2 s 51128 -960 51352 480 0 FreeSans 896 90 0 0 wbs_adr_i[6]
port 564 nsew signal input
flabel metal2 s 54488 -960 54712 480 0 FreeSans 896 90 0 0 wbs_adr_i[7]
port 565 nsew signal input
flabel metal2 s 57848 -960 58072 480 0 FreeSans 896 90 0 0 wbs_adr_i[8]
port 566 nsew signal input
flabel metal2 s 61208 -960 61432 480 0 FreeSans 896 90 0 0 wbs_adr_i[9]
port 567 nsew signal input
flabel metal2 s 23128 -960 23352 480 0 FreeSans 896 90 0 0 wbs_cyc_i
port 568 nsew signal input
flabel metal2 s 27608 -960 27832 480 0 FreeSans 896 90 0 0 wbs_dat_i[0]
port 569 nsew signal input
flabel metal2 s 65688 -960 65912 480 0 FreeSans 896 90 0 0 wbs_dat_i[10]
port 570 nsew signal input
flabel metal2 s 69048 -960 69272 480 0 FreeSans 896 90 0 0 wbs_dat_i[11]
port 571 nsew signal input
flabel metal2 s 72408 -960 72632 480 0 FreeSans 896 90 0 0 wbs_dat_i[12]
port 572 nsew signal input
flabel metal2 s 75768 -960 75992 480 0 FreeSans 896 90 0 0 wbs_dat_i[13]
port 573 nsew signal input
flabel metal2 s 79128 -960 79352 480 0 FreeSans 896 90 0 0 wbs_dat_i[14]
port 574 nsew signal input
flabel metal2 s 82488 -960 82712 480 0 FreeSans 896 90 0 0 wbs_dat_i[15]
port 575 nsew signal input
flabel metal2 s 85848 -960 86072 480 0 FreeSans 896 90 0 0 wbs_dat_i[16]
port 576 nsew signal input
flabel metal2 s 89208 -960 89432 480 0 FreeSans 896 90 0 0 wbs_dat_i[17]
port 577 nsew signal input
flabel metal2 s 92568 -960 92792 480 0 FreeSans 896 90 0 0 wbs_dat_i[18]
port 578 nsew signal input
flabel metal2 s 95928 -960 96152 480 0 FreeSans 896 90 0 0 wbs_dat_i[19]
port 579 nsew signal input
flabel metal2 s 32088 -960 32312 480 0 FreeSans 896 90 0 0 wbs_dat_i[1]
port 580 nsew signal input
flabel metal2 s 99288 -960 99512 480 0 FreeSans 896 90 0 0 wbs_dat_i[20]
port 581 nsew signal input
flabel metal2 s 102648 -960 102872 480 0 FreeSans 896 90 0 0 wbs_dat_i[21]
port 582 nsew signal input
flabel metal2 s 106008 -960 106232 480 0 FreeSans 896 90 0 0 wbs_dat_i[22]
port 583 nsew signal input
flabel metal2 s 109368 -960 109592 480 0 FreeSans 896 90 0 0 wbs_dat_i[23]
port 584 nsew signal input
flabel metal2 s 112728 -960 112952 480 0 FreeSans 896 90 0 0 wbs_dat_i[24]
port 585 nsew signal input
flabel metal2 s 116088 -960 116312 480 0 FreeSans 896 90 0 0 wbs_dat_i[25]
port 586 nsew signal input
flabel metal2 s 119448 -960 119672 480 0 FreeSans 896 90 0 0 wbs_dat_i[26]
port 587 nsew signal input
flabel metal2 s 122808 -960 123032 480 0 FreeSans 896 90 0 0 wbs_dat_i[27]
port 588 nsew signal input
flabel metal2 s 126168 -960 126392 480 0 FreeSans 896 90 0 0 wbs_dat_i[28]
port 589 nsew signal input
flabel metal2 s 129528 -960 129752 480 0 FreeSans 896 90 0 0 wbs_dat_i[29]
port 590 nsew signal input
flabel metal2 s 36568 -960 36792 480 0 FreeSans 896 90 0 0 wbs_dat_i[2]
port 591 nsew signal input
flabel metal2 s 132888 -960 133112 480 0 FreeSans 896 90 0 0 wbs_dat_i[30]
port 592 nsew signal input
flabel metal2 s 136248 -960 136472 480 0 FreeSans 896 90 0 0 wbs_dat_i[31]
port 593 nsew signal input
flabel metal2 s 41048 -960 41272 480 0 FreeSans 896 90 0 0 wbs_dat_i[3]
port 594 nsew signal input
flabel metal2 s 45528 -960 45752 480 0 FreeSans 896 90 0 0 wbs_dat_i[4]
port 595 nsew signal input
flabel metal2 s 48888 -960 49112 480 0 FreeSans 896 90 0 0 wbs_dat_i[5]
port 596 nsew signal input
flabel metal2 s 52248 -960 52472 480 0 FreeSans 896 90 0 0 wbs_dat_i[6]
port 597 nsew signal input
flabel metal2 s 55608 -960 55832 480 0 FreeSans 896 90 0 0 wbs_dat_i[7]
port 598 nsew signal input
flabel metal2 s 58968 -960 59192 480 0 FreeSans 896 90 0 0 wbs_dat_i[8]
port 599 nsew signal input
flabel metal2 s 62328 -960 62552 480 0 FreeSans 896 90 0 0 wbs_dat_i[9]
port 600 nsew signal input
flabel metal2 s 28728 -960 28952 480 0 FreeSans 896 90 0 0 wbs_dat_o[0]
port 601 nsew signal tristate
flabel metal2 s 66808 -960 67032 480 0 FreeSans 896 90 0 0 wbs_dat_o[10]
port 602 nsew signal tristate
flabel metal2 s 70168 -960 70392 480 0 FreeSans 896 90 0 0 wbs_dat_o[11]
port 603 nsew signal tristate
flabel metal2 s 73528 -960 73752 480 0 FreeSans 896 90 0 0 wbs_dat_o[12]
port 604 nsew signal tristate
flabel metal2 s 76888 -960 77112 480 0 FreeSans 896 90 0 0 wbs_dat_o[13]
port 605 nsew signal tristate
flabel metal2 s 80248 -960 80472 480 0 FreeSans 896 90 0 0 wbs_dat_o[14]
port 606 nsew signal tristate
flabel metal2 s 83608 -960 83832 480 0 FreeSans 896 90 0 0 wbs_dat_o[15]
port 607 nsew signal tristate
flabel metal2 s 86968 -960 87192 480 0 FreeSans 896 90 0 0 wbs_dat_o[16]
port 608 nsew signal tristate
flabel metal2 s 90328 -960 90552 480 0 FreeSans 896 90 0 0 wbs_dat_o[17]
port 609 nsew signal tristate
flabel metal2 s 93688 -960 93912 480 0 FreeSans 896 90 0 0 wbs_dat_o[18]
port 610 nsew signal tristate
flabel metal2 s 97048 -960 97272 480 0 FreeSans 896 90 0 0 wbs_dat_o[19]
port 611 nsew signal tristate
flabel metal2 s 33208 -960 33432 480 0 FreeSans 896 90 0 0 wbs_dat_o[1]
port 612 nsew signal tristate
flabel metal2 s 100408 -960 100632 480 0 FreeSans 896 90 0 0 wbs_dat_o[20]
port 613 nsew signal tristate
flabel metal2 s 103768 -960 103992 480 0 FreeSans 896 90 0 0 wbs_dat_o[21]
port 614 nsew signal tristate
flabel metal2 s 107128 -960 107352 480 0 FreeSans 896 90 0 0 wbs_dat_o[22]
port 615 nsew signal tristate
flabel metal2 s 110488 -960 110712 480 0 FreeSans 896 90 0 0 wbs_dat_o[23]
port 616 nsew signal tristate
flabel metal2 s 113848 -960 114072 480 0 FreeSans 896 90 0 0 wbs_dat_o[24]
port 617 nsew signal tristate
flabel metal2 s 117208 -960 117432 480 0 FreeSans 896 90 0 0 wbs_dat_o[25]
port 618 nsew signal tristate
flabel metal2 s 120568 -960 120792 480 0 FreeSans 896 90 0 0 wbs_dat_o[26]
port 619 nsew signal tristate
flabel metal2 s 123928 -960 124152 480 0 FreeSans 896 90 0 0 wbs_dat_o[27]
port 620 nsew signal tristate
flabel metal2 s 127288 -960 127512 480 0 FreeSans 896 90 0 0 wbs_dat_o[28]
port 621 nsew signal tristate
flabel metal2 s 130648 -960 130872 480 0 FreeSans 896 90 0 0 wbs_dat_o[29]
port 622 nsew signal tristate
flabel metal2 s 37688 -960 37912 480 0 FreeSans 896 90 0 0 wbs_dat_o[2]
port 623 nsew signal tristate
flabel metal2 s 134008 -960 134232 480 0 FreeSans 896 90 0 0 wbs_dat_o[30]
port 624 nsew signal tristate
flabel metal2 s 137368 -960 137592 480 0 FreeSans 896 90 0 0 wbs_dat_o[31]
port 625 nsew signal tristate
flabel metal2 s 42168 -960 42392 480 0 FreeSans 896 90 0 0 wbs_dat_o[3]
port 626 nsew signal tristate
flabel metal2 s 46648 -960 46872 480 0 FreeSans 896 90 0 0 wbs_dat_o[4]
port 627 nsew signal tristate
flabel metal2 s 50008 -960 50232 480 0 FreeSans 896 90 0 0 wbs_dat_o[5]
port 628 nsew signal tristate
flabel metal2 s 53368 -960 53592 480 0 FreeSans 896 90 0 0 wbs_dat_o[6]
port 629 nsew signal tristate
flabel metal2 s 56728 -960 56952 480 0 FreeSans 896 90 0 0 wbs_dat_o[7]
port 630 nsew signal tristate
flabel metal2 s 60088 -960 60312 480 0 FreeSans 896 90 0 0 wbs_dat_o[8]
port 631 nsew signal tristate
flabel metal2 s 63448 -960 63672 480 0 FreeSans 896 90 0 0 wbs_dat_o[9]
port 632 nsew signal tristate
flabel metal2 s 29848 -960 30072 480 0 FreeSans 896 90 0 0 wbs_sel_i[0]
port 633 nsew signal input
flabel metal2 s 34328 -960 34552 480 0 FreeSans 896 90 0 0 wbs_sel_i[1]
port 634 nsew signal input
flabel metal2 s 38808 -960 39032 480 0 FreeSans 896 90 0 0 wbs_sel_i[2]
port 635 nsew signal input
flabel metal2 s 43288 -960 43512 480 0 FreeSans 896 90 0 0 wbs_sel_i[3]
port 636 nsew signal input
flabel metal2 s 24248 -960 24472 480 0 FreeSans 896 90 0 0 wbs_stb_i
port 637 nsew signal input
flabel metal2 s 25368 -960 25592 480 0 FreeSans 896 90 0 0 wbs_we_i
port 638 nsew signal input
rlabel via4 57650 58322 57650 58322 0 vdd
rlabel via4 61370 64322 61370 64322 0 vss
rlabel metal4 196280 63224 196280 63224 0 clock_out\[0\]
rlabel metal2 67256 117558 67256 117558 0 clock_out\[1\]
rlabel metal2 68194 115864 68194 115864 0 clock_out\[2\]
rlabel metal2 69538 115864 69538 115864 0 clock_out\[3\]
rlabel metal2 70938 115864 70938 115864 0 clock_out\[4\]
rlabel metal2 76258 115864 76258 115864 0 clock_out\[8\]
rlabel metal2 77658 115864 77658 115864 0 clock_out\[9\]
rlabel metal3 520072 67802 520072 67802 0 clock_out_a
rlabel metal3 519554 84952 519554 84952 0 clock_out_b
rlabel metal3 516992 100856 516992 100856 0 clock_out_c
rlabel metal2 122696 144284 122696 144284 0 col_select_left\[0\]
rlabel metal2 190904 213696 190904 213696 0 col_select_left\[1\]
rlabel metal2 189672 235648 189672 235648 0 col_select_left\[2\]
rlabel metal2 188664 226408 188664 226408 0 col_select_left\[3\]
rlabel metal2 188552 302960 188552 302960 0 col_select_left\[4\]
rlabel metal2 188440 303072 188440 303072 0 col_select_left\[5\]
rlabel metal2 95480 116886 95480 116886 0 col_select_right\[0\]
rlabel metal2 96418 115864 96418 115864 0 col_select_right\[1\]
rlabel metal2 97818 115864 97818 115864 0 col_select_right\[2\]
rlabel metal2 99330 115864 99330 115864 0 col_select_right\[3\]
rlabel metal2 100982 115752 100982 115752 0 col_select_right\[4\]
rlabel metal2 101850 115864 101850 115864 0 col_select_right\[5\]
rlabel metal2 194936 148064 194936 148064 0 data_out_left\[0\]
rlabel metal2 146552 119350 146552 119350 0 data_out_left\[10\]
rlabel metal2 147896 118566 147896 118566 0 data_out_left\[11\]
rlabel metal2 149058 115864 149058 115864 0 data_out_left\[12\]
rlabel metal2 70392 158130 70392 158130 0 data_out_left\[13\]
rlabel metal3 195160 120008 195160 120008 0 data_out_left\[14\]
rlabel metal3 195160 124376 195160 124376 0 data_out_left\[15\]
rlabel metal2 24696 158186 24696 158186 0 data_out_left\[1\]
rlabel metal3 194600 147952 194600 147952 0 data_out_left\[2\]
rlabel metal3 89152 122584 89152 122584 0 data_out_left\[3\]
rlabel metal2 138138 115864 138138 115864 0 data_out_left\[4\]
rlabel metal2 139650 115864 139650 115864 0 data_out_left\[5\]
rlabel metal2 8232 235648 8232 235648 0 data_out_left\[6\]
rlabel metal2 142226 115864 142226 115864 0 data_out_left\[7\]
rlabel metal2 51282 160104 51282 160104 0 data_out_left\[8\]
rlabel metal2 145208 118118 145208 118118 0 data_out_left\[9\]
rlabel metal2 397880 234640 397880 234640 0 data_out_right\[0\]
rlabel metal2 125048 119294 125048 119294 0 data_out_right\[10\]
rlabel metal2 260792 153664 260792 153664 0 data_out_right\[11\]
rlabel metal2 356216 4704 356216 4704 0 data_out_right\[12\]
rlabel metal2 262136 154224 262136 154224 0 data_out_right\[13\]
rlabel metal4 195944 60144 195944 60144 0 data_out_right\[14\]
rlabel metal4 195832 146384 195832 146384 0 data_out_right\[15\]
rlabel metal2 397992 234696 397992 234696 0 data_out_right\[1\]
rlabel metal2 114296 135702 114296 135702 0 data_out_right\[2\]
rlabel metal2 115640 116830 115640 116830 0 data_out_right\[3\]
rlabel metal2 116984 117670 116984 117670 0 data_out_right\[4\]
rlabel metal2 117978 115864 117978 115864 0 data_out_right\[5\]
rlabel metal2 119490 115864 119490 115864 0 data_out_right\[6\]
rlabel metal2 121016 121086 121016 121086 0 data_out_right\[7\]
rlabel metal2 122360 120134 122360 120134 0 data_out_right\[8\]
rlabel metal2 123298 115864 123298 115864 0 data_out_right\[9\]
rlabel metal2 168056 116158 168056 116158 0 inverter_select\[0\]
rlabel metal2 168994 115864 168994 115864 0 inverter_select\[1\]
rlabel metal2 170338 115864 170338 115864 0 inverter_select\[2\]
rlabel metal2 171738 115864 171738 115864 0 inverter_select\[3\]
rlabel metal2 194600 210952 194600 210952 0 inverter_select\[4\]
rlabel metal4 195720 211848 195720 211848 0 inverter_select\[8\]
rlabel metal2 180334 115416 180334 115416 0 inverter_select\[9\]
rlabel metal3 37184 68600 37184 68600 0 io_control_trigger_oeb
rlabel metal3 1470 268856 1470 268856 0 io_in[31]
rlabel metal3 280 225176 280 225176 0 io_in[32]
rlabel metal3 1526 181832 1526 181832 0 io_in[33]
rlabel metal3 392 94472 392 94472 0 io_in[35]
rlabel metal2 35672 69538 35672 69538 0 io_in[36]
rlabel metal3 5726 29736 5726 29736 0 io_in[37]
rlabel metal3 569912 84546 569912 84546 0 io_in[8]
rlabel metal3 392 72688 392 72688 0 io_latch_data_oeb
rlabel metal3 5670 116648 5670 116648 0 io_miso_oeb
rlabel metal3 392 126728 392 126728 0 io_miso_out
rlabel metal3 3262 160104 3262 160104 0 io_mosi_oeb
rlabel metal3 589442 406728 589442 406728 0 io_oeb[10]
rlabel metal3 589386 451080 589386 451080 0 io_oeb[11]
rlabel metal3 591640 494648 591640 494648 0 io_oeb[12]
rlabel metal2 78008 69594 78008 69594 0 io_oeb[13]
rlabel metal2 75656 69538 75656 69538 0 io_oeb[14]
rlabel metal2 73304 68530 73304 68530 0 io_oeb[15]
rlabel metal2 467544 589386 467544 589386 0 io_oeb[16]
rlabel metal2 68600 69426 68600 69426 0 io_oeb[17]
rlabel metal4 190680 328216 190680 328216 0 io_oeb[20]
rlabel metal2 140728 589386 140728 589386 0 io_oeb[21]
rlabel metal2 75096 589442 75096 589442 0 io_oeb[22]
rlabel metal3 9968 587944 9968 587944 0 io_oeb[23]
rlabel metal3 4046 551208 4046 551208 0 io_oeb[24]
rlabel metal2 53816 69328 53816 69328 0 io_oeb[25]
rlabel metal2 52136 69314 52136 69314 0 io_oeb[26]
rlabel metal3 2310 420840 2310 420840 0 io_oeb[27]
rlabel metal3 2422 377384 2422 377384 0 io_oeb[28]
rlabel metal3 2590 333928 2590 333928 0 io_oeb[29]
rlabel metal2 192584 193088 192584 193088 0 io_oeb[8]
rlabel metal2 194264 189280 194264 189280 0 io_oeb[9]
rlabel metal2 403256 154770 403256 154770 0 io_out[10]
rlabel metal2 407736 317912 407736 317912 0 io_out[11]
rlabel metal2 404040 319592 404040 319592 0 io_out[12]
rlabel metal2 196504 453264 196504 453264 0 io_out[20]
rlabel metal2 189000 453264 189000 453264 0 io_out[21]
rlabel metal2 91448 589386 91448 589386 0 io_out[22]
rlabel metal2 26040 589498 26040 589498 0 io_out[23]
rlabel metal3 392 561568 392 561568 0 io_out[24]
rlabel metal3 392 518000 392 518000 0 io_out[25]
rlabel metal3 3150 475160 3150 475160 0 io_out[26]
rlabel metal3 3192 320992 3192 320992 0 io_out[27]
rlabel metal3 2366 388248 2366 388248 0 io_out[28]
rlabel metal3 2478 344792 2478 344792 0 io_out[29]
rlabel metal3 590786 351288 590786 351288 0 io_out[9]
rlabel metal3 392 7336 392 7336 0 io_reset_n_oeb
rlabel metal3 10640 30184 10640 30184 0 io_sclk_oeb
rlabel metal3 10696 54824 10696 54824 0 io_ss_n_oeb
rlabel metal3 2534 290472 2534 290472 0 io_update_cycle_complete_oeb
rlabel metal2 31192 68992 31192 68992 0 io_update_cycle_complete_out
rlabel metal2 138488 4158 138488 4158 0 la_data_in[0]
rlabel metal2 171696 392 171696 392 0 la_data_in[10]
rlabel metal2 159978 70056 159978 70056 0 la_data_in[11]
rlabel metal3 163240 65576 163240 65576 0 la_data_in[12]
rlabel metal2 165032 67410 165032 67410 0 la_data_in[13]
rlabel metal2 166866 70056 166866 70056 0 la_data_in[14]
rlabel metal2 169736 40586 169736 40586 0 la_data_in[15]
rlabel metal2 191856 392 191856 392 0 la_data_in[16]
rlabel metal2 195216 392 195216 392 0 la_data_in[17]
rlabel metal2 47880 15498 47880 15498 0 la_data_in[18]
rlabel metal2 53368 18858 53368 18858 0 la_data_in[19]
rlabel metal2 141848 4214 141848 4214 0 la_data_in[1]
rlabel metal3 202160 4536 202160 4536 0 la_data_in[20]
rlabel metal3 141512 7448 141512 7448 0 la_data_in[2]
rlabel metal3 144872 6776 144872 6776 0 la_data_in[3]
rlabel metal2 143346 70056 143346 70056 0 la_data_in[4]
rlabel metal3 147112 65912 147112 65912 0 la_data_in[5]
rlabel metal2 148218 70056 148218 70056 0 la_data_in[6]
rlabel metal2 162008 2702 162008 2702 0 la_data_in[7]
rlabel metal3 164696 4424 164696 4424 0 la_data_in[8]
rlabel metal2 168952 2254 168952 2254 0 la_data_in[9]
rlabel metal2 91434 70056 91434 70056 0 la_oenb[0]
rlabel metal3 116200 65576 116200 65576 0 la_oenb[10]
rlabel metal2 117810 70056 117810 70056 0 la_oenb[11]
rlabel metal2 119826 70056 119826 70056 0 la_oenb[12]
rlabel metal2 122696 38010 122696 38010 0 la_oenb[13]
rlabel metal2 124698 70056 124698 70056 0 la_oenb[14]
rlabel metal2 191128 4830 191128 4830 0 la_oenb[15]
rlabel metal3 192640 4088 192640 4088 0 la_oenb[16]
rlabel metal2 20440 18802 20440 18802 0 la_oenb[17]
rlabel metal2 25578 20104 25578 20104 0 la_oenb[18]
rlabel metal2 30842 20104 30842 20104 0 la_oenb[19]
rlabel metal2 94290 70056 94290 70056 0 la_oenb[1]
rlabel metal4 198968 4032 198968 4032 0 la_oenb[20]
rlabel metal2 147448 2478 147448 2478 0 la_oenb[2]
rlabel metal2 99176 45570 99176 45570 0 la_oenb[3]
rlabel metal2 101178 70056 101178 70056 0 la_oenb[4]
rlabel metal2 145320 13720 145320 13720 0 la_oenb[5]
rlabel metal2 352632 3150 352632 3150 0 la_oenb[63]
rlabel metal2 106050 70056 106050 70056 0 la_oenb[6]
rlabel metal2 164248 2646 164248 2646 0 la_oenb[7]
rlabel metal2 167608 2478 167608 2478 0 la_oenb[8]
rlabel metal3 166544 4760 166544 4760 0 la_oenb[9]
rlabel metal2 43848 134232 43848 134232 0 mem_address_left\[0\]
rlabel metal2 40376 117166 40376 117166 0 mem_address_left\[1\]
rlabel metal2 6664 232680 6664 232680 0 mem_address_left\[2\]
rlabel metal2 6440 229320 6440 229320 0 mem_address_left\[3\]
rlabel metal2 44408 119742 44408 119742 0 mem_address_left\[4\]
rlabel metal2 45752 117222 45752 117222 0 mem_address_left\[5\]
rlabel metal2 47096 118174 47096 118174 0 mem_address_left\[6\]
rlabel metal2 48090 115864 48090 115864 0 mem_address_left\[7\]
rlabel metal2 49784 117446 49784 117446 0 mem_address_left\[8\]
rlabel metal2 50778 115864 50778 115864 0 mem_address_left\[9\]
rlabel metal2 25592 117614 25592 117614 0 mem_address_right\[0\]
rlabel metal2 26936 127246 26936 127246 0 mem_address_right\[1\]
rlabel metal2 27874 115864 27874 115864 0 mem_address_right\[2\]
rlabel metal2 29218 115864 29218 115864 0 mem_address_right\[3\]
rlabel metal2 30968 118454 30968 118454 0 mem_address_right\[4\]
rlabel metal4 397656 230104 397656 230104 0 mem_address_right\[5\]
rlabel metal2 194712 61208 194712 61208 0 mem_address_right\[6\]
rlabel metal3 497448 151144 497448 151144 0 mem_address_right\[7\]
rlabel metal4 195720 61320 195720 61320 0 mem_address_right\[8\]
rlabel metal2 37338 115864 37338 115864 0 mem_address_right\[9\]
rlabel metal2 52472 116774 52472 116774 0 mem_write_n\[0\]
rlabel metal2 53816 117278 53816 117278 0 mem_write_n\[1\]
rlabel metal2 54754 115864 54754 115864 0 mem_write_n\[2\]
rlabel metal2 119602 320040 119602 320040 0 mem_write_n\[3\]
rlabel metal2 194712 219408 194712 219408 0 mem_write_n\[4\]
rlabel metal2 195720 236992 195720 236992 0 mem_write_n\[8\]
rlabel metal2 64218 115864 64218 115864 0 mem_write_n\[9\]
rlabel metal2 24248 117558 24248 117558 0 output_active_left
rlabel metal2 22498 115864 22498 115864 0 output_active_right
rlabel metal2 194152 62608 194152 62608 0 row_col_select\[0\]
rlabel metal2 155960 119686 155960 119686 0 row_col_select\[1\]
rlabel metal2 156898 115864 156898 115864 0 row_col_select\[2\]
rlabel metal2 188328 233016 188328 233016 0 row_col_select\[3\]
rlabel metal4 189224 228536 189224 228536 0 row_col_select\[4\]
rlabel metal2 165368 117222 165368 117222 0 row_col_select\[8\]
rlabel metal2 166530 115864 166530 115864 0 row_col_select\[9\]
rlabel metal2 190680 235536 190680 235536 0 row_select_left\[0\]
rlabel metal2 191016 235200 191016 235200 0 row_select_left\[1\]
rlabel metal2 161966 160104 161966 160104 0 row_select_left\[2\]
rlabel metal2 91448 120526 91448 120526 0 row_select_left\[3\]
rlabel metal2 92792 118062 92792 118062 0 row_select_left\[4\]
rlabel metal2 94136 121366 94136 121366 0 row_select_left\[5\]
rlabel metal2 544152 155274 544152 155274 0 row_select_right\[0\]
rlabel metal2 547736 155848 547736 155848 0 row_select_right\[1\]
rlabel metal2 82040 116046 82040 116046 0 row_select_right\[2\]
rlabel metal2 82978 115864 82978 115864 0 row_select_right\[3\]
rlabel metal2 84378 115864 84378 115864 0 row_select_right\[4\]
rlabel metal2 192696 63448 192696 63448 0 row_select_right\[5\]
rlabel metal2 6664 46200 6664 46200 0 spi_data\[0\]
rlabel metal4 22232 82572 22232 82572 0 spi_data\[10\]
rlabel metal3 18858 87528 18858 87528 0 spi_data\[11\]
rlabel metal3 20426 88872 20426 88872 0 spi_data\[12\]
rlabel metal3 20650 90216 20650 90216 0 spi_data\[13\]
rlabel metal3 20874 91560 20874 91560 0 spi_data\[14\]
rlabel metal3 18914 92904 18914 92904 0 spi_data\[15\]
rlabel metal3 20706 94248 20706 94248 0 spi_data\[16\]
rlabel metal3 20426 95592 20426 95592 0 spi_data\[17\]
rlabel metal3 20650 96936 20650 96936 0 spi_data\[18\]
rlabel metal3 20706 98280 20706 98280 0 spi_data\[19\]
rlabel metal2 6552 47656 6552 47656 0 spi_data\[1\]
rlabel metal3 20594 99624 20594 99624 0 spi_data\[20\]
rlabel metal3 20818 100968 20818 100968 0 spi_data\[21\]
rlabel metal3 18970 102312 18970 102312 0 spi_data\[22\]
rlabel metal3 20986 103656 20986 103656 0 spi_data\[23\]
rlabel metal3 21042 105000 21042 105000 0 spi_data\[24\]
rlabel metal3 20930 106344 20930 106344 0 spi_data\[25\]
rlabel metal3 20538 107688 20538 107688 0 spi_data\[26\]
rlabel metal3 20762 109032 20762 109032 0 spi_data\[27\]
rlabel metal3 20818 110376 20818 110376 0 spi_data\[28\]
rlabel metal3 20874 111720 20874 111720 0 spi_data\[29\]
rlabel metal3 21672 74914 21672 74914 0 spi_data\[2\]
rlabel metal3 20482 113064 20482 113064 0 spi_data\[30\]
rlabel metal3 28840 68432 28840 68432 0 spi_data\[31\]
rlabel metal3 21672 76202 21672 76202 0 spi_data\[3\]
rlabel metal3 21672 77714 21672 77714 0 spi_data\[4\]
rlabel metal2 4984 50232 4984 50232 0 spi_data\[5\]
rlabel metal3 20930 80808 20930 80808 0 spi_data\[6\]
rlabel metal4 22568 82152 22568 82152 0 spi_data\[7\]
rlabel metal3 20986 83496 20986 83496 0 spi_data\[8\]
rlabel metal3 20034 84840 20034 84840 0 spi_data\[9\]
rlabel metal4 61880 20944 61880 20944 0 spi_data_clock
rlabel metal2 568176 392 568176 392 0 user_clock2
<< properties >>
string FIXED_BBOX 0 0 592040 592040
<< end >>

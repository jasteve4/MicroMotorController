magic
tech gf180mcuC
magscale 1 5
timestamp 1670301663
<< obsm1 >>
rect 5172 6538 288820 230198
<< metal2 >>
rect 4844 295780 4956 296500
rect 13020 295780 13132 296500
rect 21196 295780 21308 296500
rect 29372 295780 29484 296500
rect 37548 295780 37660 296500
rect 45724 295780 45836 296500
rect 53900 295780 54012 296500
rect 62076 295780 62188 296500
rect 70252 295780 70364 296500
rect 78428 295780 78540 296500
rect 86604 295780 86716 296500
rect 94780 295780 94892 296500
rect 102956 295780 103068 296500
rect 111132 295780 111244 296500
rect 119308 295780 119420 296500
rect 127484 295780 127596 296500
rect 135660 295780 135772 296500
rect 143836 295780 143948 296500
rect 152012 295780 152124 296500
rect 160188 295780 160300 296500
rect 168364 295780 168476 296500
rect 176540 295780 176652 296500
rect 184716 295780 184828 296500
rect 192892 295780 193004 296500
rect 201068 295780 201180 296500
rect 209244 295780 209356 296500
rect 217420 295780 217532 296500
rect 225596 295780 225708 296500
rect 233772 295780 233884 296500
rect 241948 295780 242060 296500
rect 250124 295780 250236 296500
rect 258300 295780 258412 296500
rect 266476 295780 266588 296500
rect 274652 295780 274764 296500
rect 282828 295780 282940 296500
rect 291004 295780 291116 296500
rect 9884 -480 9996 240
rect 10444 -480 10556 240
rect 11004 -480 11116 240
rect 11564 -480 11676 240
rect 12124 -480 12236 240
rect 12684 -480 12796 240
rect 13244 -480 13356 240
rect 13804 -480 13916 240
rect 14364 -480 14476 240
rect 14924 -480 15036 240
rect 15484 -480 15596 240
rect 16044 -480 16156 240
rect 16604 -480 16716 240
rect 17164 -480 17276 240
rect 17724 -480 17836 240
rect 18284 -480 18396 240
rect 18844 -480 18956 240
rect 19404 -480 19516 240
rect 19964 -480 20076 240
rect 20524 -480 20636 240
rect 21084 -480 21196 240
rect 21644 -480 21756 240
rect 22204 -480 22316 240
rect 22764 -480 22876 240
rect 23324 -480 23436 240
rect 23884 -480 23996 240
rect 24444 -480 24556 240
rect 25004 -480 25116 240
rect 25564 -480 25676 240
rect 26124 -480 26236 240
rect 26684 -480 26796 240
rect 27244 -480 27356 240
rect 27804 -480 27916 240
rect 28364 -480 28476 240
rect 28924 -480 29036 240
rect 29484 -480 29596 240
rect 30044 -480 30156 240
rect 30604 -480 30716 240
rect 31164 -480 31276 240
rect 31724 -480 31836 240
rect 32284 -480 32396 240
rect 32844 -480 32956 240
rect 33404 -480 33516 240
rect 33964 -480 34076 240
rect 34524 -480 34636 240
rect 35084 -480 35196 240
rect 35644 -480 35756 240
rect 36204 -480 36316 240
rect 36764 -480 36876 240
rect 37324 -480 37436 240
rect 37884 -480 37996 240
rect 38444 -480 38556 240
rect 39004 -480 39116 240
rect 39564 -480 39676 240
rect 40124 -480 40236 240
rect 40684 -480 40796 240
rect 41244 -480 41356 240
rect 41804 -480 41916 240
rect 42364 -480 42476 240
rect 42924 -480 43036 240
rect 43484 -480 43596 240
rect 44044 -480 44156 240
rect 44604 -480 44716 240
rect 45164 -480 45276 240
rect 45724 -480 45836 240
rect 46284 -480 46396 240
rect 46844 -480 46956 240
rect 47404 -480 47516 240
rect 47964 -480 48076 240
rect 48524 -480 48636 240
rect 49084 -480 49196 240
rect 49644 -480 49756 240
rect 50204 -480 50316 240
rect 50764 -480 50876 240
rect 51324 -480 51436 240
rect 51884 -480 51996 240
rect 52444 -480 52556 240
rect 53004 -480 53116 240
rect 53564 -480 53676 240
rect 54124 -480 54236 240
rect 54684 -480 54796 240
rect 55244 -480 55356 240
rect 55804 -480 55916 240
rect 56364 -480 56476 240
rect 56924 -480 57036 240
rect 57484 -480 57596 240
rect 58044 -480 58156 240
rect 58604 -480 58716 240
rect 59164 -480 59276 240
rect 59724 -480 59836 240
rect 60284 -480 60396 240
rect 60844 -480 60956 240
rect 61404 -480 61516 240
rect 61964 -480 62076 240
rect 62524 -480 62636 240
rect 63084 -480 63196 240
rect 63644 -480 63756 240
rect 64204 -480 64316 240
rect 64764 -480 64876 240
rect 65324 -480 65436 240
rect 65884 -480 65996 240
rect 66444 -480 66556 240
rect 67004 -480 67116 240
rect 67564 -480 67676 240
rect 68124 -480 68236 240
rect 68684 -480 68796 240
rect 69244 -480 69356 240
rect 69804 -480 69916 240
rect 70364 -480 70476 240
rect 70924 -480 71036 240
rect 71484 -480 71596 240
rect 72044 -480 72156 240
rect 72604 -480 72716 240
rect 73164 -480 73276 240
rect 73724 -480 73836 240
rect 74284 -480 74396 240
rect 74844 -480 74956 240
rect 75404 -480 75516 240
rect 75964 -480 76076 240
rect 76524 -480 76636 240
rect 77084 -480 77196 240
rect 77644 -480 77756 240
rect 78204 -480 78316 240
rect 78764 -480 78876 240
rect 79324 -480 79436 240
rect 79884 -480 79996 240
rect 80444 -480 80556 240
rect 81004 -480 81116 240
rect 81564 -480 81676 240
rect 82124 -480 82236 240
rect 82684 -480 82796 240
rect 83244 -480 83356 240
rect 83804 -480 83916 240
rect 84364 -480 84476 240
rect 84924 -480 85036 240
rect 85484 -480 85596 240
rect 86044 -480 86156 240
rect 86604 -480 86716 240
rect 87164 -480 87276 240
rect 87724 -480 87836 240
rect 88284 -480 88396 240
rect 88844 -480 88956 240
rect 89404 -480 89516 240
rect 89964 -480 90076 240
rect 90524 -480 90636 240
rect 91084 -480 91196 240
rect 91644 -480 91756 240
rect 92204 -480 92316 240
rect 92764 -480 92876 240
rect 93324 -480 93436 240
rect 93884 -480 93996 240
rect 94444 -480 94556 240
rect 95004 -480 95116 240
rect 95564 -480 95676 240
rect 96124 -480 96236 240
rect 96684 -480 96796 240
rect 97244 -480 97356 240
rect 97804 -480 97916 240
rect 98364 -480 98476 240
rect 98924 -480 99036 240
rect 99484 -480 99596 240
rect 100044 -480 100156 240
rect 100604 -480 100716 240
rect 101164 -480 101276 240
rect 101724 -480 101836 240
rect 102284 -480 102396 240
rect 102844 -480 102956 240
rect 103404 -480 103516 240
rect 103964 -480 104076 240
rect 104524 -480 104636 240
rect 105084 -480 105196 240
rect 105644 -480 105756 240
rect 106204 -480 106316 240
rect 106764 -480 106876 240
rect 107324 -480 107436 240
rect 107884 -480 107996 240
rect 108444 -480 108556 240
rect 109004 -480 109116 240
rect 109564 -480 109676 240
rect 110124 -480 110236 240
rect 110684 -480 110796 240
rect 111244 -480 111356 240
rect 111804 -480 111916 240
rect 112364 -480 112476 240
rect 112924 -480 113036 240
rect 113484 -480 113596 240
rect 114044 -480 114156 240
rect 114604 -480 114716 240
rect 115164 -480 115276 240
rect 115724 -480 115836 240
rect 116284 -480 116396 240
rect 116844 -480 116956 240
rect 117404 -480 117516 240
rect 117964 -480 118076 240
rect 118524 -480 118636 240
rect 119084 -480 119196 240
rect 119644 -480 119756 240
rect 120204 -480 120316 240
rect 120764 -480 120876 240
rect 121324 -480 121436 240
rect 121884 -480 121996 240
rect 122444 -480 122556 240
rect 123004 -480 123116 240
rect 123564 -480 123676 240
rect 124124 -480 124236 240
rect 124684 -480 124796 240
rect 125244 -480 125356 240
rect 125804 -480 125916 240
rect 126364 -480 126476 240
rect 126924 -480 127036 240
rect 127484 -480 127596 240
rect 128044 -480 128156 240
rect 128604 -480 128716 240
rect 129164 -480 129276 240
rect 129724 -480 129836 240
rect 130284 -480 130396 240
rect 130844 -480 130956 240
rect 131404 -480 131516 240
rect 131964 -480 132076 240
rect 132524 -480 132636 240
rect 133084 -480 133196 240
rect 133644 -480 133756 240
rect 134204 -480 134316 240
rect 134764 -480 134876 240
rect 135324 -480 135436 240
rect 135884 -480 135996 240
rect 136444 -480 136556 240
rect 137004 -480 137116 240
rect 137564 -480 137676 240
rect 138124 -480 138236 240
rect 138684 -480 138796 240
rect 139244 -480 139356 240
rect 139804 -480 139916 240
rect 140364 -480 140476 240
rect 140924 -480 141036 240
rect 141484 -480 141596 240
rect 142044 -480 142156 240
rect 142604 -480 142716 240
rect 143164 -480 143276 240
rect 143724 -480 143836 240
rect 144284 -480 144396 240
rect 144844 -480 144956 240
rect 145404 -480 145516 240
rect 145964 -480 146076 240
rect 146524 -480 146636 240
rect 147084 -480 147196 240
rect 147644 -480 147756 240
rect 148204 -480 148316 240
rect 148764 -480 148876 240
rect 149324 -480 149436 240
rect 149884 -480 149996 240
rect 150444 -480 150556 240
rect 151004 -480 151116 240
rect 151564 -480 151676 240
rect 152124 -480 152236 240
rect 152684 -480 152796 240
rect 153244 -480 153356 240
rect 153804 -480 153916 240
rect 154364 -480 154476 240
rect 154924 -480 155036 240
rect 155484 -480 155596 240
rect 156044 -480 156156 240
rect 156604 -480 156716 240
rect 157164 -480 157276 240
rect 157724 -480 157836 240
rect 158284 -480 158396 240
rect 158844 -480 158956 240
rect 159404 -480 159516 240
rect 159964 -480 160076 240
rect 160524 -480 160636 240
rect 161084 -480 161196 240
rect 161644 -480 161756 240
rect 162204 -480 162316 240
rect 162764 -480 162876 240
rect 163324 -480 163436 240
rect 163884 -480 163996 240
rect 164444 -480 164556 240
rect 165004 -480 165116 240
rect 165564 -480 165676 240
rect 166124 -480 166236 240
rect 166684 -480 166796 240
rect 167244 -480 167356 240
rect 167804 -480 167916 240
rect 168364 -480 168476 240
rect 168924 -480 169036 240
rect 169484 -480 169596 240
rect 170044 -480 170156 240
rect 170604 -480 170716 240
rect 171164 -480 171276 240
rect 171724 -480 171836 240
rect 172284 -480 172396 240
rect 172844 -480 172956 240
rect 173404 -480 173516 240
rect 173964 -480 174076 240
rect 174524 -480 174636 240
rect 175084 -480 175196 240
rect 175644 -480 175756 240
rect 176204 -480 176316 240
rect 176764 -480 176876 240
rect 177324 -480 177436 240
rect 177884 -480 177996 240
rect 178444 -480 178556 240
rect 179004 -480 179116 240
rect 179564 -480 179676 240
rect 180124 -480 180236 240
rect 180684 -480 180796 240
rect 181244 -480 181356 240
rect 181804 -480 181916 240
rect 182364 -480 182476 240
rect 182924 -480 183036 240
rect 183484 -480 183596 240
rect 184044 -480 184156 240
rect 184604 -480 184716 240
rect 185164 -480 185276 240
rect 185724 -480 185836 240
rect 186284 -480 186396 240
rect 186844 -480 186956 240
rect 187404 -480 187516 240
rect 187964 -480 188076 240
rect 188524 -480 188636 240
rect 189084 -480 189196 240
rect 189644 -480 189756 240
rect 190204 -480 190316 240
rect 190764 -480 190876 240
rect 191324 -480 191436 240
rect 191884 -480 191996 240
rect 192444 -480 192556 240
rect 193004 -480 193116 240
rect 193564 -480 193676 240
rect 194124 -480 194236 240
rect 194684 -480 194796 240
rect 195244 -480 195356 240
rect 195804 -480 195916 240
rect 196364 -480 196476 240
rect 196924 -480 197036 240
rect 197484 -480 197596 240
rect 198044 -480 198156 240
rect 198604 -480 198716 240
rect 199164 -480 199276 240
rect 199724 -480 199836 240
rect 200284 -480 200396 240
rect 200844 -480 200956 240
rect 201404 -480 201516 240
rect 201964 -480 202076 240
rect 202524 -480 202636 240
rect 203084 -480 203196 240
rect 203644 -480 203756 240
rect 204204 -480 204316 240
rect 204764 -480 204876 240
rect 205324 -480 205436 240
rect 205884 -480 205996 240
rect 206444 -480 206556 240
rect 207004 -480 207116 240
rect 207564 -480 207676 240
rect 208124 -480 208236 240
rect 208684 -480 208796 240
rect 209244 -480 209356 240
rect 209804 -480 209916 240
rect 210364 -480 210476 240
rect 210924 -480 211036 240
rect 211484 -480 211596 240
rect 212044 -480 212156 240
rect 212604 -480 212716 240
rect 213164 -480 213276 240
rect 213724 -480 213836 240
rect 214284 -480 214396 240
rect 214844 -480 214956 240
rect 215404 -480 215516 240
rect 215964 -480 216076 240
rect 216524 -480 216636 240
rect 217084 -480 217196 240
rect 217644 -480 217756 240
rect 218204 -480 218316 240
rect 218764 -480 218876 240
rect 219324 -480 219436 240
rect 219884 -480 219996 240
rect 220444 -480 220556 240
rect 221004 -480 221116 240
rect 221564 -480 221676 240
rect 222124 -480 222236 240
rect 222684 -480 222796 240
rect 223244 -480 223356 240
rect 223804 -480 223916 240
rect 224364 -480 224476 240
rect 224924 -480 225036 240
rect 225484 -480 225596 240
rect 226044 -480 226156 240
rect 226604 -480 226716 240
rect 227164 -480 227276 240
rect 227724 -480 227836 240
rect 228284 -480 228396 240
rect 228844 -480 228956 240
rect 229404 -480 229516 240
rect 229964 -480 230076 240
rect 230524 -480 230636 240
rect 231084 -480 231196 240
rect 231644 -480 231756 240
rect 232204 -480 232316 240
rect 232764 -480 232876 240
rect 233324 -480 233436 240
rect 233884 -480 233996 240
rect 234444 -480 234556 240
rect 235004 -480 235116 240
rect 235564 -480 235676 240
rect 236124 -480 236236 240
rect 236684 -480 236796 240
rect 237244 -480 237356 240
rect 237804 -480 237916 240
rect 238364 -480 238476 240
rect 238924 -480 239036 240
rect 239484 -480 239596 240
rect 240044 -480 240156 240
rect 240604 -480 240716 240
rect 241164 -480 241276 240
rect 241724 -480 241836 240
rect 242284 -480 242396 240
rect 242844 -480 242956 240
rect 243404 -480 243516 240
rect 243964 -480 244076 240
rect 244524 -480 244636 240
rect 245084 -480 245196 240
rect 245644 -480 245756 240
rect 246204 -480 246316 240
rect 246764 -480 246876 240
rect 247324 -480 247436 240
rect 247884 -480 247996 240
rect 248444 -480 248556 240
rect 249004 -480 249116 240
rect 249564 -480 249676 240
rect 250124 -480 250236 240
rect 250684 -480 250796 240
rect 251244 -480 251356 240
rect 251804 -480 251916 240
rect 252364 -480 252476 240
rect 252924 -480 253036 240
rect 253484 -480 253596 240
rect 254044 -480 254156 240
rect 254604 -480 254716 240
rect 255164 -480 255276 240
rect 255724 -480 255836 240
rect 256284 -480 256396 240
rect 256844 -480 256956 240
rect 257404 -480 257516 240
rect 257964 -480 258076 240
rect 258524 -480 258636 240
rect 259084 -480 259196 240
rect 259644 -480 259756 240
rect 260204 -480 260316 240
rect 260764 -480 260876 240
rect 261324 -480 261436 240
rect 261884 -480 261996 240
rect 262444 -480 262556 240
rect 263004 -480 263116 240
rect 263564 -480 263676 240
rect 264124 -480 264236 240
rect 264684 -480 264796 240
rect 265244 -480 265356 240
rect 265804 -480 265916 240
rect 266364 -480 266476 240
rect 266924 -480 267036 240
rect 267484 -480 267596 240
rect 268044 -480 268156 240
rect 268604 -480 268716 240
rect 269164 -480 269276 240
rect 269724 -480 269836 240
rect 270284 -480 270396 240
rect 270844 -480 270956 240
rect 271404 -480 271516 240
rect 271964 -480 272076 240
rect 272524 -480 272636 240
rect 273084 -480 273196 240
rect 273644 -480 273756 240
rect 274204 -480 274316 240
rect 274764 -480 274876 240
rect 275324 -480 275436 240
rect 275884 -480 275996 240
rect 276444 -480 276556 240
rect 277004 -480 277116 240
rect 277564 -480 277676 240
rect 278124 -480 278236 240
rect 278684 -480 278796 240
rect 279244 -480 279356 240
rect 279804 -480 279916 240
rect 280364 -480 280476 240
rect 280924 -480 281036 240
rect 281484 -480 281596 240
rect 282044 -480 282156 240
rect 282604 -480 282716 240
rect 283164 -480 283276 240
rect 283724 -480 283836 240
rect 284284 -480 284396 240
rect 284844 -480 284956 240
rect 285404 -480 285516 240
rect 285964 -480 286076 240
<< obsm2 >>
rect 14 295750 4814 295834
rect 4986 295750 12990 295834
rect 13162 295750 21166 295834
rect 21338 295750 29342 295834
rect 29514 295750 37518 295834
rect 37690 295750 45694 295834
rect 45866 295750 53870 295834
rect 54042 295750 62046 295834
rect 62218 295750 70222 295834
rect 70394 295750 78398 295834
rect 78570 295750 86574 295834
rect 86746 295750 94750 295834
rect 94922 295750 102926 295834
rect 103098 295750 111102 295834
rect 111274 295750 119278 295834
rect 119450 295750 127454 295834
rect 127626 295750 135630 295834
rect 135802 295750 143806 295834
rect 143978 295750 151982 295834
rect 152154 295750 160158 295834
rect 160330 295750 168334 295834
rect 168506 295750 176510 295834
rect 176682 295750 184686 295834
rect 184858 295750 192862 295834
rect 193034 295750 201038 295834
rect 201210 295750 209214 295834
rect 209386 295750 217390 295834
rect 217562 295750 225566 295834
rect 225738 295750 233742 295834
rect 233914 295750 241918 295834
rect 242090 295750 250094 295834
rect 250266 295750 258270 295834
rect 258442 295750 266446 295834
rect 266618 295750 274622 295834
rect 274794 295750 282798 295834
rect 282970 295750 290974 295834
rect 291146 295750 295050 295834
rect 14 270 295050 295750
rect 14 182 9854 270
rect 10026 182 10414 270
rect 10586 182 10974 270
rect 11146 182 11534 270
rect 11706 182 12094 270
rect 12266 182 12654 270
rect 12826 182 13214 270
rect 13386 182 13774 270
rect 13946 182 14334 270
rect 14506 182 14894 270
rect 15066 182 15454 270
rect 15626 182 16014 270
rect 16186 182 16574 270
rect 16746 182 17134 270
rect 17306 182 17694 270
rect 17866 182 18254 270
rect 18426 182 18814 270
rect 18986 182 19374 270
rect 19546 182 19934 270
rect 20106 182 20494 270
rect 20666 182 21054 270
rect 21226 182 21614 270
rect 21786 182 22174 270
rect 22346 182 22734 270
rect 22906 182 23294 270
rect 23466 182 23854 270
rect 24026 182 24414 270
rect 24586 182 24974 270
rect 25146 182 25534 270
rect 25706 182 26094 270
rect 26266 182 26654 270
rect 26826 182 27214 270
rect 27386 182 27774 270
rect 27946 182 28334 270
rect 28506 182 28894 270
rect 29066 182 29454 270
rect 29626 182 30014 270
rect 30186 182 30574 270
rect 30746 182 31134 270
rect 31306 182 31694 270
rect 31866 182 32254 270
rect 32426 182 32814 270
rect 32986 182 33374 270
rect 33546 182 33934 270
rect 34106 182 34494 270
rect 34666 182 35054 270
rect 35226 182 35614 270
rect 35786 182 36174 270
rect 36346 182 36734 270
rect 36906 182 37294 270
rect 37466 182 37854 270
rect 38026 182 38414 270
rect 38586 182 38974 270
rect 39146 182 39534 270
rect 39706 182 40094 270
rect 40266 182 40654 270
rect 40826 182 41214 270
rect 41386 182 41774 270
rect 41946 182 42334 270
rect 42506 182 42894 270
rect 43066 182 43454 270
rect 43626 182 44014 270
rect 44186 182 44574 270
rect 44746 182 45134 270
rect 45306 182 45694 270
rect 45866 182 46254 270
rect 46426 182 46814 270
rect 46986 182 47374 270
rect 47546 182 47934 270
rect 48106 182 48494 270
rect 48666 182 49054 270
rect 49226 182 49614 270
rect 49786 182 50174 270
rect 50346 182 50734 270
rect 50906 182 51294 270
rect 51466 182 51854 270
rect 52026 182 52414 270
rect 52586 182 52974 270
rect 53146 182 53534 270
rect 53706 182 54094 270
rect 54266 182 54654 270
rect 54826 182 55214 270
rect 55386 182 55774 270
rect 55946 182 56334 270
rect 56506 182 56894 270
rect 57066 182 57454 270
rect 57626 182 58014 270
rect 58186 182 58574 270
rect 58746 182 59134 270
rect 59306 182 59694 270
rect 59866 182 60254 270
rect 60426 182 60814 270
rect 60986 182 61374 270
rect 61546 182 61934 270
rect 62106 182 62494 270
rect 62666 182 63054 270
rect 63226 182 63614 270
rect 63786 182 64174 270
rect 64346 182 64734 270
rect 64906 182 65294 270
rect 65466 182 65854 270
rect 66026 182 66414 270
rect 66586 182 66974 270
rect 67146 182 67534 270
rect 67706 182 68094 270
rect 68266 182 68654 270
rect 68826 182 69214 270
rect 69386 182 69774 270
rect 69946 182 70334 270
rect 70506 182 70894 270
rect 71066 182 71454 270
rect 71626 182 72014 270
rect 72186 182 72574 270
rect 72746 182 73134 270
rect 73306 182 73694 270
rect 73866 182 74254 270
rect 74426 182 74814 270
rect 74986 182 75374 270
rect 75546 182 75934 270
rect 76106 182 76494 270
rect 76666 182 77054 270
rect 77226 182 77614 270
rect 77786 182 78174 270
rect 78346 182 78734 270
rect 78906 182 79294 270
rect 79466 182 79854 270
rect 80026 182 80414 270
rect 80586 182 80974 270
rect 81146 182 81534 270
rect 81706 182 82094 270
rect 82266 182 82654 270
rect 82826 182 83214 270
rect 83386 182 83774 270
rect 83946 182 84334 270
rect 84506 182 84894 270
rect 85066 182 85454 270
rect 85626 182 86014 270
rect 86186 182 86574 270
rect 86746 182 87134 270
rect 87306 182 87694 270
rect 87866 182 88254 270
rect 88426 182 88814 270
rect 88986 182 89374 270
rect 89546 182 89934 270
rect 90106 182 90494 270
rect 90666 182 91054 270
rect 91226 182 91614 270
rect 91786 182 92174 270
rect 92346 182 92734 270
rect 92906 182 93294 270
rect 93466 182 93854 270
rect 94026 182 94414 270
rect 94586 182 94974 270
rect 95146 182 95534 270
rect 95706 182 96094 270
rect 96266 182 96654 270
rect 96826 182 97214 270
rect 97386 182 97774 270
rect 97946 182 98334 270
rect 98506 182 98894 270
rect 99066 182 99454 270
rect 99626 182 100014 270
rect 100186 182 100574 270
rect 100746 182 101134 270
rect 101306 182 101694 270
rect 101866 182 102254 270
rect 102426 182 102814 270
rect 102986 182 103374 270
rect 103546 182 103934 270
rect 104106 182 104494 270
rect 104666 182 105054 270
rect 105226 182 105614 270
rect 105786 182 106174 270
rect 106346 182 106734 270
rect 106906 182 107294 270
rect 107466 182 107854 270
rect 108026 182 108414 270
rect 108586 182 108974 270
rect 109146 182 109534 270
rect 109706 182 110094 270
rect 110266 182 110654 270
rect 110826 182 111214 270
rect 111386 182 111774 270
rect 111946 182 112334 270
rect 112506 182 112894 270
rect 113066 182 113454 270
rect 113626 182 114014 270
rect 114186 182 114574 270
rect 114746 182 115134 270
rect 115306 182 115694 270
rect 115866 182 116254 270
rect 116426 182 116814 270
rect 116986 182 117374 270
rect 117546 182 117934 270
rect 118106 182 118494 270
rect 118666 182 119054 270
rect 119226 182 119614 270
rect 119786 182 120174 270
rect 120346 182 120734 270
rect 120906 182 121294 270
rect 121466 182 121854 270
rect 122026 182 122414 270
rect 122586 182 122974 270
rect 123146 182 123534 270
rect 123706 182 124094 270
rect 124266 182 124654 270
rect 124826 182 125214 270
rect 125386 182 125774 270
rect 125946 182 126334 270
rect 126506 182 126894 270
rect 127066 182 127454 270
rect 127626 182 128014 270
rect 128186 182 128574 270
rect 128746 182 129134 270
rect 129306 182 129694 270
rect 129866 182 130254 270
rect 130426 182 130814 270
rect 130986 182 131374 270
rect 131546 182 131934 270
rect 132106 182 132494 270
rect 132666 182 133054 270
rect 133226 182 133614 270
rect 133786 182 134174 270
rect 134346 182 134734 270
rect 134906 182 135294 270
rect 135466 182 135854 270
rect 136026 182 136414 270
rect 136586 182 136974 270
rect 137146 182 137534 270
rect 137706 182 138094 270
rect 138266 182 138654 270
rect 138826 182 139214 270
rect 139386 182 139774 270
rect 139946 182 140334 270
rect 140506 182 140894 270
rect 141066 182 141454 270
rect 141626 182 142014 270
rect 142186 182 142574 270
rect 142746 182 143134 270
rect 143306 182 143694 270
rect 143866 182 144254 270
rect 144426 182 144814 270
rect 144986 182 145374 270
rect 145546 182 145934 270
rect 146106 182 146494 270
rect 146666 182 147054 270
rect 147226 182 147614 270
rect 147786 182 148174 270
rect 148346 182 148734 270
rect 148906 182 149294 270
rect 149466 182 149854 270
rect 150026 182 150414 270
rect 150586 182 150974 270
rect 151146 182 151534 270
rect 151706 182 152094 270
rect 152266 182 152654 270
rect 152826 182 153214 270
rect 153386 182 153774 270
rect 153946 182 154334 270
rect 154506 182 154894 270
rect 155066 182 155454 270
rect 155626 182 156014 270
rect 156186 182 156574 270
rect 156746 182 157134 270
rect 157306 182 157694 270
rect 157866 182 158254 270
rect 158426 182 158814 270
rect 158986 182 159374 270
rect 159546 182 159934 270
rect 160106 182 160494 270
rect 160666 182 161054 270
rect 161226 182 161614 270
rect 161786 182 162174 270
rect 162346 182 162734 270
rect 162906 182 163294 270
rect 163466 182 163854 270
rect 164026 182 164414 270
rect 164586 182 164974 270
rect 165146 182 165534 270
rect 165706 182 166094 270
rect 166266 182 166654 270
rect 166826 182 167214 270
rect 167386 182 167774 270
rect 167946 182 168334 270
rect 168506 182 168894 270
rect 169066 182 169454 270
rect 169626 182 170014 270
rect 170186 182 170574 270
rect 170746 182 171134 270
rect 171306 182 171694 270
rect 171866 182 172254 270
rect 172426 182 172814 270
rect 172986 182 173374 270
rect 173546 182 173934 270
rect 174106 182 174494 270
rect 174666 182 175054 270
rect 175226 182 175614 270
rect 175786 182 176174 270
rect 176346 182 176734 270
rect 176906 182 177294 270
rect 177466 182 177854 270
rect 178026 182 178414 270
rect 178586 182 178974 270
rect 179146 182 179534 270
rect 179706 182 180094 270
rect 180266 182 180654 270
rect 180826 182 181214 270
rect 181386 182 181774 270
rect 181946 182 182334 270
rect 182506 182 182894 270
rect 183066 182 183454 270
rect 183626 182 184014 270
rect 184186 182 184574 270
rect 184746 182 185134 270
rect 185306 182 185694 270
rect 185866 182 186254 270
rect 186426 182 186814 270
rect 186986 182 187374 270
rect 187546 182 187934 270
rect 188106 182 188494 270
rect 188666 182 189054 270
rect 189226 182 189614 270
rect 189786 182 190174 270
rect 190346 182 190734 270
rect 190906 182 191294 270
rect 191466 182 191854 270
rect 192026 182 192414 270
rect 192586 182 192974 270
rect 193146 182 193534 270
rect 193706 182 194094 270
rect 194266 182 194654 270
rect 194826 182 195214 270
rect 195386 182 195774 270
rect 195946 182 196334 270
rect 196506 182 196894 270
rect 197066 182 197454 270
rect 197626 182 198014 270
rect 198186 182 198574 270
rect 198746 182 199134 270
rect 199306 182 199694 270
rect 199866 182 200254 270
rect 200426 182 200814 270
rect 200986 182 201374 270
rect 201546 182 201934 270
rect 202106 182 202494 270
rect 202666 182 203054 270
rect 203226 182 203614 270
rect 203786 182 204174 270
rect 204346 182 204734 270
rect 204906 182 205294 270
rect 205466 182 205854 270
rect 206026 182 206414 270
rect 206586 182 206974 270
rect 207146 182 207534 270
rect 207706 182 208094 270
rect 208266 182 208654 270
rect 208826 182 209214 270
rect 209386 182 209774 270
rect 209946 182 210334 270
rect 210506 182 210894 270
rect 211066 182 211454 270
rect 211626 182 212014 270
rect 212186 182 212574 270
rect 212746 182 213134 270
rect 213306 182 213694 270
rect 213866 182 214254 270
rect 214426 182 214814 270
rect 214986 182 215374 270
rect 215546 182 215934 270
rect 216106 182 216494 270
rect 216666 182 217054 270
rect 217226 182 217614 270
rect 217786 182 218174 270
rect 218346 182 218734 270
rect 218906 182 219294 270
rect 219466 182 219854 270
rect 220026 182 220414 270
rect 220586 182 220974 270
rect 221146 182 221534 270
rect 221706 182 222094 270
rect 222266 182 222654 270
rect 222826 182 223214 270
rect 223386 182 223774 270
rect 223946 182 224334 270
rect 224506 182 224894 270
rect 225066 182 225454 270
rect 225626 182 226014 270
rect 226186 182 226574 270
rect 226746 182 227134 270
rect 227306 182 227694 270
rect 227866 182 228254 270
rect 228426 182 228814 270
rect 228986 182 229374 270
rect 229546 182 229934 270
rect 230106 182 230494 270
rect 230666 182 231054 270
rect 231226 182 231614 270
rect 231786 182 232174 270
rect 232346 182 232734 270
rect 232906 182 233294 270
rect 233466 182 233854 270
rect 234026 182 234414 270
rect 234586 182 234974 270
rect 235146 182 235534 270
rect 235706 182 236094 270
rect 236266 182 236654 270
rect 236826 182 237214 270
rect 237386 182 237774 270
rect 237946 182 238334 270
rect 238506 182 238894 270
rect 239066 182 239454 270
rect 239626 182 240014 270
rect 240186 182 240574 270
rect 240746 182 241134 270
rect 241306 182 241694 270
rect 241866 182 242254 270
rect 242426 182 242814 270
rect 242986 182 243374 270
rect 243546 182 243934 270
rect 244106 182 244494 270
rect 244666 182 245054 270
rect 245226 182 245614 270
rect 245786 182 246174 270
rect 246346 182 246734 270
rect 246906 182 247294 270
rect 247466 182 247854 270
rect 248026 182 248414 270
rect 248586 182 248974 270
rect 249146 182 249534 270
rect 249706 182 250094 270
rect 250266 182 250654 270
rect 250826 182 251214 270
rect 251386 182 251774 270
rect 251946 182 252334 270
rect 252506 182 252894 270
rect 253066 182 253454 270
rect 253626 182 254014 270
rect 254186 182 254574 270
rect 254746 182 255134 270
rect 255306 182 255694 270
rect 255866 182 256254 270
rect 256426 182 256814 270
rect 256986 182 257374 270
rect 257546 182 257934 270
rect 258106 182 258494 270
rect 258666 182 259054 270
rect 259226 182 259614 270
rect 259786 182 260174 270
rect 260346 182 260734 270
rect 260906 182 261294 270
rect 261466 182 261854 270
rect 262026 182 262414 270
rect 262586 182 262974 270
rect 263146 182 263534 270
rect 263706 182 264094 270
rect 264266 182 264654 270
rect 264826 182 265214 270
rect 265386 182 265774 270
rect 265946 182 266334 270
rect 266506 182 266894 270
rect 267066 182 267454 270
rect 267626 182 268014 270
rect 268186 182 268574 270
rect 268746 182 269134 270
rect 269306 182 269694 270
rect 269866 182 270254 270
rect 270426 182 270814 270
rect 270986 182 271374 270
rect 271546 182 271934 270
rect 272106 182 272494 270
rect 272666 182 273054 270
rect 273226 182 273614 270
rect 273786 182 274174 270
rect 274346 182 274734 270
rect 274906 182 275294 270
rect 275466 182 275854 270
rect 276026 182 276414 270
rect 276586 182 276974 270
rect 277146 182 277534 270
rect 277706 182 278094 270
rect 278266 182 278654 270
rect 278826 182 279214 270
rect 279386 182 279774 270
rect 279946 182 280334 270
rect 280506 182 280894 270
rect 281066 182 281454 270
rect 281626 182 282014 270
rect 282186 182 282574 270
rect 282746 182 283134 270
rect 283306 182 283694 270
rect 283866 182 284254 270
rect 284426 182 284814 270
rect 284986 182 285374 270
rect 285546 182 285934 270
rect 286106 182 295050 270
<< metal3 >>
rect 295780 292068 296500 292180
rect -480 291900 240 292012
rect -480 286468 240 286580
rect 295780 286524 296500 286636
rect -480 281036 240 281148
rect 295780 280980 296500 281092
rect -480 275604 240 275716
rect 295780 275436 296500 275548
rect -480 270172 240 270284
rect 295780 269892 296500 270004
rect -480 264740 240 264852
rect 295780 264348 296500 264460
rect -480 259308 240 259420
rect 295780 258804 296500 258916
rect -480 253876 240 253988
rect 295780 253260 296500 253372
rect -480 248444 240 248556
rect 295780 247716 296500 247828
rect -480 243012 240 243124
rect 295780 242172 296500 242284
rect -480 237580 240 237692
rect 295780 236628 296500 236740
rect -480 232148 240 232260
rect 295780 231084 296500 231196
rect -480 226716 240 226828
rect 295780 225540 296500 225652
rect -480 221284 240 221396
rect 295780 219996 296500 220108
rect -480 215852 240 215964
rect 295780 214452 296500 214564
rect -480 210420 240 210532
rect 295780 208908 296500 209020
rect -480 204988 240 205100
rect 295780 203364 296500 203476
rect -480 199556 240 199668
rect 295780 197820 296500 197932
rect -480 194124 240 194236
rect 295780 192276 296500 192388
rect -480 188692 240 188804
rect 295780 186732 296500 186844
rect -480 183260 240 183372
rect 295780 181188 296500 181300
rect -480 177828 240 177940
rect 295780 175644 296500 175756
rect -480 172396 240 172508
rect 295780 170100 296500 170212
rect -480 166964 240 167076
rect 295780 164556 296500 164668
rect -480 161532 240 161644
rect 295780 159012 296500 159124
rect -480 156100 240 156212
rect 295780 153468 296500 153580
rect -480 150668 240 150780
rect 295780 147924 296500 148036
rect -480 145236 240 145348
rect 295780 142380 296500 142492
rect -480 139804 240 139916
rect 295780 136836 296500 136948
rect -480 134372 240 134484
rect 295780 131292 296500 131404
rect -480 128940 240 129052
rect 295780 125748 296500 125860
rect -480 123508 240 123620
rect 295780 120204 296500 120316
rect -480 118076 240 118188
rect 295780 114660 296500 114772
rect -480 112644 240 112756
rect 295780 109116 296500 109228
rect -480 107212 240 107324
rect 295780 103572 296500 103684
rect -480 101780 240 101892
rect 295780 98028 296500 98140
rect -480 96348 240 96460
rect 295780 92484 296500 92596
rect -480 90916 240 91028
rect 295780 86940 296500 87052
rect -480 85484 240 85596
rect 295780 81396 296500 81508
rect -480 80052 240 80164
rect 295780 75852 296500 75964
rect -480 74620 240 74732
rect 295780 70308 296500 70420
rect -480 69188 240 69300
rect 295780 64764 296500 64876
rect -480 63756 240 63868
rect 295780 59220 296500 59332
rect -480 58324 240 58436
rect 295780 53676 296500 53788
rect -480 52892 240 53004
rect 295780 48132 296500 48244
rect -480 47460 240 47572
rect 295780 42588 296500 42700
rect -480 42028 240 42140
rect 295780 37044 296500 37156
rect -480 36596 240 36708
rect 295780 31500 296500 31612
rect -480 31164 240 31276
rect 295780 25956 296500 26068
rect -480 25732 240 25844
rect -480 20300 240 20412
rect 295780 20412 296500 20524
rect -480 14868 240 14980
rect 295780 14868 296500 14980
rect -480 9436 240 9548
rect 295780 9324 296500 9436
rect -480 4004 240 4116
rect 295780 3780 296500 3892
<< obsm3 >>
rect 9 292210 295834 293986
rect 9 292042 295750 292210
rect 270 292038 295750 292042
rect 270 291870 295834 292038
rect 9 286666 295834 291870
rect 9 286610 295750 286666
rect 270 286494 295750 286610
rect 270 286438 295834 286494
rect 9 281178 295834 286438
rect 270 281122 295834 281178
rect 270 281006 295750 281122
rect 9 280950 295750 281006
rect 9 275746 295834 280950
rect 270 275578 295834 275746
rect 270 275574 295750 275578
rect 9 275406 295750 275574
rect 9 270314 295834 275406
rect 270 270142 295834 270314
rect 9 270034 295834 270142
rect 9 269862 295750 270034
rect 9 264882 295834 269862
rect 270 264710 295834 264882
rect 9 264490 295834 264710
rect 9 264318 295750 264490
rect 9 259450 295834 264318
rect 270 259278 295834 259450
rect 9 258946 295834 259278
rect 9 258774 295750 258946
rect 9 254018 295834 258774
rect 270 253846 295834 254018
rect 9 253402 295834 253846
rect 9 253230 295750 253402
rect 9 248586 295834 253230
rect 270 248414 295834 248586
rect 9 247858 295834 248414
rect 9 247686 295750 247858
rect 9 243154 295834 247686
rect 270 242982 295834 243154
rect 9 242314 295834 242982
rect 9 242142 295750 242314
rect 9 237722 295834 242142
rect 270 237550 295834 237722
rect 9 236770 295834 237550
rect 9 236598 295750 236770
rect 9 232290 295834 236598
rect 270 232118 295834 232290
rect 9 231226 295834 232118
rect 9 231054 295750 231226
rect 9 226858 295834 231054
rect 270 226686 295834 226858
rect 9 225682 295834 226686
rect 9 225510 295750 225682
rect 9 221426 295834 225510
rect 270 221254 295834 221426
rect 9 220138 295834 221254
rect 9 219966 295750 220138
rect 9 215994 295834 219966
rect 270 215822 295834 215994
rect 9 214594 295834 215822
rect 9 214422 295750 214594
rect 9 210562 295834 214422
rect 270 210390 295834 210562
rect 9 209050 295834 210390
rect 9 208878 295750 209050
rect 9 205130 295834 208878
rect 270 204958 295834 205130
rect 9 203506 295834 204958
rect 9 203334 295750 203506
rect 9 199698 295834 203334
rect 270 199526 295834 199698
rect 9 197962 295834 199526
rect 9 197790 295750 197962
rect 9 194266 295834 197790
rect 270 194094 295834 194266
rect 9 192418 295834 194094
rect 9 192246 295750 192418
rect 9 188834 295834 192246
rect 270 188662 295834 188834
rect 9 186874 295834 188662
rect 9 186702 295750 186874
rect 9 183402 295834 186702
rect 270 183230 295834 183402
rect 9 181330 295834 183230
rect 9 181158 295750 181330
rect 9 177970 295834 181158
rect 270 177798 295834 177970
rect 9 175786 295834 177798
rect 9 175614 295750 175786
rect 9 172538 295834 175614
rect 270 172366 295834 172538
rect 9 170242 295834 172366
rect 9 170070 295750 170242
rect 9 167106 295834 170070
rect 270 166934 295834 167106
rect 9 164698 295834 166934
rect 9 164526 295750 164698
rect 9 161674 295834 164526
rect 270 161502 295834 161674
rect 9 159154 295834 161502
rect 9 158982 295750 159154
rect 9 156242 295834 158982
rect 270 156070 295834 156242
rect 9 153610 295834 156070
rect 9 153438 295750 153610
rect 9 150810 295834 153438
rect 270 150638 295834 150810
rect 9 148066 295834 150638
rect 9 147894 295750 148066
rect 9 145378 295834 147894
rect 270 145206 295834 145378
rect 9 142522 295834 145206
rect 9 142350 295750 142522
rect 9 139946 295834 142350
rect 270 139774 295834 139946
rect 9 136978 295834 139774
rect 9 136806 295750 136978
rect 9 134514 295834 136806
rect 270 134342 295834 134514
rect 9 131434 295834 134342
rect 9 131262 295750 131434
rect 9 129082 295834 131262
rect 270 128910 295834 129082
rect 9 125890 295834 128910
rect 9 125718 295750 125890
rect 9 123650 295834 125718
rect 270 123478 295834 123650
rect 9 120346 295834 123478
rect 9 120174 295750 120346
rect 9 118218 295834 120174
rect 270 118046 295834 118218
rect 9 114802 295834 118046
rect 9 114630 295750 114802
rect 9 112786 295834 114630
rect 270 112614 295834 112786
rect 9 109258 295834 112614
rect 9 109086 295750 109258
rect 9 107354 295834 109086
rect 270 107182 295834 107354
rect 9 103714 295834 107182
rect 9 103542 295750 103714
rect 9 101922 295834 103542
rect 270 101750 295834 101922
rect 9 98170 295834 101750
rect 9 97998 295750 98170
rect 9 96490 295834 97998
rect 270 96318 295834 96490
rect 9 92626 295834 96318
rect 9 92454 295750 92626
rect 9 91058 295834 92454
rect 270 90886 295834 91058
rect 9 87082 295834 90886
rect 9 86910 295750 87082
rect 9 85626 295834 86910
rect 270 85454 295834 85626
rect 9 81538 295834 85454
rect 9 81366 295750 81538
rect 9 80194 295834 81366
rect 270 80022 295834 80194
rect 9 75994 295834 80022
rect 9 75822 295750 75994
rect 9 74762 295834 75822
rect 270 74590 295834 74762
rect 9 70450 295834 74590
rect 9 70278 295750 70450
rect 9 69330 295834 70278
rect 270 69158 295834 69330
rect 9 64906 295834 69158
rect 9 64734 295750 64906
rect 9 63898 295834 64734
rect 270 63726 295834 63898
rect 9 59362 295834 63726
rect 9 59190 295750 59362
rect 9 58466 295834 59190
rect 270 58294 295834 58466
rect 9 53818 295834 58294
rect 9 53646 295750 53818
rect 9 53034 295834 53646
rect 270 52862 295834 53034
rect 9 48274 295834 52862
rect 9 48102 295750 48274
rect 9 47602 295834 48102
rect 270 47430 295834 47602
rect 9 42730 295834 47430
rect 9 42558 295750 42730
rect 9 42170 295834 42558
rect 270 41998 295834 42170
rect 9 37186 295834 41998
rect 9 37014 295750 37186
rect 9 36738 295834 37014
rect 270 36566 295834 36738
rect 9 31642 295834 36566
rect 9 31470 295750 31642
rect 9 31306 295834 31470
rect 270 31134 295834 31306
rect 9 26098 295834 31134
rect 9 25926 295750 26098
rect 9 25874 295834 25926
rect 270 25702 295834 25874
rect 9 20554 295834 25702
rect 9 20442 295750 20554
rect 270 20382 295750 20442
rect 270 20270 295834 20382
rect 9 15010 295834 20270
rect 270 14838 295750 15010
rect 9 9578 295834 14838
rect 270 9466 295834 9578
rect 270 9406 295750 9466
rect 9 9294 295750 9406
rect 9 4146 295834 9294
rect 270 3974 295834 4146
rect 9 3922 295834 3974
rect 9 3750 295750 3922
rect 9 350 295834 3750
<< metal4 >>
rect -958 -822 -648 299134
rect -478 -342 -168 298654
rect 1577 -822 1887 299134
rect 3437 -822 3747 299134
rect 10577 229171 10887 299134
rect 12437 229171 12747 299134
rect 19577 229171 19887 299134
rect 21437 229171 21747 299134
rect 28577 229171 28887 299134
rect 30437 229171 30747 299134
rect 37577 229171 37887 299134
rect 39437 229171 39747 299134
rect 46577 229171 46887 299134
rect 48437 229171 48747 299134
rect 55577 229171 55887 299134
rect 57437 229171 57747 299134
rect 64577 229171 64887 299134
rect 66437 229171 66747 299134
rect 73577 229171 73887 299134
rect 75437 229171 75747 299134
rect 82577 229171 82887 299134
rect 84437 229171 84747 299134
rect 91577 229171 91887 299134
rect 93437 229171 93747 299134
rect 12437 149171 12747 159429
rect 21437 149171 21747 159429
rect 30437 149171 30747 159429
rect 39437 149171 39747 159429
rect 48437 149171 48747 159429
rect 57437 149171 57747 159429
rect 66437 149171 66747 159429
rect 75437 149171 75747 159429
rect 84437 149171 84747 159429
rect 93437 149171 93747 159429
rect 10577 -822 10887 79429
rect 12437 -822 12747 79429
rect 19577 -822 19887 79429
rect 21437 -822 21747 79429
rect 28577 55619 28887 79429
rect 30437 55619 30747 79429
rect 37577 55619 37887 79429
rect 39437 55619 39747 79429
rect 46577 55619 46887 79429
rect 48437 55619 48747 79429
rect 55577 55619 55887 79429
rect 57437 55619 57747 79429
rect 64577 55619 64887 79429
rect 66437 55619 66747 79429
rect 73577 55619 73887 79429
rect 75437 55619 75747 79429
rect 82577 55619 82887 79429
rect 84437 55619 84747 79429
rect 28577 -822 28887 38797
rect 30437 -822 30747 38797
rect 37577 -822 37887 38797
rect 39437 -822 39747 38797
rect 46577 -822 46887 38797
rect 48437 -822 48747 38797
rect 55577 -822 55887 38797
rect 57437 -822 57747 38797
rect 64577 -822 64887 38797
rect 66437 -822 66747 38797
rect 73577 -822 73887 38797
rect 75437 -822 75747 38797
rect 82577 -822 82887 38797
rect 84437 -822 84747 38797
rect 91577 -822 91887 79429
rect 93437 -822 93747 79429
rect 100577 -822 100887 299134
rect 102437 -822 102747 299134
rect 109577 229171 109887 299134
rect 111437 229171 111747 299134
rect 118577 229171 118887 299134
rect 120437 229171 120747 299134
rect 127577 229171 127887 299134
rect 129437 229171 129747 299134
rect 136577 229171 136887 299134
rect 138437 229171 138747 299134
rect 145577 229171 145887 299134
rect 147437 229171 147747 299134
rect 154577 229171 154887 299134
rect 156437 229171 156747 299134
rect 163577 229171 163887 299134
rect 165437 229171 165747 299134
rect 172577 229171 172887 299134
rect 174437 229171 174747 299134
rect 181577 229171 181887 299134
rect 183437 229171 183747 299134
rect 111437 149171 111747 159429
rect 120437 149171 120747 159429
rect 129437 149171 129747 159429
rect 138437 149171 138747 159429
rect 147437 149171 147747 159429
rect 156437 149171 156747 159429
rect 165437 149171 165747 159429
rect 174437 149171 174747 159429
rect 183437 149171 183747 159429
rect 109577 74171 109887 79429
rect 111437 74171 111747 79429
rect 118577 74171 118887 79429
rect 120437 74171 120747 79429
rect 127577 74171 127887 79429
rect 129437 74171 129747 79429
rect 136577 74171 136887 79429
rect 138437 74171 138747 79429
rect 145577 74171 145887 79429
rect 147437 74171 147747 79429
rect 154577 74171 154887 79429
rect 156437 74171 156747 79429
rect 163577 74171 163887 79429
rect 165437 74171 165747 79429
rect 172577 74171 172887 79429
rect 174437 74171 174747 79429
rect 181577 74171 181887 79429
rect 183437 74171 183747 79429
rect 109577 -822 109887 4429
rect 118577 -822 118887 4429
rect 127577 -822 127887 4429
rect 136577 -822 136887 4429
rect 145577 -822 145887 4429
rect 154577 -822 154887 4429
rect 163577 -822 163887 4429
rect 172577 -822 172887 4429
rect 181577 -822 181887 4429
rect 190577 -822 190887 299134
rect 192437 -822 192747 299134
rect 199577 -822 199887 299134
rect 201437 -822 201747 299134
rect 208577 229171 208887 299134
rect 210437 229171 210747 299134
rect 217577 229171 217887 299134
rect 219437 229171 219747 299134
rect 226577 229171 226887 299134
rect 228437 229171 228747 299134
rect 235577 229171 235887 299134
rect 237437 229171 237747 299134
rect 244577 229171 244887 299134
rect 246437 229171 246747 299134
rect 253577 229171 253887 299134
rect 255437 229171 255747 299134
rect 262577 229171 262887 299134
rect 264437 229171 264747 299134
rect 271577 229171 271887 299134
rect 273437 229171 273747 299134
rect 280577 229171 280887 299134
rect 282437 229171 282747 299134
rect 210437 149171 210747 159429
rect 219437 149171 219747 159429
rect 228437 149171 228747 159429
rect 237437 149171 237747 159429
rect 246437 149171 246747 159429
rect 255437 149171 255747 159429
rect 264437 149171 264747 159429
rect 273437 149171 273747 159429
rect 282437 149171 282747 159429
rect 208577 -822 208887 79429
rect 210437 -822 210747 79429
rect 217577 -822 217887 79429
rect 219437 -822 219747 79429
rect 226577 -822 226887 79429
rect 228437 -822 228747 79429
rect 235577 -822 235887 79429
rect 237437 -822 237747 79429
rect 244577 -822 244887 79429
rect 246437 -822 246747 79429
rect 253577 -822 253887 79429
rect 255437 -822 255747 79429
rect 262577 -822 262887 79429
rect 264437 -822 264747 79429
rect 271577 -822 271887 79429
rect 273437 -822 273747 79429
rect 280577 -822 280887 79429
rect 282437 -822 282747 79429
rect 289577 -822 289887 299134
rect 291437 -822 291747 299134
rect 298200 -342 298510 298654
rect 298680 -822 298990 299134
<< obsm4 >>
rect 3822 229141 10547 293991
rect 10917 229141 12407 293991
rect 12777 229141 19547 293991
rect 19917 229141 21407 293991
rect 21777 229141 28547 293991
rect 28917 229141 30407 293991
rect 30777 229141 37547 293991
rect 37917 229141 39407 293991
rect 39777 229141 46547 293991
rect 46917 229141 48407 293991
rect 48777 229141 55547 293991
rect 55917 229141 57407 293991
rect 57777 229141 64547 293991
rect 64917 229141 66407 293991
rect 66777 229141 73547 293991
rect 73917 229141 75407 293991
rect 75777 229141 82547 293991
rect 82917 229141 84407 293991
rect 84777 229141 91547 293991
rect 91917 229141 93407 293991
rect 93777 229141 100547 293991
rect 3822 159459 100547 229141
rect 3822 149141 12407 159459
rect 12777 149141 21407 159459
rect 21777 149141 30407 159459
rect 30777 149141 39407 159459
rect 39777 149141 48407 159459
rect 48777 149141 57407 159459
rect 57777 149141 66407 159459
rect 66777 149141 75407 159459
rect 75777 149141 84407 159459
rect 84777 149141 93407 159459
rect 93777 149141 100547 159459
rect 3822 79459 100547 149141
rect 3822 345 10547 79459
rect 10917 345 12407 79459
rect 12777 345 19547 79459
rect 19917 345 21407 79459
rect 21777 55589 28547 79459
rect 28917 55589 30407 79459
rect 30777 55589 37547 79459
rect 37917 55589 39407 79459
rect 39777 55589 46547 79459
rect 46917 55589 48407 79459
rect 48777 55589 55547 79459
rect 55917 55589 57407 79459
rect 57777 55589 64547 79459
rect 64917 55589 66407 79459
rect 66777 55589 73547 79459
rect 73917 55589 75407 79459
rect 75777 55589 82547 79459
rect 82917 55589 84407 79459
rect 84777 55589 91547 79459
rect 21777 38827 91547 55589
rect 21777 345 28547 38827
rect 28917 345 30407 38827
rect 30777 345 37547 38827
rect 37917 345 39407 38827
rect 39777 345 46547 38827
rect 46917 345 48407 38827
rect 48777 345 55547 38827
rect 55917 345 57407 38827
rect 57777 345 64547 38827
rect 64917 345 66407 38827
rect 66777 345 73547 38827
rect 73917 345 75407 38827
rect 75777 345 82547 38827
rect 82917 345 84407 38827
rect 84777 345 91547 38827
rect 91917 345 93407 79459
rect 93777 345 100547 79459
rect 100917 345 102407 293991
rect 102777 229141 109547 293991
rect 109917 229141 111407 293991
rect 111777 229141 118547 293991
rect 118917 229141 120407 293991
rect 120777 229141 127547 293991
rect 127917 229141 129407 293991
rect 129777 229141 136547 293991
rect 136917 229141 138407 293991
rect 138777 229141 145547 293991
rect 145917 229141 147407 293991
rect 147777 229141 154547 293991
rect 154917 229141 156407 293991
rect 156777 229141 163547 293991
rect 163917 229141 165407 293991
rect 165777 229141 172547 293991
rect 172917 229141 174407 293991
rect 174777 229141 181547 293991
rect 181917 229141 183407 293991
rect 183777 229141 190547 293991
rect 102777 159459 190547 229141
rect 102777 149141 111407 159459
rect 111777 149141 120407 159459
rect 120777 149141 129407 159459
rect 129777 149141 138407 159459
rect 138777 149141 147407 159459
rect 147777 149141 156407 159459
rect 156777 149141 165407 159459
rect 165777 149141 174407 159459
rect 174777 149141 183407 159459
rect 183777 149141 190547 159459
rect 102777 79459 190547 149141
rect 102777 74141 109547 79459
rect 109917 74141 111407 79459
rect 111777 74141 118547 79459
rect 118917 74141 120407 79459
rect 120777 74141 127547 79459
rect 127917 74141 129407 79459
rect 129777 74141 136547 79459
rect 136917 74141 138407 79459
rect 138777 74141 145547 79459
rect 145917 74141 147407 79459
rect 147777 74141 154547 79459
rect 154917 74141 156407 79459
rect 156777 74141 163547 79459
rect 163917 74141 165407 79459
rect 165777 74141 172547 79459
rect 172917 74141 174407 79459
rect 174777 74141 181547 79459
rect 181917 74141 183407 79459
rect 183777 74141 190547 79459
rect 102777 4459 190547 74141
rect 102777 345 109547 4459
rect 109917 345 118547 4459
rect 118917 345 127547 4459
rect 127917 345 136547 4459
rect 136917 345 145547 4459
rect 145917 345 154547 4459
rect 154917 345 163547 4459
rect 163917 345 172547 4459
rect 172917 345 181547 4459
rect 181917 345 190547 4459
rect 190917 345 192407 293991
rect 192777 345 199547 293991
rect 199917 345 201407 293991
rect 201777 229141 208547 293991
rect 208917 229141 210407 293991
rect 210777 229141 217547 293991
rect 217917 229141 219407 293991
rect 219777 229141 226547 293991
rect 226917 229141 228407 293991
rect 228777 229141 235547 293991
rect 235917 229141 237407 293991
rect 237777 229141 244547 293991
rect 244917 229141 246407 293991
rect 246777 229141 253547 293991
rect 253917 229141 255407 293991
rect 255777 229141 262547 293991
rect 262917 229141 264407 293991
rect 264777 229141 271547 293991
rect 271917 229141 273407 293991
rect 273777 229141 280547 293991
rect 280917 229141 282407 293991
rect 282777 229141 287966 293991
rect 201777 159459 287966 229141
rect 201777 149141 210407 159459
rect 210777 149141 219407 159459
rect 219777 149141 228407 159459
rect 228777 149141 237407 159459
rect 237777 149141 246407 159459
rect 246777 149141 255407 159459
rect 255777 149141 264407 159459
rect 264777 149141 273407 159459
rect 273777 149141 282407 159459
rect 282777 149141 287966 159459
rect 201777 79459 287966 149141
rect 201777 345 208547 79459
rect 208917 345 210407 79459
rect 210777 345 217547 79459
rect 217917 345 219407 79459
rect 219777 345 226547 79459
rect 226917 345 228407 79459
rect 228777 345 235547 79459
rect 235917 345 237407 79459
rect 237777 345 244547 79459
rect 244917 345 246407 79459
rect 246777 345 253547 79459
rect 253917 345 255407 79459
rect 255777 345 262547 79459
rect 262917 345 264407 79459
rect 264777 345 271547 79459
rect 271917 345 273407 79459
rect 273777 345 280547 79459
rect 280917 345 282407 79459
rect 282777 345 287966 79459
<< metal5 >>
rect -958 298824 298990 299134
rect -478 298344 298510 298654
rect -958 292913 298990 293223
rect -958 289913 298990 290223
rect -958 283913 298990 284223
rect -958 280913 298990 281223
rect -958 274913 298990 275223
rect -958 271913 298990 272223
rect -958 265913 298990 266223
rect -958 262913 298990 263223
rect -958 256913 298990 257223
rect -958 253913 298990 254223
rect -958 247913 298990 248223
rect -958 244913 298990 245223
rect -958 238913 298990 239223
rect -958 235913 298990 236223
rect -958 229913 298990 230223
rect -958 226913 298990 227223
rect -958 220913 298990 221223
rect -958 217913 298990 218223
rect -958 211913 298990 212223
rect -958 208913 298990 209223
rect -958 202913 298990 203223
rect -958 199913 298990 200223
rect -958 193913 298990 194223
rect -958 190913 298990 191223
rect -958 184913 298990 185223
rect -958 181913 298990 182223
rect -958 175913 298990 176223
rect -958 172913 298990 173223
rect -958 166913 298990 167223
rect -958 163913 298990 164223
rect -958 157913 298990 158223
rect -958 154913 298990 155223
rect -958 148913 298990 149223
rect -958 145913 298990 146223
rect -958 139913 298990 140223
rect -958 136913 298990 137223
rect -958 130913 298990 131223
rect -958 127913 298990 128223
rect -958 121913 298990 122223
rect -958 118913 298990 119223
rect -958 112913 298990 113223
rect -958 109913 298990 110223
rect -958 103913 298990 104223
rect -958 100913 298990 101223
rect -958 94913 298990 95223
rect -958 91913 298990 92223
rect -958 85913 298990 86223
rect -958 82913 298990 83223
rect -958 76913 298990 77223
rect -958 73913 298990 74223
rect -958 67913 298990 68223
rect -958 64913 298990 65223
rect -958 58913 298990 59223
rect -958 55913 298990 56223
rect -958 49913 298990 50223
rect -958 46913 298990 47223
rect -958 40913 298990 41223
rect -958 37913 298990 38223
rect -958 31913 298990 32223
rect -958 28913 298990 29223
rect -958 22913 298990 23223
rect -958 19913 298990 20223
rect -958 13913 298990 14223
rect -958 10913 298990 11223
rect -958 4913 298990 5223
rect -958 1913 298990 2223
rect -478 -342 298510 -32
rect -958 -822 298990 -512
<< labels >>
rlabel metal3 s 295780 120204 296500 120316 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 225596 295780 225708 296500 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 192892 295780 193004 296500 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 160188 295780 160300 296500 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 127484 295780 127596 296500 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 94780 295780 94892 296500 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 62076 295780 62188 296500 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 29372 295780 29484 296500 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s -480 291900 240 292012 4 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s -480 270172 240 270284 4 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s -480 248444 240 248556 4 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 295780 142380 296500 142492 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s -480 226716 240 226828 4 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s -480 204988 240 205100 4 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s -480 183260 240 183372 4 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s -480 161532 240 161644 4 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s -480 139804 240 139916 4 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s -480 118076 240 118188 4 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s -480 96348 240 96460 4 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s -480 74620 240 74732 4 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s -480 52892 240 53004 4 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 295780 164556 296500 164668 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 295780 186732 296500 186844 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 295780 208908 296500 209020 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 295780 231084 296500 231196 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 295780 253260 296500 253372 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 295780 275436 296500 275548 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 291004 295780 291116 296500 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 258300 295780 258412 296500 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 295780 3780 296500 3892 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 295780 192276 296500 192388 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 295780 214452 296500 214564 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 295780 236628 296500 236740 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 295780 258804 296500 258916 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 295780 280980 296500 281092 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 282828 295780 282940 296500 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 250124 295780 250236 296500 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 217420 295780 217532 296500 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 184716 295780 184828 296500 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 152012 295780 152124 296500 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 295780 20412 296500 20524 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 119308 295780 119420 296500 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 86604 295780 86716 296500 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 53900 295780 54012 296500 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 21196 295780 21308 296500 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s -480 286468 240 286580 4 io_in[24]
port 46 nsew signal input
rlabel metal3 s -480 264740 240 264852 4 io_in[25]
port 47 nsew signal input
rlabel metal3 s -480 243012 240 243124 4 io_in[26]
port 48 nsew signal input
rlabel metal3 s -480 221284 240 221396 4 io_in[27]
port 49 nsew signal input
rlabel metal3 s -480 199556 240 199668 4 io_in[28]
port 50 nsew signal input
rlabel metal3 s -480 177828 240 177940 4 io_in[29]
port 51 nsew signal input
rlabel metal3 s 295780 37044 296500 37156 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s -480 156100 240 156212 4 io_in[30]
port 53 nsew signal input
rlabel metal3 s -480 134372 240 134484 4 io_in[31]
port 54 nsew signal input
rlabel metal3 s -480 112644 240 112756 4 io_in[32]
port 55 nsew signal input
rlabel metal3 s -480 90916 240 91028 4 io_in[33]
port 56 nsew signal input
rlabel metal3 s -480 69188 240 69300 4 io_in[34]
port 57 nsew signal input
rlabel metal3 s -480 47460 240 47572 4 io_in[35]
port 58 nsew signal input
rlabel metal3 s -480 31164 240 31276 4 io_in[36]
port 59 nsew signal input
rlabel metal3 s -480 14868 240 14980 4 io_in[37]
port 60 nsew signal input
rlabel metal3 s 295780 53676 296500 53788 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 295780 70308 296500 70420 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 295780 86940 296500 87052 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 295780 103572 296500 103684 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 295780 125748 296500 125860 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 295780 147924 296500 148036 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 295780 170100 296500 170212 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 295780 14868 296500 14980 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 295780 203364 296500 203476 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 295780 225540 296500 225652 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 295780 247716 296500 247828 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 295780 269892 296500 270004 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 295780 292068 296500 292180 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 266476 295780 266588 296500 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 233772 295780 233884 296500 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 201068 295780 201180 296500 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 168364 295780 168476 296500 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 135660 295780 135772 296500 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 295780 31500 296500 31612 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 102956 295780 103068 296500 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 70252 295780 70364 296500 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 37548 295780 37660 296500 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 4844 295780 4956 296500 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s -480 275604 240 275716 4 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s -480 253876 240 253988 4 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s -480 232148 240 232260 4 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s -480 210420 240 210532 4 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s -480 188692 240 188804 4 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s -480 166964 240 167076 4 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 295780 48132 296500 48244 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s -480 145236 240 145348 4 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s -480 123508 240 123620 4 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s -480 101780 240 101892 4 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s -480 80052 240 80164 4 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s -480 58324 240 58436 4 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s -480 36596 240 36708 4 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s -480 20300 240 20412 4 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s -480 4004 240 4116 4 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 295780 64764 296500 64876 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 295780 81396 296500 81508 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 295780 98028 296500 98140 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 295780 114660 296500 114772 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 295780 136836 296500 136948 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 295780 159012 296500 159124 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 295780 181188 296500 181300 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 295780 9324 296500 9436 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 295780 197820 296500 197932 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 295780 219996 296500 220108 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 295780 242172 296500 242284 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 295780 264348 296500 264460 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 295780 286524 296500 286636 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 274652 295780 274764 296500 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 241948 295780 242060 296500 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 209244 295780 209356 296500 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 176540 295780 176652 296500 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 143836 295780 143948 296500 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 295780 25956 296500 26068 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 111132 295780 111244 296500 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 78428 295780 78540 296500 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 45724 295780 45836 296500 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 13020 295780 13132 296500 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s -480 281036 240 281148 4 io_out[24]
port 122 nsew signal output
rlabel metal3 s -480 259308 240 259420 4 io_out[25]
port 123 nsew signal output
rlabel metal3 s -480 237580 240 237692 4 io_out[26]
port 124 nsew signal output
rlabel metal3 s -480 215852 240 215964 4 io_out[27]
port 125 nsew signal output
rlabel metal3 s -480 194124 240 194236 4 io_out[28]
port 126 nsew signal output
rlabel metal3 s -480 172396 240 172508 4 io_out[29]
port 127 nsew signal output
rlabel metal3 s 295780 42588 296500 42700 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s -480 150668 240 150780 4 io_out[30]
port 129 nsew signal output
rlabel metal3 s -480 128940 240 129052 4 io_out[31]
port 130 nsew signal output
rlabel metal3 s -480 107212 240 107324 4 io_out[32]
port 131 nsew signal output
rlabel metal3 s -480 85484 240 85596 4 io_out[33]
port 132 nsew signal output
rlabel metal3 s -480 63756 240 63868 4 io_out[34]
port 133 nsew signal output
rlabel metal3 s -480 42028 240 42140 4 io_out[35]
port 134 nsew signal output
rlabel metal3 s -480 25732 240 25844 4 io_out[36]
port 135 nsew signal output
rlabel metal3 s -480 9436 240 9548 4 io_out[37]
port 136 nsew signal output
rlabel metal3 s 295780 59220 296500 59332 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 295780 75852 296500 75964 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 295780 92484 296500 92596 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 295780 109116 296500 109228 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 295780 131292 296500 131404 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 295780 153468 296500 153580 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 295780 175644 296500 175756 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 69244 -480 69356 240 8 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 237244 -480 237356 240 8 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 238924 -480 239036 240 8 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 240604 -480 240716 240 8 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 242284 -480 242396 240 8 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 243964 -480 244076 240 8 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 245644 -480 245756 240 8 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 247324 -480 247436 240 8 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 249004 -480 249116 240 8 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 250684 -480 250796 240 8 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 252364 -480 252476 240 8 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 86044 -480 86156 240 8 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 254044 -480 254156 240 8 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 255724 -480 255836 240 8 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 257404 -480 257516 240 8 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 259084 -480 259196 240 8 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 260764 -480 260876 240 8 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 262444 -480 262556 240 8 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 264124 -480 264236 240 8 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 265804 -480 265916 240 8 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 267484 -480 267596 240 8 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 269164 -480 269276 240 8 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 87724 -480 87836 240 8 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 270844 -480 270956 240 8 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 272524 -480 272636 240 8 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 274204 -480 274316 240 8 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 275884 -480 275996 240 8 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 277564 -480 277676 240 8 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 279244 -480 279356 240 8 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 280924 -480 281036 240 8 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 282604 -480 282716 240 8 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 89404 -480 89516 240 8 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 91084 -480 91196 240 8 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 92764 -480 92876 240 8 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 94444 -480 94556 240 8 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 96124 -480 96236 240 8 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 97804 -480 97916 240 8 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 99484 -480 99596 240 8 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 101164 -480 101276 240 8 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 70924 -480 71036 240 8 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 102844 -480 102956 240 8 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 104524 -480 104636 240 8 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 106204 -480 106316 240 8 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 107884 -480 107996 240 8 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 109564 -480 109676 240 8 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 111244 -480 111356 240 8 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 112924 -480 113036 240 8 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 114604 -480 114716 240 8 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 116284 -480 116396 240 8 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 117964 -480 118076 240 8 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 72604 -480 72716 240 8 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 119644 -480 119756 240 8 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 121324 -480 121436 240 8 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 123004 -480 123116 240 8 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 124684 -480 124796 240 8 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 126364 -480 126476 240 8 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 128044 -480 128156 240 8 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 129724 -480 129836 240 8 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 131404 -480 131516 240 8 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 133084 -480 133196 240 8 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 134764 -480 134876 240 8 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 74284 -480 74396 240 8 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 136444 -480 136556 240 8 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 138124 -480 138236 240 8 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 139804 -480 139916 240 8 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 141484 -480 141596 240 8 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 143164 -480 143276 240 8 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 144844 -480 144956 240 8 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 146524 -480 146636 240 8 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 148204 -480 148316 240 8 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 149884 -480 149996 240 8 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 151564 -480 151676 240 8 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 75964 -480 76076 240 8 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 153244 -480 153356 240 8 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 154924 -480 155036 240 8 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 156604 -480 156716 240 8 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 158284 -480 158396 240 8 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 159964 -480 160076 240 8 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 161644 -480 161756 240 8 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 163324 -480 163436 240 8 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 165004 -480 165116 240 8 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 166684 -480 166796 240 8 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 168364 -480 168476 240 8 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 77644 -480 77756 240 8 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 170044 -480 170156 240 8 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 171724 -480 171836 240 8 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 173404 -480 173516 240 8 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 175084 -480 175196 240 8 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 176764 -480 176876 240 8 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 178444 -480 178556 240 8 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 180124 -480 180236 240 8 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 181804 -480 181916 240 8 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 183484 -480 183596 240 8 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 185164 -480 185276 240 8 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 79324 -480 79436 240 8 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 186844 -480 186956 240 8 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 188524 -480 188636 240 8 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 190204 -480 190316 240 8 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 191884 -480 191996 240 8 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 193564 -480 193676 240 8 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 195244 -480 195356 240 8 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 196924 -480 197036 240 8 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 198604 -480 198716 240 8 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 200284 -480 200396 240 8 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 201964 -480 202076 240 8 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 81004 -480 81116 240 8 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 203644 -480 203756 240 8 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 205324 -480 205436 240 8 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 207004 -480 207116 240 8 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 208684 -480 208796 240 8 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 210364 -480 210476 240 8 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 212044 -480 212156 240 8 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 213724 -480 213836 240 8 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 215404 -480 215516 240 8 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 217084 -480 217196 240 8 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 218764 -480 218876 240 8 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 82684 -480 82796 240 8 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 220444 -480 220556 240 8 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 222124 -480 222236 240 8 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 223804 -480 223916 240 8 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 225484 -480 225596 240 8 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 227164 -480 227276 240 8 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 228844 -480 228956 240 8 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 230524 -480 230636 240 8 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 232204 -480 232316 240 8 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 233884 -480 233996 240 8 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 235564 -480 235676 240 8 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 84364 -480 84476 240 8 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 69804 -480 69916 240 8 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 237804 -480 237916 240 8 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 239484 -480 239596 240 8 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 241164 -480 241276 240 8 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 242844 -480 242956 240 8 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 244524 -480 244636 240 8 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 246204 -480 246316 240 8 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 247884 -480 247996 240 8 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 249564 -480 249676 240 8 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 251244 -480 251356 240 8 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 252924 -480 253036 240 8 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 86604 -480 86716 240 8 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 254604 -480 254716 240 8 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 256284 -480 256396 240 8 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 257964 -480 258076 240 8 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 259644 -480 259756 240 8 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 261324 -480 261436 240 8 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 263004 -480 263116 240 8 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 264684 -480 264796 240 8 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 266364 -480 266476 240 8 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 268044 -480 268156 240 8 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 269724 -480 269836 240 8 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 88284 -480 88396 240 8 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 271404 -480 271516 240 8 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 273084 -480 273196 240 8 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 274764 -480 274876 240 8 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 276444 -480 276556 240 8 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 278124 -480 278236 240 8 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 279804 -480 279916 240 8 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 281484 -480 281596 240 8 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 283164 -480 283276 240 8 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 89964 -480 90076 240 8 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 91644 -480 91756 240 8 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 93324 -480 93436 240 8 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 95004 -480 95116 240 8 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 96684 -480 96796 240 8 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 98364 -480 98476 240 8 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 100044 -480 100156 240 8 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 101724 -480 101836 240 8 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 71484 -480 71596 240 8 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 103404 -480 103516 240 8 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 105084 -480 105196 240 8 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 106764 -480 106876 240 8 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 108444 -480 108556 240 8 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 110124 -480 110236 240 8 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 111804 -480 111916 240 8 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 113484 -480 113596 240 8 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 115164 -480 115276 240 8 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 116844 -480 116956 240 8 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 118524 -480 118636 240 8 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 73164 -480 73276 240 8 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 120204 -480 120316 240 8 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 121884 -480 121996 240 8 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 123564 -480 123676 240 8 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 125244 -480 125356 240 8 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 126924 -480 127036 240 8 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 128604 -480 128716 240 8 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 130284 -480 130396 240 8 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 131964 -480 132076 240 8 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 133644 -480 133756 240 8 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 135324 -480 135436 240 8 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 74844 -480 74956 240 8 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 137004 -480 137116 240 8 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 138684 -480 138796 240 8 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 140364 -480 140476 240 8 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 142044 -480 142156 240 8 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 143724 -480 143836 240 8 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 145404 -480 145516 240 8 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 147084 -480 147196 240 8 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 148764 -480 148876 240 8 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 150444 -480 150556 240 8 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 152124 -480 152236 240 8 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 76524 -480 76636 240 8 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 153804 -480 153916 240 8 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 155484 -480 155596 240 8 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 157164 -480 157276 240 8 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 158844 -480 158956 240 8 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 160524 -480 160636 240 8 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 162204 -480 162316 240 8 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 163884 -480 163996 240 8 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 165564 -480 165676 240 8 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 167244 -480 167356 240 8 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 168924 -480 169036 240 8 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 78204 -480 78316 240 8 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 170604 -480 170716 240 8 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 172284 -480 172396 240 8 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 173964 -480 174076 240 8 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 175644 -480 175756 240 8 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 177324 -480 177436 240 8 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 179004 -480 179116 240 8 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 180684 -480 180796 240 8 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 182364 -480 182476 240 8 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 184044 -480 184156 240 8 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 185724 -480 185836 240 8 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 79884 -480 79996 240 8 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 187404 -480 187516 240 8 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 189084 -480 189196 240 8 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 190764 -480 190876 240 8 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 192444 -480 192556 240 8 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 194124 -480 194236 240 8 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 195804 -480 195916 240 8 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 197484 -480 197596 240 8 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 199164 -480 199276 240 8 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 200844 -480 200956 240 8 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 202524 -480 202636 240 8 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 81564 -480 81676 240 8 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 204204 -480 204316 240 8 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 205884 -480 205996 240 8 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 207564 -480 207676 240 8 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 209244 -480 209356 240 8 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 210924 -480 211036 240 8 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 212604 -480 212716 240 8 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 214284 -480 214396 240 8 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 215964 -480 216076 240 8 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 217644 -480 217756 240 8 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 219324 -480 219436 240 8 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 83244 -480 83356 240 8 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 221004 -480 221116 240 8 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 222684 -480 222796 240 8 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 224364 -480 224476 240 8 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 226044 -480 226156 240 8 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 227724 -480 227836 240 8 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 229404 -480 229516 240 8 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 231084 -480 231196 240 8 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 232764 -480 232876 240 8 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 234444 -480 234556 240 8 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 236124 -480 236236 240 8 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 84924 -480 85036 240 8 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 70364 -480 70476 240 8 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 238364 -480 238476 240 8 la_oenb[100]
port 401 nsew signal input
rlabel metal2 s 240044 -480 240156 240 8 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 241724 -480 241836 240 8 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 243404 -480 243516 240 8 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 245084 -480 245196 240 8 la_oenb[104]
port 405 nsew signal input
rlabel metal2 s 246764 -480 246876 240 8 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 248444 -480 248556 240 8 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 250124 -480 250236 240 8 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 251804 -480 251916 240 8 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 253484 -480 253596 240 8 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 87164 -480 87276 240 8 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 255164 -480 255276 240 8 la_oenb[110]
port 412 nsew signal input
rlabel metal2 s 256844 -480 256956 240 8 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 258524 -480 258636 240 8 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 260204 -480 260316 240 8 la_oenb[113]
port 415 nsew signal input
rlabel metal2 s 261884 -480 261996 240 8 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 263564 -480 263676 240 8 la_oenb[115]
port 417 nsew signal input
rlabel metal2 s 265244 -480 265356 240 8 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 266924 -480 267036 240 8 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 268604 -480 268716 240 8 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 270284 -480 270396 240 8 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 88844 -480 88956 240 8 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 271964 -480 272076 240 8 la_oenb[120]
port 423 nsew signal input
rlabel metal2 s 273644 -480 273756 240 8 la_oenb[121]
port 424 nsew signal input
rlabel metal2 s 275324 -480 275436 240 8 la_oenb[122]
port 425 nsew signal input
rlabel metal2 s 277004 -480 277116 240 8 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 278684 -480 278796 240 8 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 280364 -480 280476 240 8 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 282044 -480 282156 240 8 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 283724 -480 283836 240 8 la_oenb[127]
port 430 nsew signal input
rlabel metal2 s 90524 -480 90636 240 8 la_oenb[12]
port 431 nsew signal input
rlabel metal2 s 92204 -480 92316 240 8 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 93884 -480 93996 240 8 la_oenb[14]
port 433 nsew signal input
rlabel metal2 s 95564 -480 95676 240 8 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 97244 -480 97356 240 8 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 98924 -480 99036 240 8 la_oenb[17]
port 436 nsew signal input
rlabel metal2 s 100604 -480 100716 240 8 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 102284 -480 102396 240 8 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 72044 -480 72156 240 8 la_oenb[1]
port 439 nsew signal input
rlabel metal2 s 103964 -480 104076 240 8 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 105644 -480 105756 240 8 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 107324 -480 107436 240 8 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 109004 -480 109116 240 8 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 110684 -480 110796 240 8 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 112364 -480 112476 240 8 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 114044 -480 114156 240 8 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 115724 -480 115836 240 8 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 117404 -480 117516 240 8 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 119084 -480 119196 240 8 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 73724 -480 73836 240 8 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 120764 -480 120876 240 8 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 122444 -480 122556 240 8 la_oenb[31]
port 452 nsew signal input
rlabel metal2 s 124124 -480 124236 240 8 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 125804 -480 125916 240 8 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 127484 -480 127596 240 8 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 129164 -480 129276 240 8 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 130844 -480 130956 240 8 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 132524 -480 132636 240 8 la_oenb[37]
port 458 nsew signal input
rlabel metal2 s 134204 -480 134316 240 8 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 135884 -480 135996 240 8 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 75404 -480 75516 240 8 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 137564 -480 137676 240 8 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 139244 -480 139356 240 8 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 140924 -480 141036 240 8 la_oenb[42]
port 464 nsew signal input
rlabel metal2 s 142604 -480 142716 240 8 la_oenb[43]
port 465 nsew signal input
rlabel metal2 s 144284 -480 144396 240 8 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 145964 -480 146076 240 8 la_oenb[45]
port 467 nsew signal input
rlabel metal2 s 147644 -480 147756 240 8 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 149324 -480 149436 240 8 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 151004 -480 151116 240 8 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 152684 -480 152796 240 8 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 77084 -480 77196 240 8 la_oenb[4]
port 472 nsew signal input
rlabel metal2 s 154364 -480 154476 240 8 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 156044 -480 156156 240 8 la_oenb[51]
port 474 nsew signal input
rlabel metal2 s 157724 -480 157836 240 8 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 159404 -480 159516 240 8 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 161084 -480 161196 240 8 la_oenb[54]
port 477 nsew signal input
rlabel metal2 s 162764 -480 162876 240 8 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 164444 -480 164556 240 8 la_oenb[56]
port 479 nsew signal input
rlabel metal2 s 166124 -480 166236 240 8 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 167804 -480 167916 240 8 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 169484 -480 169596 240 8 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 78764 -480 78876 240 8 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 171164 -480 171276 240 8 la_oenb[60]
port 484 nsew signal input
rlabel metal2 s 172844 -480 172956 240 8 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 174524 -480 174636 240 8 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 176204 -480 176316 240 8 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 177884 -480 177996 240 8 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 179564 -480 179676 240 8 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 181244 -480 181356 240 8 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 182924 -480 183036 240 8 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 184604 -480 184716 240 8 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 186284 -480 186396 240 8 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 80444 -480 80556 240 8 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 187964 -480 188076 240 8 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 189644 -480 189756 240 8 la_oenb[71]
port 496 nsew signal input
rlabel metal2 s 191324 -480 191436 240 8 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 193004 -480 193116 240 8 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 194684 -480 194796 240 8 la_oenb[74]
port 499 nsew signal input
rlabel metal2 s 196364 -480 196476 240 8 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 198044 -480 198156 240 8 la_oenb[76]
port 501 nsew signal input
rlabel metal2 s 199724 -480 199836 240 8 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 201404 -480 201516 240 8 la_oenb[78]
port 503 nsew signal input
rlabel metal2 s 203084 -480 203196 240 8 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 82124 -480 82236 240 8 la_oenb[7]
port 505 nsew signal input
rlabel metal2 s 204764 -480 204876 240 8 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 206444 -480 206556 240 8 la_oenb[81]
port 507 nsew signal input
rlabel metal2 s 208124 -480 208236 240 8 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 209804 -480 209916 240 8 la_oenb[83]
port 509 nsew signal input
rlabel metal2 s 211484 -480 211596 240 8 la_oenb[84]
port 510 nsew signal input
rlabel metal2 s 213164 -480 213276 240 8 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 214844 -480 214956 240 8 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 216524 -480 216636 240 8 la_oenb[87]
port 513 nsew signal input
rlabel metal2 s 218204 -480 218316 240 8 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 219884 -480 219996 240 8 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 83804 -480 83916 240 8 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 221564 -480 221676 240 8 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 223244 -480 223356 240 8 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 224924 -480 225036 240 8 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 226604 -480 226716 240 8 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 228284 -480 228396 240 8 la_oenb[94]
port 521 nsew signal input
rlabel metal2 s 229964 -480 230076 240 8 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 231644 -480 231756 240 8 la_oenb[96]
port 523 nsew signal input
rlabel metal2 s 233324 -480 233436 240 8 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 235004 -480 235116 240 8 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 236684 -480 236796 240 8 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 85484 -480 85596 240 8 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 284284 -480 284396 240 8 user_clock2
port 528 nsew signal input
rlabel metal2 s 284844 -480 284956 240 8 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 285404 -480 285516 240 8 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 285964 -480 286076 240 8 user_irq[2]
port 531 nsew signal output
rlabel metal4 s -478 -342 -168 298654 4 vdd
port 532 nsew power bidirectional
rlabel metal5 s -478 -342 298510 -32 8 vdd
port 532 nsew power bidirectional
rlabel metal5 s -478 298344 298510 298654 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 298200 -342 298510 298654 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 1577 -822 1887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 10577 -822 10887 79429 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 10577 229171 10887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 19577 -822 19887 79429 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 19577 229171 19887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 28577 -822 28887 38797 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 28577 55619 28887 79429 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 28577 229171 28887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 37577 -822 37887 38797 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 37577 55619 37887 79429 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 37577 229171 37887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 46577 -822 46887 38797 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 46577 55619 46887 79429 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 46577 229171 46887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 55577 -822 55887 38797 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 55577 55619 55887 79429 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 55577 229171 55887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 64577 -822 64887 38797 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 64577 55619 64887 79429 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 64577 229171 64887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 73577 -822 73887 38797 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 73577 55619 73887 79429 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 73577 229171 73887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 82577 -822 82887 38797 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 82577 55619 82887 79429 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 82577 229171 82887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 91577 -822 91887 79429 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 91577 229171 91887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 100577 -822 100887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 109577 -822 109887 4429 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 109577 74171 109887 79429 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 109577 229171 109887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 118577 -822 118887 4429 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 118577 74171 118887 79429 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 118577 229171 118887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 127577 -822 127887 4429 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 127577 74171 127887 79429 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 127577 229171 127887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 136577 -822 136887 4429 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 136577 74171 136887 79429 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 136577 229171 136887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 145577 -822 145887 4429 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 145577 74171 145887 79429 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 145577 229171 145887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 154577 -822 154887 4429 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 154577 74171 154887 79429 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 154577 229171 154887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 163577 -822 163887 4429 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 163577 74171 163887 79429 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 163577 229171 163887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 172577 -822 172887 4429 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 172577 74171 172887 79429 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 172577 229171 172887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 181577 -822 181887 4429 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 181577 74171 181887 79429 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 181577 229171 181887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 190577 -822 190887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 199577 -822 199887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 208577 -822 208887 79429 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 208577 229171 208887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 217577 -822 217887 79429 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 217577 229171 217887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 226577 -822 226887 79429 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 226577 229171 226887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 235577 -822 235887 79429 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 235577 229171 235887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 244577 -822 244887 79429 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 244577 229171 244887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 253577 -822 253887 79429 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 253577 229171 253887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 262577 -822 262887 79429 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 262577 229171 262887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 271577 -822 271887 79429 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 271577 229171 271887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 280577 -822 280887 79429 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 280577 229171 280887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 289577 -822 289887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 1913 298990 2223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 10913 298990 11223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 19913 298990 20223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 28913 298990 29223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 37913 298990 38223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 46913 298990 47223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 55913 298990 56223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 64913 298990 65223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 73913 298990 74223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 82913 298990 83223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 91913 298990 92223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 100913 298990 101223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 109913 298990 110223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 118913 298990 119223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 127913 298990 128223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 136913 298990 137223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 145913 298990 146223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 154913 298990 155223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 163913 298990 164223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 172913 298990 173223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 181913 298990 182223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 190913 298990 191223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 199913 298990 200223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 208913 298990 209223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 217913 298990 218223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 226913 298990 227223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 235913 298990 236223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 244913 298990 245223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 253913 298990 254223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 262913 298990 263223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 271913 298990 272223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 280913 298990 281223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 289913 298990 290223 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s -958 -822 -648 299134 4 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 -822 298990 -512 8 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 298824 298990 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 298680 -822 298990 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 3437 -822 3747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 12437 -822 12747 79429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 12437 149171 12747 159429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 12437 229171 12747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 21437 -822 21747 79429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 21437 149171 21747 159429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 21437 229171 21747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 30437 -822 30747 38797 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 30437 55619 30747 79429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 30437 149171 30747 159429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 30437 229171 30747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 39437 -822 39747 38797 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 39437 55619 39747 79429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 39437 149171 39747 159429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 39437 229171 39747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 48437 -822 48747 38797 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 48437 55619 48747 79429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 48437 149171 48747 159429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 48437 229171 48747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 57437 -822 57747 38797 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 57437 55619 57747 79429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 57437 149171 57747 159429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 57437 229171 57747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 66437 -822 66747 38797 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 66437 55619 66747 79429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 66437 149171 66747 159429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 66437 229171 66747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 75437 -822 75747 38797 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 75437 55619 75747 79429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 75437 149171 75747 159429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 75437 229171 75747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 84437 -822 84747 38797 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 84437 55619 84747 79429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 84437 149171 84747 159429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 84437 229171 84747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 93437 -822 93747 79429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 93437 149171 93747 159429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 93437 229171 93747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 102437 -822 102747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 111437 74171 111747 79429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 111437 149171 111747 159429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 111437 229171 111747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 120437 74171 120747 79429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 120437 149171 120747 159429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 120437 229171 120747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 129437 74171 129747 79429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 129437 149171 129747 159429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 129437 229171 129747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 138437 74171 138747 79429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 138437 149171 138747 159429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 138437 229171 138747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 147437 74171 147747 79429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 147437 149171 147747 159429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 147437 229171 147747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 156437 74171 156747 79429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 156437 149171 156747 159429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 156437 229171 156747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 165437 74171 165747 79429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 165437 149171 165747 159429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 165437 229171 165747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 174437 74171 174747 79429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 174437 149171 174747 159429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 174437 229171 174747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 183437 74171 183747 79429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 183437 149171 183747 159429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 183437 229171 183747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 192437 -822 192747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 201437 -822 201747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 210437 -822 210747 79429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 210437 149171 210747 159429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 210437 229171 210747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 219437 -822 219747 79429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 219437 149171 219747 159429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 219437 229171 219747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 228437 -822 228747 79429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 228437 149171 228747 159429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 228437 229171 228747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 237437 -822 237747 79429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 237437 149171 237747 159429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 237437 229171 237747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 246437 -822 246747 79429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 246437 149171 246747 159429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 246437 229171 246747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 255437 -822 255747 79429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 255437 149171 255747 159429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 255437 229171 255747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 264437 -822 264747 79429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 264437 149171 264747 159429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 264437 229171 264747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 273437 -822 273747 79429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 273437 149171 273747 159429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 273437 229171 273747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 282437 -822 282747 79429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 282437 149171 282747 159429 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 282437 229171 282747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 291437 -822 291747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 4913 298990 5223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 13913 298990 14223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 22913 298990 23223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 31913 298990 32223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 40913 298990 41223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 49913 298990 50223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 58913 298990 59223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 67913 298990 68223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 76913 298990 77223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 85913 298990 86223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 94913 298990 95223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 103913 298990 104223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 112913 298990 113223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 121913 298990 122223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 130913 298990 131223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 139913 298990 140223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 148913 298990 149223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 157913 298990 158223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 166913 298990 167223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 175913 298990 176223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 184913 298990 185223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 193913 298990 194223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 202913 298990 203223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 211913 298990 212223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 220913 298990 221223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 229913 298990 230223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 238913 298990 239223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 247913 298990 248223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 256913 298990 257223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 265913 298990 266223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 274913 298990 275223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 283913 298990 284223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 292913 298990 293223 6 vss
port 533 nsew ground bidirectional
rlabel metal2 s 9884 -480 9996 240 8 wb_clk_i
port 534 nsew signal input
rlabel metal2 s 10444 -480 10556 240 8 wb_rst_i
port 535 nsew signal input
rlabel metal2 s 11004 -480 11116 240 8 wbs_ack_o
port 536 nsew signal output
rlabel metal2 s 13244 -480 13356 240 8 wbs_adr_i[0]
port 537 nsew signal input
rlabel metal2 s 32284 -480 32396 240 8 wbs_adr_i[10]
port 538 nsew signal input
rlabel metal2 s 33964 -480 34076 240 8 wbs_adr_i[11]
port 539 nsew signal input
rlabel metal2 s 35644 -480 35756 240 8 wbs_adr_i[12]
port 540 nsew signal input
rlabel metal2 s 37324 -480 37436 240 8 wbs_adr_i[13]
port 541 nsew signal input
rlabel metal2 s 39004 -480 39116 240 8 wbs_adr_i[14]
port 542 nsew signal input
rlabel metal2 s 40684 -480 40796 240 8 wbs_adr_i[15]
port 543 nsew signal input
rlabel metal2 s 42364 -480 42476 240 8 wbs_adr_i[16]
port 544 nsew signal input
rlabel metal2 s 44044 -480 44156 240 8 wbs_adr_i[17]
port 545 nsew signal input
rlabel metal2 s 45724 -480 45836 240 8 wbs_adr_i[18]
port 546 nsew signal input
rlabel metal2 s 47404 -480 47516 240 8 wbs_adr_i[19]
port 547 nsew signal input
rlabel metal2 s 15484 -480 15596 240 8 wbs_adr_i[1]
port 548 nsew signal input
rlabel metal2 s 49084 -480 49196 240 8 wbs_adr_i[20]
port 549 nsew signal input
rlabel metal2 s 50764 -480 50876 240 8 wbs_adr_i[21]
port 550 nsew signal input
rlabel metal2 s 52444 -480 52556 240 8 wbs_adr_i[22]
port 551 nsew signal input
rlabel metal2 s 54124 -480 54236 240 8 wbs_adr_i[23]
port 552 nsew signal input
rlabel metal2 s 55804 -480 55916 240 8 wbs_adr_i[24]
port 553 nsew signal input
rlabel metal2 s 57484 -480 57596 240 8 wbs_adr_i[25]
port 554 nsew signal input
rlabel metal2 s 59164 -480 59276 240 8 wbs_adr_i[26]
port 555 nsew signal input
rlabel metal2 s 60844 -480 60956 240 8 wbs_adr_i[27]
port 556 nsew signal input
rlabel metal2 s 62524 -480 62636 240 8 wbs_adr_i[28]
port 557 nsew signal input
rlabel metal2 s 64204 -480 64316 240 8 wbs_adr_i[29]
port 558 nsew signal input
rlabel metal2 s 17724 -480 17836 240 8 wbs_adr_i[2]
port 559 nsew signal input
rlabel metal2 s 65884 -480 65996 240 8 wbs_adr_i[30]
port 560 nsew signal input
rlabel metal2 s 67564 -480 67676 240 8 wbs_adr_i[31]
port 561 nsew signal input
rlabel metal2 s 19964 -480 20076 240 8 wbs_adr_i[3]
port 562 nsew signal input
rlabel metal2 s 22204 -480 22316 240 8 wbs_adr_i[4]
port 563 nsew signal input
rlabel metal2 s 23884 -480 23996 240 8 wbs_adr_i[5]
port 564 nsew signal input
rlabel metal2 s 25564 -480 25676 240 8 wbs_adr_i[6]
port 565 nsew signal input
rlabel metal2 s 27244 -480 27356 240 8 wbs_adr_i[7]
port 566 nsew signal input
rlabel metal2 s 28924 -480 29036 240 8 wbs_adr_i[8]
port 567 nsew signal input
rlabel metal2 s 30604 -480 30716 240 8 wbs_adr_i[9]
port 568 nsew signal input
rlabel metal2 s 11564 -480 11676 240 8 wbs_cyc_i
port 569 nsew signal input
rlabel metal2 s 13804 -480 13916 240 8 wbs_dat_i[0]
port 570 nsew signal input
rlabel metal2 s 32844 -480 32956 240 8 wbs_dat_i[10]
port 571 nsew signal input
rlabel metal2 s 34524 -480 34636 240 8 wbs_dat_i[11]
port 572 nsew signal input
rlabel metal2 s 36204 -480 36316 240 8 wbs_dat_i[12]
port 573 nsew signal input
rlabel metal2 s 37884 -480 37996 240 8 wbs_dat_i[13]
port 574 nsew signal input
rlabel metal2 s 39564 -480 39676 240 8 wbs_dat_i[14]
port 575 nsew signal input
rlabel metal2 s 41244 -480 41356 240 8 wbs_dat_i[15]
port 576 nsew signal input
rlabel metal2 s 42924 -480 43036 240 8 wbs_dat_i[16]
port 577 nsew signal input
rlabel metal2 s 44604 -480 44716 240 8 wbs_dat_i[17]
port 578 nsew signal input
rlabel metal2 s 46284 -480 46396 240 8 wbs_dat_i[18]
port 579 nsew signal input
rlabel metal2 s 47964 -480 48076 240 8 wbs_dat_i[19]
port 580 nsew signal input
rlabel metal2 s 16044 -480 16156 240 8 wbs_dat_i[1]
port 581 nsew signal input
rlabel metal2 s 49644 -480 49756 240 8 wbs_dat_i[20]
port 582 nsew signal input
rlabel metal2 s 51324 -480 51436 240 8 wbs_dat_i[21]
port 583 nsew signal input
rlabel metal2 s 53004 -480 53116 240 8 wbs_dat_i[22]
port 584 nsew signal input
rlabel metal2 s 54684 -480 54796 240 8 wbs_dat_i[23]
port 585 nsew signal input
rlabel metal2 s 56364 -480 56476 240 8 wbs_dat_i[24]
port 586 nsew signal input
rlabel metal2 s 58044 -480 58156 240 8 wbs_dat_i[25]
port 587 nsew signal input
rlabel metal2 s 59724 -480 59836 240 8 wbs_dat_i[26]
port 588 nsew signal input
rlabel metal2 s 61404 -480 61516 240 8 wbs_dat_i[27]
port 589 nsew signal input
rlabel metal2 s 63084 -480 63196 240 8 wbs_dat_i[28]
port 590 nsew signal input
rlabel metal2 s 64764 -480 64876 240 8 wbs_dat_i[29]
port 591 nsew signal input
rlabel metal2 s 18284 -480 18396 240 8 wbs_dat_i[2]
port 592 nsew signal input
rlabel metal2 s 66444 -480 66556 240 8 wbs_dat_i[30]
port 593 nsew signal input
rlabel metal2 s 68124 -480 68236 240 8 wbs_dat_i[31]
port 594 nsew signal input
rlabel metal2 s 20524 -480 20636 240 8 wbs_dat_i[3]
port 595 nsew signal input
rlabel metal2 s 22764 -480 22876 240 8 wbs_dat_i[4]
port 596 nsew signal input
rlabel metal2 s 24444 -480 24556 240 8 wbs_dat_i[5]
port 597 nsew signal input
rlabel metal2 s 26124 -480 26236 240 8 wbs_dat_i[6]
port 598 nsew signal input
rlabel metal2 s 27804 -480 27916 240 8 wbs_dat_i[7]
port 599 nsew signal input
rlabel metal2 s 29484 -480 29596 240 8 wbs_dat_i[8]
port 600 nsew signal input
rlabel metal2 s 31164 -480 31276 240 8 wbs_dat_i[9]
port 601 nsew signal input
rlabel metal2 s 14364 -480 14476 240 8 wbs_dat_o[0]
port 602 nsew signal output
rlabel metal2 s 33404 -480 33516 240 8 wbs_dat_o[10]
port 603 nsew signal output
rlabel metal2 s 35084 -480 35196 240 8 wbs_dat_o[11]
port 604 nsew signal output
rlabel metal2 s 36764 -480 36876 240 8 wbs_dat_o[12]
port 605 nsew signal output
rlabel metal2 s 38444 -480 38556 240 8 wbs_dat_o[13]
port 606 nsew signal output
rlabel metal2 s 40124 -480 40236 240 8 wbs_dat_o[14]
port 607 nsew signal output
rlabel metal2 s 41804 -480 41916 240 8 wbs_dat_o[15]
port 608 nsew signal output
rlabel metal2 s 43484 -480 43596 240 8 wbs_dat_o[16]
port 609 nsew signal output
rlabel metal2 s 45164 -480 45276 240 8 wbs_dat_o[17]
port 610 nsew signal output
rlabel metal2 s 46844 -480 46956 240 8 wbs_dat_o[18]
port 611 nsew signal output
rlabel metal2 s 48524 -480 48636 240 8 wbs_dat_o[19]
port 612 nsew signal output
rlabel metal2 s 16604 -480 16716 240 8 wbs_dat_o[1]
port 613 nsew signal output
rlabel metal2 s 50204 -480 50316 240 8 wbs_dat_o[20]
port 614 nsew signal output
rlabel metal2 s 51884 -480 51996 240 8 wbs_dat_o[21]
port 615 nsew signal output
rlabel metal2 s 53564 -480 53676 240 8 wbs_dat_o[22]
port 616 nsew signal output
rlabel metal2 s 55244 -480 55356 240 8 wbs_dat_o[23]
port 617 nsew signal output
rlabel metal2 s 56924 -480 57036 240 8 wbs_dat_o[24]
port 618 nsew signal output
rlabel metal2 s 58604 -480 58716 240 8 wbs_dat_o[25]
port 619 nsew signal output
rlabel metal2 s 60284 -480 60396 240 8 wbs_dat_o[26]
port 620 nsew signal output
rlabel metal2 s 61964 -480 62076 240 8 wbs_dat_o[27]
port 621 nsew signal output
rlabel metal2 s 63644 -480 63756 240 8 wbs_dat_o[28]
port 622 nsew signal output
rlabel metal2 s 65324 -480 65436 240 8 wbs_dat_o[29]
port 623 nsew signal output
rlabel metal2 s 18844 -480 18956 240 8 wbs_dat_o[2]
port 624 nsew signal output
rlabel metal2 s 67004 -480 67116 240 8 wbs_dat_o[30]
port 625 nsew signal output
rlabel metal2 s 68684 -480 68796 240 8 wbs_dat_o[31]
port 626 nsew signal output
rlabel metal2 s 21084 -480 21196 240 8 wbs_dat_o[3]
port 627 nsew signal output
rlabel metal2 s 23324 -480 23436 240 8 wbs_dat_o[4]
port 628 nsew signal output
rlabel metal2 s 25004 -480 25116 240 8 wbs_dat_o[5]
port 629 nsew signal output
rlabel metal2 s 26684 -480 26796 240 8 wbs_dat_o[6]
port 630 nsew signal output
rlabel metal2 s 28364 -480 28476 240 8 wbs_dat_o[7]
port 631 nsew signal output
rlabel metal2 s 30044 -480 30156 240 8 wbs_dat_o[8]
port 632 nsew signal output
rlabel metal2 s 31724 -480 31836 240 8 wbs_dat_o[9]
port 633 nsew signal output
rlabel metal2 s 14924 -480 15036 240 8 wbs_sel_i[0]
port 634 nsew signal input
rlabel metal2 s 17164 -480 17276 240 8 wbs_sel_i[1]
port 635 nsew signal input
rlabel metal2 s 19404 -480 19516 240 8 wbs_sel_i[2]
port 636 nsew signal input
rlabel metal2 s 21644 -480 21756 240 8 wbs_sel_i[3]
port 637 nsew signal input
rlabel metal2 s 12124 -480 12236 240 8 wbs_stb_i
port 638 nsew signal input
rlabel metal2 s 12684 -480 12796 240 8 wbs_we_i
port 639 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 296020 296020
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 24981256
string GDS_FILE /home/jasteve4/Documents/MicroMotorController/openlane/user_project_wrapper/runs/22_12_05_23_39/results/signoff/user_project_wrapper.magic.gds
string GDS_START 23065200
<< end >>


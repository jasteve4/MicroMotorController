* NGSPICE file created from user_project_wrapper.ext - technology: gf180mcuC

* Black-box entry subcircuit for controller_core abstract view
.subckt controller_core clock clock_out[0] clock_out[1] clock_out[2] clock_out[3]
+ clock_out[4] clock_out[5] clock_out[6] clock_out[7] clock_out[8] clock_out[9] col_select_left[0]
+ col_select_left[1] col_select_left[2] col_select_left[3] col_select_left[4] col_select_left[5]
+ col_select_right[0] col_select_right[1] col_select_right[2] col_select_right[3]
+ col_select_right[4] col_select_right[5] data_out_left[0] data_out_left[10] data_out_left[11]
+ data_out_left[12] data_out_left[13] data_out_left[14] data_out_left[15] data_out_left[1]
+ data_out_left[2] data_out_left[3] data_out_left[4] data_out_left[5] data_out_left[6]
+ data_out_left[7] data_out_left[8] data_out_left[9] data_out_right[0] data_out_right[10]
+ data_out_right[11] data_out_right[12] data_out_right[13] data_out_right[14] data_out_right[15]
+ data_out_right[1] data_out_right[2] data_out_right[3] data_out_right[4] data_out_right[5]
+ data_out_right[6] data_out_right[7] data_out_right[8] data_out_right[9] inverter_select[0]
+ inverter_select[1] inverter_select[2] inverter_select[3] inverter_select[4] inverter_select[5]
+ inverter_select[6] inverter_select[7] inverter_select[8] inverter_select[9] io_control_trigger_in
+ io_control_trigger_oeb io_driver_io_oeb[0] io_driver_io_oeb[10] io_driver_io_oeb[11]
+ io_driver_io_oeb[12] io_driver_io_oeb[13] io_driver_io_oeb[14] io_driver_io_oeb[15]
+ io_driver_io_oeb[16] io_driver_io_oeb[17] io_driver_io_oeb[18] io_driver_io_oeb[19]
+ io_driver_io_oeb[1] io_driver_io_oeb[2] io_driver_io_oeb[3] io_driver_io_oeb[4]
+ io_driver_io_oeb[5] io_driver_io_oeb[6] io_driver_io_oeb[7] io_driver_io_oeb[8]
+ io_driver_io_oeb[9] io_latch_data_in io_latch_data_oeb io_reset_n_in io_reset_n_oeb
+ io_update_cycle_complete_oeb io_update_cycle_complete_out la_data_in[0] la_data_in[10]
+ la_data_in[11] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[1] la_data_in[2] la_data_in[3] la_data_in[4] la_data_in[5]
+ la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9] la_oenb[0] la_oenb[10] la_oenb[11]
+ la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[1]
+ la_oenb[2] la_oenb[3] la_oenb[4] la_oenb[5] la_oenb[6] la_oenb[7] la_oenb[8] la_oenb[9]
+ mem_address_left[0] mem_address_left[1] mem_address_left[2] mem_address_left[3]
+ mem_address_left[4] mem_address_left[5] mem_address_left[6] mem_address_left[7]
+ mem_address_left[8] mem_address_left[9] mem_address_right[0] mem_address_right[1]
+ mem_address_right[2] mem_address_right[3] mem_address_right[4] mem_address_right[5]
+ mem_address_right[6] mem_address_right[7] mem_address_right[8] mem_address_right[9]
+ mem_write_n[0] mem_write_n[1] mem_write_n[2] mem_write_n[3] mem_write_n[4] mem_write_n[5]
+ mem_write_n[6] mem_write_n[7] mem_write_n[8] mem_write_n[9] output_active_left output_active_right
+ row_col_select[0] row_col_select[1] row_col_select[2] row_col_select[3] row_col_select[4]
+ row_col_select[5] row_col_select[6] row_col_select[7] row_col_select[8] row_col_select[9]
+ row_select_left[0] row_select_left[1] row_select_left[2] row_select_left[3] row_select_left[4]
+ row_select_left[5] row_select_right[0] row_select_right[1] row_select_right[2] row_select_right[3]
+ row_select_right[4] row_select_right[5] spi_data[0] spi_data[10] spi_data[11] spi_data[12]
+ spi_data[13] spi_data[14] spi_data[15] spi_data[16] spi_data[17] spi_data[18] spi_data[19]
+ spi_data[1] spi_data[20] spi_data[21] spi_data[22] spi_data[23] spi_data[24] spi_data[25]
+ spi_data[26] spi_data[27] spi_data[28] spi_data[29] spi_data[2] spi_data[30] spi_data[31]
+ spi_data[3] spi_data[4] spi_data[5] spi_data[6] spi_data[7] spi_data[8] spi_data[9]
+ spi_data_clock vccd1 vssd1
.ends

* Black-box entry subcircuit for driver_core abstract view
.subckt driver_core clock clock_a col_select_a[0] col_select_a[1] col_select_a[2]
+ col_select_a[3] col_select_a[4] col_select_a[5] data_in_a[0] data_in_a[10] data_in_a[11]
+ data_in_a[12] data_in_a[13] data_in_a[14] data_in_a[15] data_in_a[1] data_in_a[2]
+ data_in_a[3] data_in_a[4] data_in_a[5] data_in_a[6] data_in_a[7] data_in_a[8] data_in_a[9]
+ driver_io[0] driver_io[1] inverter_select_a mem_address_a[0] mem_address_a[1] mem_address_a[2]
+ mem_address_a[3] mem_address_a[4] mem_address_a[5] mem_address_a[6] mem_address_a[7]
+ mem_address_a[8] mem_address_a[9] mem_write_n_a output_active_a row_col_select_a
+ row_select_a[0] row_select_a[1] row_select_a[2] row_select_a[3] row_select_a[4]
+ row_select_a[5] vccd1 vssd1
.ends

* Black-box entry subcircuit for clock_mux abstract view
.subckt clock_mux clock_out_a clock_out_b clock_out_c core_clock io_clock la_oenb
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for spi_core abstract view
.subckt spi_core clock clock_out data_out[0] data_out[10] data_out[11] data_out[12]
+ data_out[13] data_out[14] data_out[15] data_out[16] data_out[17] data_out[18] data_out[19]
+ data_out[1] data_out[20] data_out[21] data_out[22] data_out[23] data_out[24] data_out[25]
+ data_out[26] data_out[27] data_out[28] data_out[29] data_out[2] data_out[30] data_out[31]
+ data_out[3] data_out[4] data_out[5] data_out[6] data_out[7] data_out[8] data_out[9]
+ la_data_in[0] la_data_in[1] la_data_in[2] la_data_in[3] la_oenb[0] la_oenb[1] la_oenb[2]
+ la_oenb[3] miso miso_oeb mosi mosi_oeb sclk sclk_oeb ss_n ss_n_oeb vccd1 vssd1
.ends

.subckt user_project_wrapper analog_io[0] analog_io[10] analog_io[11] analog_io[12]
+ analog_io[13] analog_io[14] analog_io[15] analog_io[16] analog_io[17] analog_io[18]
+ analog_io[19] analog_io[1] analog_io[20] analog_io[21] analog_io[22] analog_io[23]
+ analog_io[24] analog_io[25] analog_io[26] analog_io[27] analog_io[28] analog_io[2]
+ analog_io[3] analog_io[4] analog_io[5] analog_io[6] analog_io[7] analog_io[8] analog_io[9]
+ io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36]
+ io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30]
+ io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100]
+ la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105]
+ la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110]
+ la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115]
+ la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120]
+ la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125]
+ la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15]
+ la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20]
+ la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42]
+ la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48]
+ la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53]
+ la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59]
+ la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64]
+ la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6]
+ la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75]
+ la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80]
+ la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86]
+ la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91]
+ la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97]
+ la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101]
+ la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106]
+ la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110]
+ la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115]
+ la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11]
+ la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124]
+ la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18]
+ la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28]
+ la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33]
+ la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38]
+ la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43]
+ la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48]
+ la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58]
+ la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63]
+ la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68]
+ la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73]
+ la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78]
+ la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83]
+ la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88]
+ la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93]
+ la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98]
+ la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102]
+ la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109]
+ la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115]
+ la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121]
+ la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12]
+ la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19]
+ la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25]
+ la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31]
+ la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38]
+ la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44]
+ la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50]
+ la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57]
+ la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63]
+ la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6]
+ la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76]
+ la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82]
+ la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89]
+ la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95]
+ la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0]
+ user_irq[1] user_irq[2] vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
Xcontroller_core_mod clock_out_c clock_out\[0\] clock_out\[1\] clock_out\[2\] clock_out\[3\]
+ clock_out\[4\] clock_out\[5\] clock_out\[6\] clock_out\[7\] clock_out\[8\] clock_out\[9\]
+ col_select_left\[0\] col_select_left\[1\] col_select_left\[2\] col_select_left\[3\]
+ col_select_left\[4\] col_select_left\[5\] col_select_right\[0\] col_select_right\[1\]
+ col_select_right\[2\] col_select_right\[3\] col_select_right\[4\] col_select_right\[5\]
+ data_out_left\[0\] data_out_left\[10\] data_out_left\[11\] data_out_left\[12\] data_out_left\[13\]
+ data_out_left\[14\] data_out_left\[15\] data_out_left\[1\] data_out_left\[2\] data_out_left\[3\]
+ data_out_left\[4\] data_out_left\[5\] data_out_left\[6\] data_out_left\[7\] data_out_left\[8\]
+ data_out_left\[9\] data_out_right\[0\] data_out_right\[10\] data_out_right\[11\]
+ data_out_right\[12\] data_out_right\[13\] data_out_right\[14\] data_out_right\[15\]
+ data_out_right\[1\] data_out_right\[2\] data_out_right\[3\] data_out_right\[4\]
+ data_out_right\[5\] data_out_right\[6\] data_out_right\[7\] data_out_right\[8\]
+ data_out_right\[9\] inverter_select\[0\] inverter_select\[1\] inverter_select\[2\]
+ inverter_select\[3\] inverter_select\[4\] inverter_select\[5\] inverter_select\[6\]
+ inverter_select\[7\] inverter_select\[8\] inverter_select\[9\] io_in[36] io_oeb[36]
+ io_oeb[29] io_oeb[17] io_oeb[16] io_oeb[15] io_oeb[14] io_oeb[13] io_oeb[12] io_oeb[11]
+ io_oeb[10] io_oeb[9] io_oeb[8] io_oeb[28] io_oeb[27] io_oeb[26] io_oeb[25] io_oeb[24]
+ io_oeb[23] io_oeb[22] io_oeb[21] io_oeb[20] io_in[35] io_oeb[35] io_in[37] io_oeb[37]
+ io_oeb[30] io_out[30] la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12]
+ la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[1]
+ la_data_in[2] la_data_in[3] la_data_in[4] la_data_in[5] la_data_in[6] la_data_in[7]
+ la_data_in[8] la_data_in[9] la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13]
+ la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[1] la_oenb[2] la_oenb[3]
+ la_oenb[4] la_oenb[5] la_oenb[6] la_oenb[7] la_oenb[8] la_oenb[9] mem_address_left\[0\]
+ mem_address_left\[1\] mem_address_left\[2\] mem_address_left\[3\] mem_address_left\[4\]
+ mem_address_left\[5\] mem_address_left\[6\] mem_address_left\[7\] mem_address_left\[8\]
+ mem_address_left\[9\] mem_address_right\[0\] mem_address_right\[1\] mem_address_right\[2\]
+ mem_address_right\[3\] mem_address_right\[4\] mem_address_right\[5\] mem_address_right\[6\]
+ mem_address_right\[7\] mem_address_right\[8\] mem_address_right\[9\] mem_write_n\[0\]
+ mem_write_n\[1\] mem_write_n\[2\] mem_write_n\[3\] mem_write_n\[4\] mem_write_n\[5\]
+ mem_write_n\[6\] mem_write_n\[7\] mem_write_n\[8\] mem_write_n\[9\] output_active_left
+ output_active_right row_col_select\[0\] row_col_select\[1\] row_col_select\[2\]
+ row_col_select\[3\] row_col_select\[4\] row_col_select\[5\] row_col_select\[6\]
+ row_col_select\[7\] row_col_select\[8\] row_col_select\[9\] row_select_left\[0\]
+ row_select_left\[1\] row_select_left\[2\] row_select_left\[3\] row_select_left\[4\]
+ row_select_left\[5\] row_select_right\[0\] row_select_right\[1\] row_select_right\[2\]
+ row_select_right\[3\] row_select_right\[4\] row_select_right\[5\] spi_data\[0\]
+ spi_data\[10\] spi_data\[11\] spi_data\[12\] spi_data\[13\] spi_data\[14\] spi_data\[15\]
+ spi_data\[16\] spi_data\[17\] spi_data\[18\] spi_data\[19\] spi_data\[1\] spi_data\[20\]
+ spi_data\[21\] spi_data\[22\] spi_data\[23\] spi_data\[24\] spi_data\[25\] spi_data\[26\]
+ spi_data\[27\] spi_data\[28\] spi_data\[29\] spi_data\[2\] spi_data\[30\] spi_data\[31\]
+ spi_data\[3\] spi_data\[4\] spi_data\[5\] spi_data\[6\] spi_data\[7\] spi_data\[8\]
+ spi_data\[9\] spi_data_clock vccd1 vssd1 controller_core
Xdriver_core_0 clock_out_c clock_out\[0\] col_select_left\[0\] col_select_left\[1\]
+ col_select_left\[2\] col_select_left\[3\] col_select_left\[4\] col_select_left\[5\]
+ data_out_left\[0\] data_out_left\[10\] data_out_left\[11\] data_out_left\[12\] data_out_left\[13\]
+ data_out_left\[14\] data_out_left\[15\] data_out_left\[1\] data_out_left\[2\] data_out_left\[3\]
+ data_out_left\[4\] data_out_left\[5\] data_out_left\[6\] data_out_left\[7\] data_out_left\[8\]
+ data_out_left\[9\] io_out[29] io_out[28] inverter_select\[0\] mem_address_left\[0\]
+ mem_address_left\[1\] mem_address_left\[2\] mem_address_left\[3\] mem_address_left\[4\]
+ mem_address_left\[5\] mem_address_left\[6\] mem_address_left\[7\] mem_address_left\[8\]
+ mem_address_left\[9\] mem_write_n\[0\] output_active_left row_col_select\[0\] row_select_left\[0\]
+ row_select_left\[1\] row_select_left\[2\] row_select_left\[3\] row_select_left\[4\]
+ row_select_left\[5\] driver_core_0/vccd1 driver_core_0/vssd1 driver_core
Xdriver_core_1 clock_out_a clock_out\[1\] col_select_left\[0\] col_select_left\[1\]
+ col_select_left\[2\] col_select_left\[3\] col_select_left\[4\] col_select_left\[5\]
+ data_out_left\[0\] data_out_left\[10\] data_out_left\[11\] data_out_left\[12\] data_out_left\[13\]
+ data_out_left\[14\] data_out_left\[15\] data_out_left\[1\] data_out_left\[2\] data_out_left\[3\]
+ data_out_left\[4\] data_out_left\[5\] data_out_left\[6\] data_out_left\[7\] data_out_left\[8\]
+ data_out_left\[9\] io_out[27] io_out[26] inverter_select\[1\] mem_address_left\[0\]
+ mem_address_left\[1\] mem_address_left\[2\] mem_address_left\[3\] mem_address_left\[4\]
+ mem_address_left\[5\] mem_address_left\[6\] mem_address_left\[7\] mem_address_left\[8\]
+ mem_address_left\[9\] mem_write_n\[1\] output_active_left row_col_select\[1\] row_select_left\[0\]
+ row_select_left\[1\] row_select_left\[2\] row_select_left\[3\] row_select_left\[4\]
+ row_select_left\[5\] driver_core_1/vccd1 driver_core_1/vssd1 driver_core
Xdriver_core_2 clock_out_a clock_out\[2\] col_select_left\[0\] col_select_left\[1\]
+ col_select_left\[2\] col_select_left\[3\] col_select_left\[4\] col_select_left\[5\]
+ data_out_left\[0\] data_out_left\[10\] data_out_left\[11\] data_out_left\[12\] data_out_left\[13\]
+ data_out_left\[14\] data_out_left\[15\] data_out_left\[1\] data_out_left\[2\] data_out_left\[3\]
+ data_out_left\[4\] data_out_left\[5\] data_out_left\[6\] data_out_left\[7\] data_out_left\[8\]
+ data_out_left\[9\] io_out[25] io_out[24] inverter_select\[2\] mem_address_left\[0\]
+ mem_address_left\[1\] mem_address_left\[2\] mem_address_left\[3\] mem_address_left\[4\]
+ mem_address_left\[5\] mem_address_left\[6\] mem_address_left\[7\] mem_address_left\[8\]
+ mem_address_left\[9\] mem_write_n\[2\] output_active_left row_col_select\[2\] row_select_left\[0\]
+ row_select_left\[1\] row_select_left\[2\] row_select_left\[3\] row_select_left\[4\]
+ row_select_left\[5\] driver_core_2/vccd1 driver_core_2/vssd1 driver_core
Xdriver_core_3 clock_out_a clock_out\[3\] col_select_left\[0\] col_select_left\[1\]
+ col_select_left\[2\] col_select_left\[3\] col_select_left\[4\] col_select_left\[5\]
+ data_out_left\[0\] data_out_left\[10\] data_out_left\[11\] data_out_left\[12\] data_out_left\[13\]
+ data_out_left\[14\] data_out_left\[15\] data_out_left\[1\] data_out_left\[2\] data_out_left\[3\]
+ data_out_left\[4\] data_out_left\[5\] data_out_left\[6\] data_out_left\[7\] data_out_left\[8\]
+ data_out_left\[9\] io_out[23] io_out[22] inverter_select\[3\] mem_address_left\[0\]
+ mem_address_left\[1\] mem_address_left\[2\] mem_address_left\[3\] mem_address_left\[4\]
+ mem_address_left\[5\] mem_address_left\[6\] mem_address_left\[7\] mem_address_left\[8\]
+ mem_address_left\[9\] mem_write_n\[3\] output_active_left row_col_select\[3\] row_select_left\[0\]
+ row_select_left\[1\] row_select_left\[2\] row_select_left\[3\] row_select_left\[4\]
+ row_select_left\[5\] driver_core_3/vccd1 driver_core_3/vssd1 driver_core
Xdriver_core_4 clock_out_a clock_out\[4\] col_select_left\[0\] col_select_left\[1\]
+ col_select_left\[2\] col_select_left\[3\] col_select_left\[4\] col_select_left\[5\]
+ data_out_left\[0\] data_out_left\[10\] data_out_left\[11\] data_out_left\[12\] data_out_left\[13\]
+ data_out_left\[14\] data_out_left\[15\] data_out_left\[1\] data_out_left\[2\] data_out_left\[3\]
+ data_out_left\[4\] data_out_left\[5\] data_out_left\[6\] data_out_left\[7\] data_out_left\[8\]
+ data_out_left\[9\] io_out[21] io_out[20] inverter_select\[4\] mem_address_left\[0\]
+ mem_address_left\[1\] mem_address_left\[2\] mem_address_left\[3\] mem_address_left\[4\]
+ mem_address_left\[5\] mem_address_left\[6\] mem_address_left\[7\] mem_address_left\[8\]
+ mem_address_left\[9\] mem_write_n\[4\] output_active_left row_col_select\[4\] row_select_left\[0\]
+ row_select_left\[1\] row_select_left\[2\] row_select_left\[3\] row_select_left\[4\]
+ row_select_left\[5\] driver_core_4/vccd1 driver_core_4/vssd1 driver_core
Xdriver_core_5 clock_out_b clock_out\[5\] col_select_right\[0\] col_select_right\[1\]
+ col_select_right\[2\] col_select_right\[3\] col_select_right\[4\] col_select_right\[5\]
+ data_out_right\[0\] data_out_right\[10\] data_out_right\[11\] data_out_right\[12\]
+ data_out_right\[13\] data_out_right\[14\] data_out_right\[15\] data_out_right\[1\]
+ data_out_right\[2\] data_out_right\[3\] data_out_right\[4\] data_out_right\[5\]
+ data_out_right\[6\] data_out_right\[7\] data_out_right\[8\] data_out_right\[9\]
+ io_out[18] io_out[17] inverter_select\[5\] mem_address_right\[0\] mem_address_right\[1\]
+ mem_address_right\[2\] mem_address_right\[3\] mem_address_right\[4\] mem_address_right\[5\]
+ mem_address_right\[6\] mem_address_right\[7\] mem_address_right\[8\] mem_address_right\[9\]
+ mem_write_n\[5\] output_active_right row_col_select\[5\] row_select_right\[0\] row_select_right\[1\]
+ row_select_right\[2\] row_select_right\[3\] row_select_right\[4\] row_select_right\[5\]
+ driver_core_5/vccd1 driver_core_5/vssd1 driver_core
Xdriver_core_6 clock_out_b clock_out\[6\] col_select_right\[0\] col_select_right\[1\]
+ col_select_right\[2\] col_select_right\[3\] col_select_right\[4\] col_select_right\[5\]
+ data_out_right\[0\] data_out_right\[10\] data_out_right\[11\] data_out_right\[12\]
+ data_out_right\[13\] data_out_right\[14\] data_out_right\[15\] data_out_right\[1\]
+ data_out_right\[2\] data_out_right\[3\] data_out_right\[4\] data_out_right\[5\]
+ data_out_right\[6\] data_out_right\[7\] data_out_right\[8\] data_out_right\[9\]
+ io_out[16] io_out[15] inverter_select\[6\] mem_address_right\[0\] mem_address_right\[1\]
+ mem_address_right\[2\] mem_address_right\[3\] mem_address_right\[4\] mem_address_right\[5\]
+ mem_address_right\[6\] mem_address_right\[7\] mem_address_right\[8\] mem_address_right\[9\]
+ mem_write_n\[6\] output_active_right row_col_select\[6\] row_select_right\[0\] row_select_right\[1\]
+ row_select_right\[2\] row_select_right\[3\] row_select_right\[4\] row_select_right\[5\]
+ driver_core_6/vccd1 driver_core_6/vssd1 driver_core
Xdriver_core_7 clock_out_b clock_out\[7\] col_select_right\[0\] col_select_right\[1\]
+ col_select_right\[2\] col_select_right\[3\] col_select_right\[4\] col_select_right\[5\]
+ data_out_right\[0\] data_out_right\[10\] data_out_right\[11\] data_out_right\[12\]
+ data_out_right\[13\] data_out_right\[14\] data_out_right\[15\] data_out_right\[1\]
+ data_out_right\[2\] data_out_right\[3\] data_out_right\[4\] data_out_right\[5\]
+ data_out_right\[6\] data_out_right\[7\] data_out_right\[8\] data_out_right\[9\]
+ io_out[14] io_out[13] inverter_select\[7\] mem_address_right\[0\] mem_address_right\[1\]
+ mem_address_right\[2\] mem_address_right\[3\] mem_address_right\[4\] mem_address_right\[5\]
+ mem_address_right\[6\] mem_address_right\[7\] mem_address_right\[8\] mem_address_right\[9\]
+ mem_write_n\[7\] output_active_right row_col_select\[7\] row_select_right\[0\] row_select_right\[1\]
+ row_select_right\[2\] row_select_right\[3\] row_select_right\[4\] row_select_right\[5\]
+ driver_core_7/vccd1 driver_core_7/vssd1 driver_core
Xdriver_core_8 clock_out_b clock_out\[8\] col_select_right\[0\] col_select_right\[1\]
+ col_select_right\[2\] col_select_right\[3\] col_select_right\[4\] col_select_right\[5\]
+ data_out_right\[0\] data_out_right\[10\] data_out_right\[11\] data_out_right\[12\]
+ data_out_right\[13\] data_out_right\[14\] data_out_right\[15\] data_out_right\[1\]
+ data_out_right\[2\] data_out_right\[3\] data_out_right\[4\] data_out_right\[5\]
+ data_out_right\[6\] data_out_right\[7\] data_out_right\[8\] data_out_right\[9\]
+ io_out[12] io_out[11] inverter_select\[8\] mem_address_right\[0\] mem_address_right\[1\]
+ mem_address_right\[2\] mem_address_right\[3\] mem_address_right\[4\] mem_address_right\[5\]
+ mem_address_right\[6\] mem_address_right\[7\] mem_address_right\[8\] mem_address_right\[9\]
+ mem_write_n\[8\] output_active_right row_col_select\[8\] row_select_right\[0\] row_select_right\[1\]
+ row_select_right\[2\] row_select_right\[3\] row_select_right\[4\] row_select_right\[5\]
+ driver_core_8/vccd1 driver_core_8/vssd1 driver_core
Xclock_mux_mod clock_out_a clock_out_b clock_out_c user_clock2 io_in[8] la_oenb[63]
+ clock_mux_mod/vccd1 clock_mux_mod/vssd1 clock_mux
Xdriver_core_9 clock_out_c clock_out\[9\] col_select_right\[0\] col_select_right\[1\]
+ col_select_right\[2\] col_select_right\[3\] col_select_right\[4\] col_select_right\[5\]
+ data_out_right\[0\] data_out_right\[10\] data_out_right\[11\] data_out_right\[12\]
+ data_out_right\[13\] data_out_right\[14\] data_out_right\[15\] data_out_right\[1\]
+ data_out_right\[2\] data_out_right\[3\] data_out_right\[4\] data_out_right\[5\]
+ data_out_right\[6\] data_out_right\[7\] data_out_right\[8\] data_out_right\[9\]
+ io_out[10] io_out[9] inverter_select\[9\] mem_address_right\[0\] mem_address_right\[1\]
+ mem_address_right\[2\] mem_address_right\[3\] mem_address_right\[4\] mem_address_right\[5\]
+ mem_address_right\[6\] mem_address_right\[7\] mem_address_right\[8\] mem_address_right\[9\]
+ mem_write_n\[9\] output_active_right row_col_select\[9\] row_select_right\[0\] row_select_right\[1\]
+ row_select_right\[2\] row_select_right\[3\] row_select_right\[4\] row_select_right\[5\]
+ driver_core_9/vccd1 driver_core_9/vssd1 driver_core
Xspi_core_mod clock_out_c spi_data_clock spi_data\[0\] spi_data\[10\] spi_data\[11\]
+ spi_data\[12\] spi_data\[13\] spi_data\[14\] spi_data\[15\] spi_data\[16\] spi_data\[17\]
+ spi_data\[18\] spi_data\[19\] spi_data\[1\] spi_data\[20\] spi_data\[21\] spi_data\[22\]
+ spi_data\[23\] spi_data\[24\] spi_data\[25\] spi_data\[26\] spi_data\[27\] spi_data\[28\]
+ spi_data\[29\] spi_data\[2\] spi_data\[30\] spi_data\[31\] spi_data\[3\] spi_data\[4\]
+ spi_data\[5\] spi_data\[6\] spi_data\[7\] spi_data\[8\] spi_data\[9\] la_data_in[17]
+ la_data_in[18] la_data_in[19] la_data_in[20] la_oenb[17] la_oenb[18] la_oenb[19]
+ la_oenb[20] io_out[34] io_oeb[34] io_in[33] io_oeb[33] io_in[31] io_oeb[31] io_in[32]
+ io_oeb[32] spi_core_mod/vccd1 spi_core_mod/vssd1 spi_core
.ends


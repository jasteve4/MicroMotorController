VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO clock_mux
  CLASS BLOCK ;
  FOREIGN clock_mux ;
  ORIGIN 0.000 0.000 ;
  SIZE 250.000 BY 250.000 ;
  PIN clock_out_a
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 41.440 4.000 42.000 ;
    END
  END clock_out_a
  PIN clock_out_b
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 124.320 4.000 124.880 ;
    END
  END clock_out_b
  PIN clock_out_c
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 207.200 4.000 207.760 ;
    END
  END clock_out_c
  PIN core_clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 62.160 0.000 62.720 4.000 ;
    END
  END core_clock
  PIN io_clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 124.320 250.000 124.880 ;
    END
  END io_clock
  PIN la_oenb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 187.040 0.000 187.600 4.000 ;
    END
  END la_oenb
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 231.580 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 231.580 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 231.580 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 243.040 231.580 ;
      LAYER Metal2 ;
        RECT 8.540 4.300 224.420 231.470 ;
        RECT 8.540 3.500 61.860 4.300 ;
        RECT 63.020 3.500 186.740 4.300 ;
        RECT 187.900 3.500 224.420 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 208.060 246.000 231.420 ;
        RECT 4.300 206.900 246.000 208.060 ;
        RECT 4.000 125.180 246.000 206.900 ;
        RECT 4.300 124.020 245.700 125.180 ;
        RECT 4.000 42.300 246.000 124.020 ;
        RECT 4.300 41.140 246.000 42.300 ;
        RECT 4.000 15.540 246.000 41.140 ;
  END
END clock_mux
END LIBRARY


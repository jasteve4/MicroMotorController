magic
tech gf180mcuC
magscale 1 5
timestamp 1670271749
<< obsm1 >>
rect 5672 6538 294320 295198
<< metal2 >>
rect 4900 299760 5012 300480
rect 13188 299760 13300 300480
rect 21476 299760 21588 300480
rect 29764 299760 29876 300480
rect 38052 299760 38164 300480
rect 46340 299760 46452 300480
rect 54628 299760 54740 300480
rect 62916 299760 63028 300480
rect 71204 299760 71316 300480
rect 79492 299760 79604 300480
rect 87780 299760 87892 300480
rect 96068 299760 96180 300480
rect 104356 299760 104468 300480
rect 112644 299760 112756 300480
rect 120932 299760 121044 300480
rect 129220 299760 129332 300480
rect 137508 299760 137620 300480
rect 145796 299760 145908 300480
rect 154084 299760 154196 300480
rect 162372 299760 162484 300480
rect 170660 299760 170772 300480
rect 178948 299760 179060 300480
rect 187236 299760 187348 300480
rect 195524 299760 195636 300480
rect 203812 299760 203924 300480
rect 212100 299760 212212 300480
rect 220388 299760 220500 300480
rect 228676 299760 228788 300480
rect 236964 299760 237076 300480
rect 245252 299760 245364 300480
rect 253540 299760 253652 300480
rect 261828 299760 261940 300480
rect 270116 299760 270228 300480
rect 278404 299760 278516 300480
rect 286692 299760 286804 300480
rect 294980 299760 295092 300480
rect 11900 -480 12012 240
rect 12460 -480 12572 240
rect 13020 -480 13132 240
rect 13580 -480 13692 240
rect 14140 -480 14252 240
rect 14700 -480 14812 240
rect 15260 -480 15372 240
rect 15820 -480 15932 240
rect 16380 -480 16492 240
rect 16940 -480 17052 240
rect 17500 -480 17612 240
rect 18060 -480 18172 240
rect 18620 -480 18732 240
rect 19180 -480 19292 240
rect 19740 -480 19852 240
rect 20300 -480 20412 240
rect 20860 -480 20972 240
rect 21420 -480 21532 240
rect 21980 -480 22092 240
rect 22540 -480 22652 240
rect 23100 -480 23212 240
rect 23660 -480 23772 240
rect 24220 -480 24332 240
rect 24780 -480 24892 240
rect 25340 -480 25452 240
rect 25900 -480 26012 240
rect 26460 -480 26572 240
rect 27020 -480 27132 240
rect 27580 -480 27692 240
rect 28140 -480 28252 240
rect 28700 -480 28812 240
rect 29260 -480 29372 240
rect 29820 -480 29932 240
rect 30380 -480 30492 240
rect 30940 -480 31052 240
rect 31500 -480 31612 240
rect 32060 -480 32172 240
rect 32620 -480 32732 240
rect 33180 -480 33292 240
rect 33740 -480 33852 240
rect 34300 -480 34412 240
rect 34860 -480 34972 240
rect 35420 -480 35532 240
rect 35980 -480 36092 240
rect 36540 -480 36652 240
rect 37100 -480 37212 240
rect 37660 -480 37772 240
rect 38220 -480 38332 240
rect 38780 -480 38892 240
rect 39340 -480 39452 240
rect 39900 -480 40012 240
rect 40460 -480 40572 240
rect 41020 -480 41132 240
rect 41580 -480 41692 240
rect 42140 -480 42252 240
rect 42700 -480 42812 240
rect 43260 -480 43372 240
rect 43820 -480 43932 240
rect 44380 -480 44492 240
rect 44940 -480 45052 240
rect 45500 -480 45612 240
rect 46060 -480 46172 240
rect 46620 -480 46732 240
rect 47180 -480 47292 240
rect 47740 -480 47852 240
rect 48300 -480 48412 240
rect 48860 -480 48972 240
rect 49420 -480 49532 240
rect 49980 -480 50092 240
rect 50540 -480 50652 240
rect 51100 -480 51212 240
rect 51660 -480 51772 240
rect 52220 -480 52332 240
rect 52780 -480 52892 240
rect 53340 -480 53452 240
rect 53900 -480 54012 240
rect 54460 -480 54572 240
rect 55020 -480 55132 240
rect 55580 -480 55692 240
rect 56140 -480 56252 240
rect 56700 -480 56812 240
rect 57260 -480 57372 240
rect 57820 -480 57932 240
rect 58380 -480 58492 240
rect 58940 -480 59052 240
rect 59500 -480 59612 240
rect 60060 -480 60172 240
rect 60620 -480 60732 240
rect 61180 -480 61292 240
rect 61740 -480 61852 240
rect 62300 -480 62412 240
rect 62860 -480 62972 240
rect 63420 -480 63532 240
rect 63980 -480 64092 240
rect 64540 -480 64652 240
rect 65100 -480 65212 240
rect 65660 -480 65772 240
rect 66220 -480 66332 240
rect 66780 -480 66892 240
rect 67340 -480 67452 240
rect 67900 -480 68012 240
rect 68460 -480 68572 240
rect 69020 -480 69132 240
rect 69580 -480 69692 240
rect 70140 -480 70252 240
rect 70700 -480 70812 240
rect 71260 -480 71372 240
rect 71820 -480 71932 240
rect 72380 -480 72492 240
rect 72940 -480 73052 240
rect 73500 -480 73612 240
rect 74060 -480 74172 240
rect 74620 -480 74732 240
rect 75180 -480 75292 240
rect 75740 -480 75852 240
rect 76300 -480 76412 240
rect 76860 -480 76972 240
rect 77420 -480 77532 240
rect 77980 -480 78092 240
rect 78540 -480 78652 240
rect 79100 -480 79212 240
rect 79660 -480 79772 240
rect 80220 -480 80332 240
rect 80780 -480 80892 240
rect 81340 -480 81452 240
rect 81900 -480 82012 240
rect 82460 -480 82572 240
rect 83020 -480 83132 240
rect 83580 -480 83692 240
rect 84140 -480 84252 240
rect 84700 -480 84812 240
rect 85260 -480 85372 240
rect 85820 -480 85932 240
rect 86380 -480 86492 240
rect 86940 -480 87052 240
rect 87500 -480 87612 240
rect 88060 -480 88172 240
rect 88620 -480 88732 240
rect 89180 -480 89292 240
rect 89740 -480 89852 240
rect 90300 -480 90412 240
rect 90860 -480 90972 240
rect 91420 -480 91532 240
rect 91980 -480 92092 240
rect 92540 -480 92652 240
rect 93100 -480 93212 240
rect 93660 -480 93772 240
rect 94220 -480 94332 240
rect 94780 -480 94892 240
rect 95340 -480 95452 240
rect 95900 -480 96012 240
rect 96460 -480 96572 240
rect 97020 -480 97132 240
rect 97580 -480 97692 240
rect 98140 -480 98252 240
rect 98700 -480 98812 240
rect 99260 -480 99372 240
rect 99820 -480 99932 240
rect 100380 -480 100492 240
rect 100940 -480 101052 240
rect 101500 -480 101612 240
rect 102060 -480 102172 240
rect 102620 -480 102732 240
rect 103180 -480 103292 240
rect 103740 -480 103852 240
rect 104300 -480 104412 240
rect 104860 -480 104972 240
rect 105420 -480 105532 240
rect 105980 -480 106092 240
rect 106540 -480 106652 240
rect 107100 -480 107212 240
rect 107660 -480 107772 240
rect 108220 -480 108332 240
rect 108780 -480 108892 240
rect 109340 -480 109452 240
rect 109900 -480 110012 240
rect 110460 -480 110572 240
rect 111020 -480 111132 240
rect 111580 -480 111692 240
rect 112140 -480 112252 240
rect 112700 -480 112812 240
rect 113260 -480 113372 240
rect 113820 -480 113932 240
rect 114380 -480 114492 240
rect 114940 -480 115052 240
rect 115500 -480 115612 240
rect 116060 -480 116172 240
rect 116620 -480 116732 240
rect 117180 -480 117292 240
rect 117740 -480 117852 240
rect 118300 -480 118412 240
rect 118860 -480 118972 240
rect 119420 -480 119532 240
rect 119980 -480 120092 240
rect 120540 -480 120652 240
rect 121100 -480 121212 240
rect 121660 -480 121772 240
rect 122220 -480 122332 240
rect 122780 -480 122892 240
rect 123340 -480 123452 240
rect 123900 -480 124012 240
rect 124460 -480 124572 240
rect 125020 -480 125132 240
rect 125580 -480 125692 240
rect 126140 -480 126252 240
rect 126700 -480 126812 240
rect 127260 -480 127372 240
rect 127820 -480 127932 240
rect 128380 -480 128492 240
rect 128940 -480 129052 240
rect 129500 -480 129612 240
rect 130060 -480 130172 240
rect 130620 -480 130732 240
rect 131180 -480 131292 240
rect 131740 -480 131852 240
rect 132300 -480 132412 240
rect 132860 -480 132972 240
rect 133420 -480 133532 240
rect 133980 -480 134092 240
rect 134540 -480 134652 240
rect 135100 -480 135212 240
rect 135660 -480 135772 240
rect 136220 -480 136332 240
rect 136780 -480 136892 240
rect 137340 -480 137452 240
rect 137900 -480 138012 240
rect 138460 -480 138572 240
rect 139020 -480 139132 240
rect 139580 -480 139692 240
rect 140140 -480 140252 240
rect 140700 -480 140812 240
rect 141260 -480 141372 240
rect 141820 -480 141932 240
rect 142380 -480 142492 240
rect 142940 -480 143052 240
rect 143500 -480 143612 240
rect 144060 -480 144172 240
rect 144620 -480 144732 240
rect 145180 -480 145292 240
rect 145740 -480 145852 240
rect 146300 -480 146412 240
rect 146860 -480 146972 240
rect 147420 -480 147532 240
rect 147980 -480 148092 240
rect 148540 -480 148652 240
rect 149100 -480 149212 240
rect 149660 -480 149772 240
rect 150220 -480 150332 240
rect 150780 -480 150892 240
rect 151340 -480 151452 240
rect 151900 -480 152012 240
rect 152460 -480 152572 240
rect 153020 -480 153132 240
rect 153580 -480 153692 240
rect 154140 -480 154252 240
rect 154700 -480 154812 240
rect 155260 -480 155372 240
rect 155820 -480 155932 240
rect 156380 -480 156492 240
rect 156940 -480 157052 240
rect 157500 -480 157612 240
rect 158060 -480 158172 240
rect 158620 -480 158732 240
rect 159180 -480 159292 240
rect 159740 -480 159852 240
rect 160300 -480 160412 240
rect 160860 -480 160972 240
rect 161420 -480 161532 240
rect 161980 -480 162092 240
rect 162540 -480 162652 240
rect 163100 -480 163212 240
rect 163660 -480 163772 240
rect 164220 -480 164332 240
rect 164780 -480 164892 240
rect 165340 -480 165452 240
rect 165900 -480 166012 240
rect 166460 -480 166572 240
rect 167020 -480 167132 240
rect 167580 -480 167692 240
rect 168140 -480 168252 240
rect 168700 -480 168812 240
rect 169260 -480 169372 240
rect 169820 -480 169932 240
rect 170380 -480 170492 240
rect 170940 -480 171052 240
rect 171500 -480 171612 240
rect 172060 -480 172172 240
rect 172620 -480 172732 240
rect 173180 -480 173292 240
rect 173740 -480 173852 240
rect 174300 -480 174412 240
rect 174860 -480 174972 240
rect 175420 -480 175532 240
rect 175980 -480 176092 240
rect 176540 -480 176652 240
rect 177100 -480 177212 240
rect 177660 -480 177772 240
rect 178220 -480 178332 240
rect 178780 -480 178892 240
rect 179340 -480 179452 240
rect 179900 -480 180012 240
rect 180460 -480 180572 240
rect 181020 -480 181132 240
rect 181580 -480 181692 240
rect 182140 -480 182252 240
rect 182700 -480 182812 240
rect 183260 -480 183372 240
rect 183820 -480 183932 240
rect 184380 -480 184492 240
rect 184940 -480 185052 240
rect 185500 -480 185612 240
rect 186060 -480 186172 240
rect 186620 -480 186732 240
rect 187180 -480 187292 240
rect 187740 -480 187852 240
rect 188300 -480 188412 240
rect 188860 -480 188972 240
rect 189420 -480 189532 240
rect 189980 -480 190092 240
rect 190540 -480 190652 240
rect 191100 -480 191212 240
rect 191660 -480 191772 240
rect 192220 -480 192332 240
rect 192780 -480 192892 240
rect 193340 -480 193452 240
rect 193900 -480 194012 240
rect 194460 -480 194572 240
rect 195020 -480 195132 240
rect 195580 -480 195692 240
rect 196140 -480 196252 240
rect 196700 -480 196812 240
rect 197260 -480 197372 240
rect 197820 -480 197932 240
rect 198380 -480 198492 240
rect 198940 -480 199052 240
rect 199500 -480 199612 240
rect 200060 -480 200172 240
rect 200620 -480 200732 240
rect 201180 -480 201292 240
rect 201740 -480 201852 240
rect 202300 -480 202412 240
rect 202860 -480 202972 240
rect 203420 -480 203532 240
rect 203980 -480 204092 240
rect 204540 -480 204652 240
rect 205100 -480 205212 240
rect 205660 -480 205772 240
rect 206220 -480 206332 240
rect 206780 -480 206892 240
rect 207340 -480 207452 240
rect 207900 -480 208012 240
rect 208460 -480 208572 240
rect 209020 -480 209132 240
rect 209580 -480 209692 240
rect 210140 -480 210252 240
rect 210700 -480 210812 240
rect 211260 -480 211372 240
rect 211820 -480 211932 240
rect 212380 -480 212492 240
rect 212940 -480 213052 240
rect 213500 -480 213612 240
rect 214060 -480 214172 240
rect 214620 -480 214732 240
rect 215180 -480 215292 240
rect 215740 -480 215852 240
rect 216300 -480 216412 240
rect 216860 -480 216972 240
rect 217420 -480 217532 240
rect 217980 -480 218092 240
rect 218540 -480 218652 240
rect 219100 -480 219212 240
rect 219660 -480 219772 240
rect 220220 -480 220332 240
rect 220780 -480 220892 240
rect 221340 -480 221452 240
rect 221900 -480 222012 240
rect 222460 -480 222572 240
rect 223020 -480 223132 240
rect 223580 -480 223692 240
rect 224140 -480 224252 240
rect 224700 -480 224812 240
rect 225260 -480 225372 240
rect 225820 -480 225932 240
rect 226380 -480 226492 240
rect 226940 -480 227052 240
rect 227500 -480 227612 240
rect 228060 -480 228172 240
rect 228620 -480 228732 240
rect 229180 -480 229292 240
rect 229740 -480 229852 240
rect 230300 -480 230412 240
rect 230860 -480 230972 240
rect 231420 -480 231532 240
rect 231980 -480 232092 240
rect 232540 -480 232652 240
rect 233100 -480 233212 240
rect 233660 -480 233772 240
rect 234220 -480 234332 240
rect 234780 -480 234892 240
rect 235340 -480 235452 240
rect 235900 -480 236012 240
rect 236460 -480 236572 240
rect 237020 -480 237132 240
rect 237580 -480 237692 240
rect 238140 -480 238252 240
rect 238700 -480 238812 240
rect 239260 -480 239372 240
rect 239820 -480 239932 240
rect 240380 -480 240492 240
rect 240940 -480 241052 240
rect 241500 -480 241612 240
rect 242060 -480 242172 240
rect 242620 -480 242732 240
rect 243180 -480 243292 240
rect 243740 -480 243852 240
rect 244300 -480 244412 240
rect 244860 -480 244972 240
rect 245420 -480 245532 240
rect 245980 -480 246092 240
rect 246540 -480 246652 240
rect 247100 -480 247212 240
rect 247660 -480 247772 240
rect 248220 -480 248332 240
rect 248780 -480 248892 240
rect 249340 -480 249452 240
rect 249900 -480 250012 240
rect 250460 -480 250572 240
rect 251020 -480 251132 240
rect 251580 -480 251692 240
rect 252140 -480 252252 240
rect 252700 -480 252812 240
rect 253260 -480 253372 240
rect 253820 -480 253932 240
rect 254380 -480 254492 240
rect 254940 -480 255052 240
rect 255500 -480 255612 240
rect 256060 -480 256172 240
rect 256620 -480 256732 240
rect 257180 -480 257292 240
rect 257740 -480 257852 240
rect 258300 -480 258412 240
rect 258860 -480 258972 240
rect 259420 -480 259532 240
rect 259980 -480 260092 240
rect 260540 -480 260652 240
rect 261100 -480 261212 240
rect 261660 -480 261772 240
rect 262220 -480 262332 240
rect 262780 -480 262892 240
rect 263340 -480 263452 240
rect 263900 -480 264012 240
rect 264460 -480 264572 240
rect 265020 -480 265132 240
rect 265580 -480 265692 240
rect 266140 -480 266252 240
rect 266700 -480 266812 240
rect 267260 -480 267372 240
rect 267820 -480 267932 240
rect 268380 -480 268492 240
rect 268940 -480 269052 240
rect 269500 -480 269612 240
rect 270060 -480 270172 240
rect 270620 -480 270732 240
rect 271180 -480 271292 240
rect 271740 -480 271852 240
rect 272300 -480 272412 240
rect 272860 -480 272972 240
rect 273420 -480 273532 240
rect 273980 -480 274092 240
rect 274540 -480 274652 240
rect 275100 -480 275212 240
rect 275660 -480 275772 240
rect 276220 -480 276332 240
rect 276780 -480 276892 240
rect 277340 -480 277452 240
rect 277900 -480 278012 240
rect 278460 -480 278572 240
rect 279020 -480 279132 240
rect 279580 -480 279692 240
rect 280140 -480 280252 240
rect 280700 -480 280812 240
rect 281260 -480 281372 240
rect 281820 -480 281932 240
rect 282380 -480 282492 240
rect 282940 -480 283052 240
rect 283500 -480 283612 240
rect 284060 -480 284172 240
rect 284620 -480 284732 240
rect 285180 -480 285292 240
rect 285740 -480 285852 240
rect 286300 -480 286412 240
rect 286860 -480 286972 240
rect 287420 -480 287532 240
rect 287980 -480 288092 240
<< obsm2 >>
rect 14 299730 4870 299796
rect 5042 299730 13158 299796
rect 13330 299730 21446 299796
rect 21618 299730 29734 299796
rect 29906 299730 38022 299796
rect 38194 299730 46310 299796
rect 46482 299730 54598 299796
rect 54770 299730 62886 299796
rect 63058 299730 71174 299796
rect 71346 299730 79462 299796
rect 79634 299730 87750 299796
rect 87922 299730 96038 299796
rect 96210 299730 104326 299796
rect 104498 299730 112614 299796
rect 112786 299730 120902 299796
rect 121074 299730 129190 299796
rect 129362 299730 137478 299796
rect 137650 299730 145766 299796
rect 145938 299730 154054 299796
rect 154226 299730 162342 299796
rect 162514 299730 170630 299796
rect 170802 299730 178918 299796
rect 179090 299730 187206 299796
rect 187378 299730 195494 299796
rect 195666 299730 203782 299796
rect 203954 299730 212070 299796
rect 212242 299730 220358 299796
rect 220530 299730 228646 299796
rect 228818 299730 236934 299796
rect 237106 299730 245222 299796
rect 245394 299730 253510 299796
rect 253682 299730 261798 299796
rect 261970 299730 270086 299796
rect 270258 299730 278374 299796
rect 278546 299730 286662 299796
rect 286834 299730 294950 299796
rect 295122 299730 299586 299796
rect 14 270 299586 299730
rect 14 9 11870 270
rect 12042 9 12430 270
rect 12602 9 12990 270
rect 13162 9 13550 270
rect 13722 9 14110 270
rect 14282 9 14670 270
rect 14842 9 15230 270
rect 15402 9 15790 270
rect 15962 9 16350 270
rect 16522 9 16910 270
rect 17082 9 17470 270
rect 17642 9 18030 270
rect 18202 9 18590 270
rect 18762 9 19150 270
rect 19322 9 19710 270
rect 19882 9 20270 270
rect 20442 9 20830 270
rect 21002 9 21390 270
rect 21562 9 21950 270
rect 22122 9 22510 270
rect 22682 9 23070 270
rect 23242 9 23630 270
rect 23802 9 24190 270
rect 24362 9 24750 270
rect 24922 9 25310 270
rect 25482 9 25870 270
rect 26042 9 26430 270
rect 26602 9 26990 270
rect 27162 9 27550 270
rect 27722 9 28110 270
rect 28282 9 28670 270
rect 28842 9 29230 270
rect 29402 9 29790 270
rect 29962 9 30350 270
rect 30522 9 30910 270
rect 31082 9 31470 270
rect 31642 9 32030 270
rect 32202 9 32590 270
rect 32762 9 33150 270
rect 33322 9 33710 270
rect 33882 9 34270 270
rect 34442 9 34830 270
rect 35002 9 35390 270
rect 35562 9 35950 270
rect 36122 9 36510 270
rect 36682 9 37070 270
rect 37242 9 37630 270
rect 37802 9 38190 270
rect 38362 9 38750 270
rect 38922 9 39310 270
rect 39482 9 39870 270
rect 40042 9 40430 270
rect 40602 9 40990 270
rect 41162 9 41550 270
rect 41722 9 42110 270
rect 42282 9 42670 270
rect 42842 9 43230 270
rect 43402 9 43790 270
rect 43962 9 44350 270
rect 44522 9 44910 270
rect 45082 9 45470 270
rect 45642 9 46030 270
rect 46202 9 46590 270
rect 46762 9 47150 270
rect 47322 9 47710 270
rect 47882 9 48270 270
rect 48442 9 48830 270
rect 49002 9 49390 270
rect 49562 9 49950 270
rect 50122 9 50510 270
rect 50682 9 51070 270
rect 51242 9 51630 270
rect 51802 9 52190 270
rect 52362 9 52750 270
rect 52922 9 53310 270
rect 53482 9 53870 270
rect 54042 9 54430 270
rect 54602 9 54990 270
rect 55162 9 55550 270
rect 55722 9 56110 270
rect 56282 9 56670 270
rect 56842 9 57230 270
rect 57402 9 57790 270
rect 57962 9 58350 270
rect 58522 9 58910 270
rect 59082 9 59470 270
rect 59642 9 60030 270
rect 60202 9 60590 270
rect 60762 9 61150 270
rect 61322 9 61710 270
rect 61882 9 62270 270
rect 62442 9 62830 270
rect 63002 9 63390 270
rect 63562 9 63950 270
rect 64122 9 64510 270
rect 64682 9 65070 270
rect 65242 9 65630 270
rect 65802 9 66190 270
rect 66362 9 66750 270
rect 66922 9 67310 270
rect 67482 9 67870 270
rect 68042 9 68430 270
rect 68602 9 68990 270
rect 69162 9 69550 270
rect 69722 9 70110 270
rect 70282 9 70670 270
rect 70842 9 71230 270
rect 71402 9 71790 270
rect 71962 9 72350 270
rect 72522 9 72910 270
rect 73082 9 73470 270
rect 73642 9 74030 270
rect 74202 9 74590 270
rect 74762 9 75150 270
rect 75322 9 75710 270
rect 75882 9 76270 270
rect 76442 9 76830 270
rect 77002 9 77390 270
rect 77562 9 77950 270
rect 78122 9 78510 270
rect 78682 9 79070 270
rect 79242 9 79630 270
rect 79802 9 80190 270
rect 80362 9 80750 270
rect 80922 9 81310 270
rect 81482 9 81870 270
rect 82042 9 82430 270
rect 82602 9 82990 270
rect 83162 9 83550 270
rect 83722 9 84110 270
rect 84282 9 84670 270
rect 84842 9 85230 270
rect 85402 9 85790 270
rect 85962 9 86350 270
rect 86522 9 86910 270
rect 87082 9 87470 270
rect 87642 9 88030 270
rect 88202 9 88590 270
rect 88762 9 89150 270
rect 89322 9 89710 270
rect 89882 9 90270 270
rect 90442 9 90830 270
rect 91002 9 91390 270
rect 91562 9 91950 270
rect 92122 9 92510 270
rect 92682 9 93070 270
rect 93242 9 93630 270
rect 93802 9 94190 270
rect 94362 9 94750 270
rect 94922 9 95310 270
rect 95482 9 95870 270
rect 96042 9 96430 270
rect 96602 9 96990 270
rect 97162 9 97550 270
rect 97722 9 98110 270
rect 98282 9 98670 270
rect 98842 9 99230 270
rect 99402 9 99790 270
rect 99962 9 100350 270
rect 100522 9 100910 270
rect 101082 9 101470 270
rect 101642 9 102030 270
rect 102202 9 102590 270
rect 102762 9 103150 270
rect 103322 9 103710 270
rect 103882 9 104270 270
rect 104442 9 104830 270
rect 105002 9 105390 270
rect 105562 9 105950 270
rect 106122 9 106510 270
rect 106682 9 107070 270
rect 107242 9 107630 270
rect 107802 9 108190 270
rect 108362 9 108750 270
rect 108922 9 109310 270
rect 109482 9 109870 270
rect 110042 9 110430 270
rect 110602 9 110990 270
rect 111162 9 111550 270
rect 111722 9 112110 270
rect 112282 9 112670 270
rect 112842 9 113230 270
rect 113402 9 113790 270
rect 113962 9 114350 270
rect 114522 9 114910 270
rect 115082 9 115470 270
rect 115642 9 116030 270
rect 116202 9 116590 270
rect 116762 9 117150 270
rect 117322 9 117710 270
rect 117882 9 118270 270
rect 118442 9 118830 270
rect 119002 9 119390 270
rect 119562 9 119950 270
rect 120122 9 120510 270
rect 120682 9 121070 270
rect 121242 9 121630 270
rect 121802 9 122190 270
rect 122362 9 122750 270
rect 122922 9 123310 270
rect 123482 9 123870 270
rect 124042 9 124430 270
rect 124602 9 124990 270
rect 125162 9 125550 270
rect 125722 9 126110 270
rect 126282 9 126670 270
rect 126842 9 127230 270
rect 127402 9 127790 270
rect 127962 9 128350 270
rect 128522 9 128910 270
rect 129082 9 129470 270
rect 129642 9 130030 270
rect 130202 9 130590 270
rect 130762 9 131150 270
rect 131322 9 131710 270
rect 131882 9 132270 270
rect 132442 9 132830 270
rect 133002 9 133390 270
rect 133562 9 133950 270
rect 134122 9 134510 270
rect 134682 9 135070 270
rect 135242 9 135630 270
rect 135802 9 136190 270
rect 136362 9 136750 270
rect 136922 9 137310 270
rect 137482 9 137870 270
rect 138042 9 138430 270
rect 138602 9 138990 270
rect 139162 9 139550 270
rect 139722 9 140110 270
rect 140282 9 140670 270
rect 140842 9 141230 270
rect 141402 9 141790 270
rect 141962 9 142350 270
rect 142522 9 142910 270
rect 143082 9 143470 270
rect 143642 9 144030 270
rect 144202 9 144590 270
rect 144762 9 145150 270
rect 145322 9 145710 270
rect 145882 9 146270 270
rect 146442 9 146830 270
rect 147002 9 147390 270
rect 147562 9 147950 270
rect 148122 9 148510 270
rect 148682 9 149070 270
rect 149242 9 149630 270
rect 149802 9 150190 270
rect 150362 9 150750 270
rect 150922 9 151310 270
rect 151482 9 151870 270
rect 152042 9 152430 270
rect 152602 9 152990 270
rect 153162 9 153550 270
rect 153722 9 154110 270
rect 154282 9 154670 270
rect 154842 9 155230 270
rect 155402 9 155790 270
rect 155962 9 156350 270
rect 156522 9 156910 270
rect 157082 9 157470 270
rect 157642 9 158030 270
rect 158202 9 158590 270
rect 158762 9 159150 270
rect 159322 9 159710 270
rect 159882 9 160270 270
rect 160442 9 160830 270
rect 161002 9 161390 270
rect 161562 9 161950 270
rect 162122 9 162510 270
rect 162682 9 163070 270
rect 163242 9 163630 270
rect 163802 9 164190 270
rect 164362 9 164750 270
rect 164922 9 165310 270
rect 165482 9 165870 270
rect 166042 9 166430 270
rect 166602 9 166990 270
rect 167162 9 167550 270
rect 167722 9 168110 270
rect 168282 9 168670 270
rect 168842 9 169230 270
rect 169402 9 169790 270
rect 169962 9 170350 270
rect 170522 9 170910 270
rect 171082 9 171470 270
rect 171642 9 172030 270
rect 172202 9 172590 270
rect 172762 9 173150 270
rect 173322 9 173710 270
rect 173882 9 174270 270
rect 174442 9 174830 270
rect 175002 9 175390 270
rect 175562 9 175950 270
rect 176122 9 176510 270
rect 176682 9 177070 270
rect 177242 9 177630 270
rect 177802 9 178190 270
rect 178362 9 178750 270
rect 178922 9 179310 270
rect 179482 9 179870 270
rect 180042 9 180430 270
rect 180602 9 180990 270
rect 181162 9 181550 270
rect 181722 9 182110 270
rect 182282 9 182670 270
rect 182842 9 183230 270
rect 183402 9 183790 270
rect 183962 9 184350 270
rect 184522 9 184910 270
rect 185082 9 185470 270
rect 185642 9 186030 270
rect 186202 9 186590 270
rect 186762 9 187150 270
rect 187322 9 187710 270
rect 187882 9 188270 270
rect 188442 9 188830 270
rect 189002 9 189390 270
rect 189562 9 189950 270
rect 190122 9 190510 270
rect 190682 9 191070 270
rect 191242 9 191630 270
rect 191802 9 192190 270
rect 192362 9 192750 270
rect 192922 9 193310 270
rect 193482 9 193870 270
rect 194042 9 194430 270
rect 194602 9 194990 270
rect 195162 9 195550 270
rect 195722 9 196110 270
rect 196282 9 196670 270
rect 196842 9 197230 270
rect 197402 9 197790 270
rect 197962 9 198350 270
rect 198522 9 198910 270
rect 199082 9 199470 270
rect 199642 9 200030 270
rect 200202 9 200590 270
rect 200762 9 201150 270
rect 201322 9 201710 270
rect 201882 9 202270 270
rect 202442 9 202830 270
rect 203002 9 203390 270
rect 203562 9 203950 270
rect 204122 9 204510 270
rect 204682 9 205070 270
rect 205242 9 205630 270
rect 205802 9 206190 270
rect 206362 9 206750 270
rect 206922 9 207310 270
rect 207482 9 207870 270
rect 208042 9 208430 270
rect 208602 9 208990 270
rect 209162 9 209550 270
rect 209722 9 210110 270
rect 210282 9 210670 270
rect 210842 9 211230 270
rect 211402 9 211790 270
rect 211962 9 212350 270
rect 212522 9 212910 270
rect 213082 9 213470 270
rect 213642 9 214030 270
rect 214202 9 214590 270
rect 214762 9 215150 270
rect 215322 9 215710 270
rect 215882 9 216270 270
rect 216442 9 216830 270
rect 217002 9 217390 270
rect 217562 9 217950 270
rect 218122 9 218510 270
rect 218682 9 219070 270
rect 219242 9 219630 270
rect 219802 9 220190 270
rect 220362 9 220750 270
rect 220922 9 221310 270
rect 221482 9 221870 270
rect 222042 9 222430 270
rect 222602 9 222990 270
rect 223162 9 223550 270
rect 223722 9 224110 270
rect 224282 9 224670 270
rect 224842 9 225230 270
rect 225402 9 225790 270
rect 225962 9 226350 270
rect 226522 9 226910 270
rect 227082 9 227470 270
rect 227642 9 228030 270
rect 228202 9 228590 270
rect 228762 9 229150 270
rect 229322 9 229710 270
rect 229882 9 230270 270
rect 230442 9 230830 270
rect 231002 9 231390 270
rect 231562 9 231950 270
rect 232122 9 232510 270
rect 232682 9 233070 270
rect 233242 9 233630 270
rect 233802 9 234190 270
rect 234362 9 234750 270
rect 234922 9 235310 270
rect 235482 9 235870 270
rect 236042 9 236430 270
rect 236602 9 236990 270
rect 237162 9 237550 270
rect 237722 9 238110 270
rect 238282 9 238670 270
rect 238842 9 239230 270
rect 239402 9 239790 270
rect 239962 9 240350 270
rect 240522 9 240910 270
rect 241082 9 241470 270
rect 241642 9 242030 270
rect 242202 9 242590 270
rect 242762 9 243150 270
rect 243322 9 243710 270
rect 243882 9 244270 270
rect 244442 9 244830 270
rect 245002 9 245390 270
rect 245562 9 245950 270
rect 246122 9 246510 270
rect 246682 9 247070 270
rect 247242 9 247630 270
rect 247802 9 248190 270
rect 248362 9 248750 270
rect 248922 9 249310 270
rect 249482 9 249870 270
rect 250042 9 250430 270
rect 250602 9 250990 270
rect 251162 9 251550 270
rect 251722 9 252110 270
rect 252282 9 252670 270
rect 252842 9 253230 270
rect 253402 9 253790 270
rect 253962 9 254350 270
rect 254522 9 254910 270
rect 255082 9 255470 270
rect 255642 9 256030 270
rect 256202 9 256590 270
rect 256762 9 257150 270
rect 257322 9 257710 270
rect 257882 9 258270 270
rect 258442 9 258830 270
rect 259002 9 259390 270
rect 259562 9 259950 270
rect 260122 9 260510 270
rect 260682 9 261070 270
rect 261242 9 261630 270
rect 261802 9 262190 270
rect 262362 9 262750 270
rect 262922 9 263310 270
rect 263482 9 263870 270
rect 264042 9 264430 270
rect 264602 9 264990 270
rect 265162 9 265550 270
rect 265722 9 266110 270
rect 266282 9 266670 270
rect 266842 9 267230 270
rect 267402 9 267790 270
rect 267962 9 268350 270
rect 268522 9 268910 270
rect 269082 9 269470 270
rect 269642 9 270030 270
rect 270202 9 270590 270
rect 270762 9 271150 270
rect 271322 9 271710 270
rect 271882 9 272270 270
rect 272442 9 272830 270
rect 273002 9 273390 270
rect 273562 9 273950 270
rect 274122 9 274510 270
rect 274682 9 275070 270
rect 275242 9 275630 270
rect 275802 9 276190 270
rect 276362 9 276750 270
rect 276922 9 277310 270
rect 277482 9 277870 270
rect 278042 9 278430 270
rect 278602 9 278990 270
rect 279162 9 279550 270
rect 279722 9 280110 270
rect 280282 9 280670 270
rect 280842 9 281230 270
rect 281402 9 281790 270
rect 281962 9 282350 270
rect 282522 9 282910 270
rect 283082 9 283470 270
rect 283642 9 284030 270
rect 284202 9 284590 270
rect 284762 9 285150 270
rect 285322 9 285710 270
rect 285882 9 286270 270
rect 286442 9 286830 270
rect 287002 9 287390 270
rect 287562 9 287950 270
rect 288122 9 299586 270
<< metal3 >>
rect 299760 296996 300480 297108
rect -480 296828 240 296940
rect -480 291284 240 291396
rect 299760 291340 300480 291452
rect -480 285740 240 285852
rect 299760 285684 300480 285796
rect -480 280196 240 280308
rect 299760 280028 300480 280140
rect -480 274652 240 274764
rect 299760 274372 300480 274484
rect -480 269108 240 269220
rect 299760 268716 300480 268828
rect -480 263564 240 263676
rect 299760 263060 300480 263172
rect -480 258020 240 258132
rect 299760 257404 300480 257516
rect -480 252476 240 252588
rect 299760 251748 300480 251860
rect -480 246932 240 247044
rect 299760 246092 300480 246204
rect -480 241388 240 241500
rect 299760 240436 300480 240548
rect -480 235844 240 235956
rect 299760 234780 300480 234892
rect -480 230300 240 230412
rect 299760 229124 300480 229236
rect -480 224756 240 224868
rect 299760 223468 300480 223580
rect -480 219212 240 219324
rect 299760 217812 300480 217924
rect -480 213668 240 213780
rect 299760 212156 300480 212268
rect -480 208124 240 208236
rect 299760 206500 300480 206612
rect -480 202580 240 202692
rect 299760 200844 300480 200956
rect -480 197036 240 197148
rect 299760 195188 300480 195300
rect -480 191492 240 191604
rect 299760 189532 300480 189644
rect -480 185948 240 186060
rect 299760 183876 300480 183988
rect -480 180404 240 180516
rect 299760 178220 300480 178332
rect -480 174860 240 174972
rect 299760 172564 300480 172676
rect -480 169316 240 169428
rect 299760 166908 300480 167020
rect -480 163772 240 163884
rect 299760 161252 300480 161364
rect -480 158228 240 158340
rect 299760 155596 300480 155708
rect -480 152684 240 152796
rect 299760 149940 300480 150052
rect -480 147140 240 147252
rect 299760 144284 300480 144396
rect -480 141596 240 141708
rect 299760 138628 300480 138740
rect -480 136052 240 136164
rect 299760 132972 300480 133084
rect -480 130508 240 130620
rect 299760 127316 300480 127428
rect -480 124964 240 125076
rect 299760 121660 300480 121772
rect -480 119420 240 119532
rect 299760 116004 300480 116116
rect -480 113876 240 113988
rect 299760 110348 300480 110460
rect -480 108332 240 108444
rect 299760 104692 300480 104804
rect -480 102788 240 102900
rect 299760 99036 300480 99148
rect -480 97244 240 97356
rect 299760 93380 300480 93492
rect -480 91700 240 91812
rect 299760 87724 300480 87836
rect -480 86156 240 86268
rect 299760 82068 300480 82180
rect -480 80612 240 80724
rect 299760 76412 300480 76524
rect -480 75068 240 75180
rect 299760 70756 300480 70868
rect -480 69524 240 69636
rect 299760 65100 300480 65212
rect -480 63980 240 64092
rect 299760 59444 300480 59556
rect -480 58436 240 58548
rect 299760 53788 300480 53900
rect -480 52892 240 53004
rect 299760 48132 300480 48244
rect -480 47348 240 47460
rect 299760 42476 300480 42588
rect -480 41804 240 41916
rect 299760 36820 300480 36932
rect -480 36260 240 36372
rect 299760 31164 300480 31276
rect -480 30716 240 30828
rect 299760 25508 300480 25620
rect -480 25172 240 25284
rect 299760 19852 300480 19964
rect -480 19628 240 19740
rect -480 14084 240 14196
rect 299760 14196 300480 14308
rect -480 8540 240 8652
rect 299760 8540 300480 8652
rect -480 2996 240 3108
rect 299760 2884 300480 2996
<< obsm3 >>
rect 9 297138 299796 298018
rect 9 296970 299730 297138
rect 270 296966 299730 296970
rect 270 296798 299796 296966
rect 9 291482 299796 296798
rect 9 291426 299730 291482
rect 270 291310 299730 291426
rect 270 291254 299796 291310
rect 9 285882 299796 291254
rect 270 285826 299796 285882
rect 270 285710 299730 285826
rect 9 285654 299730 285710
rect 9 280338 299796 285654
rect 270 280170 299796 280338
rect 270 280166 299730 280170
rect 9 279998 299730 280166
rect 9 274794 299796 279998
rect 270 274622 299796 274794
rect 9 274514 299796 274622
rect 9 274342 299730 274514
rect 9 269250 299796 274342
rect 270 269078 299796 269250
rect 9 268858 299796 269078
rect 9 268686 299730 268858
rect 9 263706 299796 268686
rect 270 263534 299796 263706
rect 9 263202 299796 263534
rect 9 263030 299730 263202
rect 9 258162 299796 263030
rect 270 257990 299796 258162
rect 9 257546 299796 257990
rect 9 257374 299730 257546
rect 9 252618 299796 257374
rect 270 252446 299796 252618
rect 9 251890 299796 252446
rect 9 251718 299730 251890
rect 9 247074 299796 251718
rect 270 246902 299796 247074
rect 9 246234 299796 246902
rect 9 246062 299730 246234
rect 9 241530 299796 246062
rect 270 241358 299796 241530
rect 9 240578 299796 241358
rect 9 240406 299730 240578
rect 9 235986 299796 240406
rect 270 235814 299796 235986
rect 9 234922 299796 235814
rect 9 234750 299730 234922
rect 9 230442 299796 234750
rect 270 230270 299796 230442
rect 9 229266 299796 230270
rect 9 229094 299730 229266
rect 9 224898 299796 229094
rect 270 224726 299796 224898
rect 9 223610 299796 224726
rect 9 223438 299730 223610
rect 9 219354 299796 223438
rect 270 219182 299796 219354
rect 9 217954 299796 219182
rect 9 217782 299730 217954
rect 9 213810 299796 217782
rect 270 213638 299796 213810
rect 9 212298 299796 213638
rect 9 212126 299730 212298
rect 9 208266 299796 212126
rect 270 208094 299796 208266
rect 9 206642 299796 208094
rect 9 206470 299730 206642
rect 9 202722 299796 206470
rect 270 202550 299796 202722
rect 9 200986 299796 202550
rect 9 200814 299730 200986
rect 9 197178 299796 200814
rect 270 197006 299796 197178
rect 9 195330 299796 197006
rect 9 195158 299730 195330
rect 9 191634 299796 195158
rect 270 191462 299796 191634
rect 9 189674 299796 191462
rect 9 189502 299730 189674
rect 9 186090 299796 189502
rect 270 185918 299796 186090
rect 9 184018 299796 185918
rect 9 183846 299730 184018
rect 9 180546 299796 183846
rect 270 180374 299796 180546
rect 9 178362 299796 180374
rect 9 178190 299730 178362
rect 9 175002 299796 178190
rect 270 174830 299796 175002
rect 9 172706 299796 174830
rect 9 172534 299730 172706
rect 9 169458 299796 172534
rect 270 169286 299796 169458
rect 9 167050 299796 169286
rect 9 166878 299730 167050
rect 9 163914 299796 166878
rect 270 163742 299796 163914
rect 9 161394 299796 163742
rect 9 161222 299730 161394
rect 9 158370 299796 161222
rect 270 158198 299796 158370
rect 9 155738 299796 158198
rect 9 155566 299730 155738
rect 9 152826 299796 155566
rect 270 152654 299796 152826
rect 9 150082 299796 152654
rect 9 149910 299730 150082
rect 9 147282 299796 149910
rect 270 147110 299796 147282
rect 9 144426 299796 147110
rect 9 144254 299730 144426
rect 9 141738 299796 144254
rect 270 141566 299796 141738
rect 9 138770 299796 141566
rect 9 138598 299730 138770
rect 9 136194 299796 138598
rect 270 136022 299796 136194
rect 9 133114 299796 136022
rect 9 132942 299730 133114
rect 9 130650 299796 132942
rect 270 130478 299796 130650
rect 9 127458 299796 130478
rect 9 127286 299730 127458
rect 9 125106 299796 127286
rect 270 124934 299796 125106
rect 9 121802 299796 124934
rect 9 121630 299730 121802
rect 9 119562 299796 121630
rect 270 119390 299796 119562
rect 9 116146 299796 119390
rect 9 115974 299730 116146
rect 9 114018 299796 115974
rect 270 113846 299796 114018
rect 9 110490 299796 113846
rect 9 110318 299730 110490
rect 9 108474 299796 110318
rect 270 108302 299796 108474
rect 9 104834 299796 108302
rect 9 104662 299730 104834
rect 9 102930 299796 104662
rect 270 102758 299796 102930
rect 9 99178 299796 102758
rect 9 99006 299730 99178
rect 9 97386 299796 99006
rect 270 97214 299796 97386
rect 9 93522 299796 97214
rect 9 93350 299730 93522
rect 9 91842 299796 93350
rect 270 91670 299796 91842
rect 9 87866 299796 91670
rect 9 87694 299730 87866
rect 9 86298 299796 87694
rect 270 86126 299796 86298
rect 9 82210 299796 86126
rect 9 82038 299730 82210
rect 9 80754 299796 82038
rect 270 80582 299796 80754
rect 9 76554 299796 80582
rect 9 76382 299730 76554
rect 9 75210 299796 76382
rect 270 75038 299796 75210
rect 9 70898 299796 75038
rect 9 70726 299730 70898
rect 9 69666 299796 70726
rect 270 69494 299796 69666
rect 9 65242 299796 69494
rect 9 65070 299730 65242
rect 9 64122 299796 65070
rect 270 63950 299796 64122
rect 9 59586 299796 63950
rect 9 59414 299730 59586
rect 9 58578 299796 59414
rect 270 58406 299796 58578
rect 9 53930 299796 58406
rect 9 53758 299730 53930
rect 9 53034 299796 53758
rect 270 52862 299796 53034
rect 9 48274 299796 52862
rect 9 48102 299730 48274
rect 9 47490 299796 48102
rect 270 47318 299796 47490
rect 9 42618 299796 47318
rect 9 42446 299730 42618
rect 9 41946 299796 42446
rect 270 41774 299796 41946
rect 9 36962 299796 41774
rect 9 36790 299730 36962
rect 9 36402 299796 36790
rect 270 36230 299796 36402
rect 9 31306 299796 36230
rect 9 31134 299730 31306
rect 9 30858 299796 31134
rect 270 30686 299796 30858
rect 9 25650 299796 30686
rect 9 25478 299730 25650
rect 9 25314 299796 25478
rect 270 25142 299796 25314
rect 9 19994 299796 25142
rect 9 19822 299730 19994
rect 9 19770 299796 19822
rect 270 19598 299796 19770
rect 9 14338 299796 19598
rect 9 14226 299730 14338
rect 270 14166 299730 14226
rect 270 14054 299796 14166
rect 9 8682 299796 14054
rect 270 8510 299730 8682
rect 9 3138 299796 8510
rect 270 3026 299796 3138
rect 270 2966 299730 3026
rect 9 2854 299730 2966
rect 9 14 299796 2854
<< metal4 >>
rect -4243 -3347 -3933 303227
rect -3763 -2867 -3453 302747
rect -3283 -2387 -2973 302267
rect -2803 -1907 -2493 301787
rect -2323 -1427 -2013 301307
rect -1843 -947 -1533 300827
rect -1363 -467 -1053 300347
rect -883 13 -573 299867
rect 1017 -3347 1327 303227
rect 2877 -3347 3187 303227
rect 4737 -3347 5047 303227
rect 6597 -3347 6907 303227
rect 8457 -3347 8767 303227
rect 10317 -3347 10627 303227
rect 20877 291987 21187 303227
rect 22737 291987 23047 303227
rect 24597 291987 24907 303227
rect 26457 291987 26767 303227
rect 38877 291987 39187 303227
rect 40737 291987 41047 303227
rect 42597 291987 42907 303227
rect 44457 291987 44767 303227
rect 56877 291987 57187 303227
rect 58737 291987 59047 303227
rect 60597 291987 60907 303227
rect 62457 291987 62767 303227
rect 74877 291987 75187 303227
rect 76737 291987 77047 303227
rect 78597 291987 78907 303227
rect 80457 291987 80767 303227
rect 92877 291987 93187 303227
rect 94737 291987 95047 303227
rect 96597 291987 96907 303227
rect 19017 216987 19327 224429
rect 20877 216987 21187 224429
rect 22737 216987 23047 224429
rect 37017 216987 37327 224429
rect 38877 216987 39187 224429
rect 40737 216987 41047 224429
rect 55017 216987 55327 224429
rect 56877 216987 57187 224429
rect 58737 216987 59047 224429
rect 73017 216987 73327 224429
rect 74877 216987 75187 224429
rect 76737 216987 77047 224429
rect 91017 216987 91327 224429
rect 92877 216987 93187 224429
rect 94737 216987 95047 224429
rect 19017 144487 19327 149429
rect 20877 144487 21187 149429
rect 37017 144487 37327 149429
rect 38877 144487 39187 149429
rect 55017 144487 55327 149429
rect 56877 144487 57187 149429
rect 73017 144487 73327 149429
rect 74877 144487 75187 149429
rect 91017 144487 91327 149429
rect 92877 144487 93187 149429
rect 12177 -3347 12487 76929
rect 14037 -3347 14347 76929
rect 19017 26175 19327 76929
rect 20877 26175 21187 76929
rect 22737 26175 23047 76929
rect 24597 26175 24907 76929
rect 26457 26175 26767 76929
rect 28317 26175 28627 76929
rect 30177 26175 30487 76929
rect 32037 26175 32347 76929
rect 37017 26175 37327 76929
rect 38877 26175 39187 76929
rect 40737 26175 41047 76929
rect 42597 26175 42907 76929
rect 44457 26175 44767 76929
rect 46317 26175 46627 76929
rect 48177 52751 48487 76929
rect 48177 26175 48487 50209
rect 50037 26175 50347 76929
rect 55017 26175 55327 76929
rect 56877 26175 57187 76929
rect 58737 26175 59047 76929
rect 60597 26175 60907 76929
rect 62457 26175 62767 76929
rect 64317 26175 64627 76929
rect 66177 26175 66487 76929
rect 68037 26175 68347 76929
rect 73017 26175 73327 76929
rect 19017 -3347 19327 6217
rect 20877 -3347 21187 6217
rect 22737 -3347 23047 6217
rect 37017 -3347 37327 6217
rect 38877 -3347 39187 6217
rect 40737 -3347 41047 6217
rect 55017 -3347 55327 6217
rect 56877 -3347 57187 6217
rect 58737 -3347 59047 6217
rect 73017 -3347 73327 6217
rect 74877 -3347 75187 76929
rect 76737 -3347 77047 76929
rect 78597 -3347 78907 76929
rect 80457 -3347 80767 76929
rect 82317 -3347 82627 76929
rect 84177 -3347 84487 76929
rect 86037 -3347 86347 76929
rect 91017 -3347 91327 76929
rect 92877 -3347 93187 76929
rect 94737 -3347 95047 76929
rect 96597 -3347 96907 76929
rect 98457 -3347 98767 303227
rect 100317 -3347 100627 303227
rect 102177 -3347 102487 303227
rect 104037 -3347 104347 303227
rect 110877 291987 111187 303227
rect 112737 291987 113047 303227
rect 114597 291987 114907 303227
rect 116457 291987 116767 303227
rect 128877 291987 129187 303227
rect 130737 291987 131047 303227
rect 132597 291987 132907 303227
rect 134457 291987 134767 303227
rect 146877 291987 147187 303227
rect 148737 291987 149047 303227
rect 150597 291987 150907 303227
rect 152457 291987 152767 303227
rect 164877 291987 165187 303227
rect 166737 291987 167047 303227
rect 168597 291987 168907 303227
rect 170457 291987 170767 303227
rect 182877 291987 183187 303227
rect 184737 291987 185047 303227
rect 186597 291987 186907 303227
rect 188457 291987 188767 303227
rect 109017 216987 109327 224429
rect 110877 216987 111187 224429
rect 112737 216987 113047 224429
rect 127017 216987 127327 224429
rect 128877 216987 129187 224429
rect 130737 216987 131047 224429
rect 145017 216987 145327 224429
rect 146877 216987 147187 224429
rect 148737 216987 149047 224429
rect 163017 216987 163327 224429
rect 164877 216987 165187 224429
rect 166737 216987 167047 224429
rect 181017 216987 181327 224429
rect 182877 216987 183187 224429
rect 184737 216987 185047 224429
rect 109017 144487 109327 149429
rect 110877 144487 111187 149429
rect 127017 144487 127327 149429
rect 128877 144487 129187 149429
rect 145017 144487 145327 149429
rect 146877 144487 147187 149429
rect 163017 144487 163327 149429
rect 164877 144487 165187 149429
rect 181017 144487 181327 149429
rect 182877 144487 183187 149429
rect 109017 -3347 109327 76929
rect 110877 -3347 111187 76929
rect 112737 -3347 113047 76929
rect 114597 -3347 114907 76929
rect 116457 -3347 116767 76929
rect 118317 -3347 118627 76929
rect 120177 -3347 120487 76929
rect 127017 71987 127327 76929
rect 128877 71987 129187 76929
rect 145017 71987 145327 76929
rect 146877 71987 147187 76929
rect 163017 71987 163327 76929
rect 164877 71987 165187 76929
rect 181017 71987 181327 76929
rect 182877 71987 183187 76929
rect 194037 71987 194347 303227
rect 199017 71987 199327 303227
rect 200877 71987 201187 303227
rect 202737 71987 203047 303227
rect 204597 71987 204907 303227
rect 206457 71987 206767 303227
rect 218877 291987 219187 303227
rect 220737 291987 221047 303227
rect 222597 291987 222907 303227
rect 224457 291987 224767 303227
rect 236877 291987 237187 303227
rect 238737 291987 239047 303227
rect 240597 291987 240907 303227
rect 242457 291987 242767 303227
rect 254877 291987 255187 303227
rect 256737 291987 257047 303227
rect 258597 291987 258907 303227
rect 260457 291987 260767 303227
rect 272877 291987 273187 303227
rect 274737 291987 275047 303227
rect 276597 291987 276907 303227
rect 278457 291987 278767 303227
rect 290877 291987 291187 303227
rect 217017 216987 217327 224429
rect 218877 216987 219187 224429
rect 220737 216987 221047 224429
rect 235017 216987 235327 224429
rect 236877 216987 237187 224429
rect 238737 216987 239047 224429
rect 253017 216987 253327 224429
rect 254877 216987 255187 224429
rect 256737 216987 257047 224429
rect 271017 216987 271327 224429
rect 272877 216987 273187 224429
rect 274737 216987 275047 224429
rect 289017 216987 289327 224429
rect 290877 216987 291187 224429
rect 217017 144487 217327 149429
rect 218877 144487 219187 149429
rect 235017 144487 235327 149429
rect 236877 144487 237187 149429
rect 253017 144487 253327 149429
rect 254877 144487 255187 149429
rect 271017 144487 271327 149429
rect 272877 144487 273187 149429
rect 289017 144487 289327 149429
rect 290877 144487 291187 149429
rect 127017 -3347 127327 4429
rect 128877 -3347 129187 4429
rect 145017 -3347 145327 4429
rect 146877 -3347 147187 4429
rect 163017 -3347 163327 4429
rect 164877 -3347 165187 4429
rect 181017 -3347 181327 4429
rect 182877 -3347 183187 4429
rect 199017 -3347 199327 4429
rect 200877 -3347 201187 4429
rect 208317 -3347 208627 76929
rect 210177 -3347 210487 76929
rect 212037 -3347 212347 76929
rect 217017 -3347 217327 76929
rect 218877 -3347 219187 76929
rect 220737 -3347 221047 76929
rect 222597 -3347 222907 76929
rect 224457 -3347 224767 76929
rect 226317 -3347 226627 76929
rect 228177 -3347 228487 76929
rect 230037 -3347 230347 76929
rect 235017 -3347 235327 76929
rect 236877 -3347 237187 76929
rect 238737 -3347 239047 76929
rect 240597 -3347 240907 76929
rect 242457 -3347 242767 76929
rect 244317 -3347 244627 76929
rect 246177 -3347 246487 76929
rect 248037 -3347 248347 76929
rect 253017 -3347 253327 76929
rect 254877 -3347 255187 76929
rect 256737 -3347 257047 76929
rect 258597 -3347 258907 76929
rect 260457 -3347 260767 76929
rect 262317 -3347 262627 76929
rect 264177 -3347 264487 76929
rect 266037 -3347 266347 76929
rect 271017 -3347 271327 76929
rect 272877 -3347 273187 76929
rect 274737 -3347 275047 76929
rect 276597 -3347 276907 76929
rect 278457 -3347 278767 76929
rect 280317 -3347 280627 76929
rect 282177 -3347 282487 76929
rect 284037 -3347 284347 76929
rect 289017 -3347 289327 76929
rect 290877 -3347 291187 76929
rect 292737 -3347 293047 303227
rect 294597 -3347 294907 303227
rect 296457 -3347 296767 303227
rect 298317 -3347 298627 303227
rect 300565 13 300875 299867
rect 301045 -467 301355 300347
rect 301525 -947 301835 300827
rect 302005 -1427 302315 301307
rect 302485 -1907 302795 301787
rect 302965 -2387 303275 302267
rect 303445 -2867 303755 302747
rect 303925 -3347 304235 303227
<< obsm4 >>
rect 2702 345 2847 297855
rect 3217 345 4707 297855
rect 5077 345 6567 297855
rect 6937 345 8427 297855
rect 8797 345 10287 297855
rect 10657 291957 20847 297855
rect 21217 291957 22707 297855
rect 23077 291957 24567 297855
rect 24937 291957 26427 297855
rect 26797 291957 38847 297855
rect 39217 291957 40707 297855
rect 41077 291957 42567 297855
rect 42937 291957 44427 297855
rect 44797 291957 56847 297855
rect 57217 291957 58707 297855
rect 59077 291957 60567 297855
rect 60937 291957 62427 297855
rect 62797 291957 74847 297855
rect 75217 291957 76707 297855
rect 77077 291957 78567 297855
rect 78937 291957 80427 297855
rect 80797 291957 92847 297855
rect 93217 291957 94707 297855
rect 95077 291957 96567 297855
rect 96937 291957 98427 297855
rect 10657 224459 98427 291957
rect 10657 216957 18987 224459
rect 19357 216957 20847 224459
rect 21217 216957 22707 224459
rect 23077 216957 36987 224459
rect 37357 216957 38847 224459
rect 39217 216957 40707 224459
rect 41077 216957 54987 224459
rect 55357 216957 56847 224459
rect 57217 216957 58707 224459
rect 59077 216957 72987 224459
rect 73357 216957 74847 224459
rect 75217 216957 76707 224459
rect 77077 216957 90987 224459
rect 91357 216957 92847 224459
rect 93217 216957 94707 224459
rect 95077 216957 98427 224459
rect 10657 149459 98427 216957
rect 10657 144457 18987 149459
rect 19357 144457 20847 149459
rect 21217 144457 36987 149459
rect 37357 144457 38847 149459
rect 39217 144457 54987 149459
rect 55357 144457 56847 149459
rect 57217 144457 72987 149459
rect 73357 144457 74847 149459
rect 75217 144457 90987 149459
rect 91357 144457 92847 149459
rect 93217 144457 98427 149459
rect 10657 76959 98427 144457
rect 10657 345 12147 76959
rect 12517 345 14007 76959
rect 14377 26145 18987 76959
rect 19357 26145 20847 76959
rect 21217 26145 22707 76959
rect 23077 26145 24567 76959
rect 24937 26145 26427 76959
rect 26797 26145 28287 76959
rect 28657 26145 30147 76959
rect 30517 26145 32007 76959
rect 32377 26145 36987 76959
rect 37357 26145 38847 76959
rect 39217 26145 40707 76959
rect 41077 26145 42567 76959
rect 42937 26145 44427 76959
rect 44797 26145 46287 76959
rect 46657 52721 48147 76959
rect 48517 52721 50007 76959
rect 46657 50239 50007 52721
rect 46657 26145 48147 50239
rect 48517 26145 50007 50239
rect 50377 26145 54987 76959
rect 55357 26145 56847 76959
rect 57217 26145 58707 76959
rect 59077 26145 60567 76959
rect 60937 26145 62427 76959
rect 62797 26145 64287 76959
rect 64657 26145 66147 76959
rect 66517 26145 68007 76959
rect 68377 26145 72987 76959
rect 73357 26145 74847 76959
rect 14377 6247 74847 26145
rect 14377 345 18987 6247
rect 19357 345 20847 6247
rect 21217 345 22707 6247
rect 23077 345 36987 6247
rect 37357 345 38847 6247
rect 39217 345 40707 6247
rect 41077 345 54987 6247
rect 55357 345 56847 6247
rect 57217 345 58707 6247
rect 59077 345 72987 6247
rect 73357 345 74847 6247
rect 75217 345 76707 76959
rect 77077 345 78567 76959
rect 78937 345 80427 76959
rect 80797 345 82287 76959
rect 82657 345 84147 76959
rect 84517 345 86007 76959
rect 86377 345 90987 76959
rect 91357 345 92847 76959
rect 93217 345 94707 76959
rect 95077 345 96567 76959
rect 96937 345 98427 76959
rect 98797 345 100287 297855
rect 100657 345 102147 297855
rect 102517 345 104007 297855
rect 104377 291957 110847 297855
rect 111217 291957 112707 297855
rect 113077 291957 114567 297855
rect 114937 291957 116427 297855
rect 116797 291957 128847 297855
rect 129217 291957 130707 297855
rect 131077 291957 132567 297855
rect 132937 291957 134427 297855
rect 134797 291957 146847 297855
rect 147217 291957 148707 297855
rect 149077 291957 150567 297855
rect 150937 291957 152427 297855
rect 152797 291957 164847 297855
rect 165217 291957 166707 297855
rect 167077 291957 168567 297855
rect 168937 291957 170427 297855
rect 170797 291957 182847 297855
rect 183217 291957 184707 297855
rect 185077 291957 186567 297855
rect 186937 291957 188427 297855
rect 188797 291957 194007 297855
rect 104377 224459 194007 291957
rect 104377 216957 108987 224459
rect 109357 216957 110847 224459
rect 111217 216957 112707 224459
rect 113077 216957 126987 224459
rect 127357 216957 128847 224459
rect 129217 216957 130707 224459
rect 131077 216957 144987 224459
rect 145357 216957 146847 224459
rect 147217 216957 148707 224459
rect 149077 216957 162987 224459
rect 163357 216957 164847 224459
rect 165217 216957 166707 224459
rect 167077 216957 180987 224459
rect 181357 216957 182847 224459
rect 183217 216957 184707 224459
rect 185077 216957 194007 224459
rect 104377 149459 194007 216957
rect 104377 144457 108987 149459
rect 109357 144457 110847 149459
rect 111217 144457 126987 149459
rect 127357 144457 128847 149459
rect 129217 144457 144987 149459
rect 145357 144457 146847 149459
rect 147217 144457 162987 149459
rect 163357 144457 164847 149459
rect 165217 144457 180987 149459
rect 181357 144457 182847 149459
rect 183217 144457 194007 149459
rect 104377 76959 194007 144457
rect 104377 345 108987 76959
rect 109357 345 110847 76959
rect 111217 345 112707 76959
rect 113077 345 114567 76959
rect 114937 345 116427 76959
rect 116797 345 118287 76959
rect 118657 345 120147 76959
rect 120517 71957 126987 76959
rect 127357 71957 128847 76959
rect 129217 71957 144987 76959
rect 145357 71957 146847 76959
rect 147217 71957 162987 76959
rect 163357 71957 164847 76959
rect 165217 71957 180987 76959
rect 181357 71957 182847 76959
rect 183217 71957 194007 76959
rect 194377 71957 198987 297855
rect 199357 71957 200847 297855
rect 201217 71957 202707 297855
rect 203077 71957 204567 297855
rect 204937 71957 206427 297855
rect 206797 291957 218847 297855
rect 219217 291957 220707 297855
rect 221077 291957 222567 297855
rect 222937 291957 224427 297855
rect 224797 291957 236847 297855
rect 237217 291957 238707 297855
rect 239077 291957 240567 297855
rect 240937 291957 242427 297855
rect 242797 291957 254847 297855
rect 255217 291957 256707 297855
rect 257077 291957 258567 297855
rect 258937 291957 260427 297855
rect 260797 291957 272847 297855
rect 273217 291957 274707 297855
rect 275077 291957 276567 297855
rect 276937 291957 278427 297855
rect 278797 291957 290847 297855
rect 291217 291957 292707 297855
rect 206797 224459 292707 291957
rect 206797 216957 216987 224459
rect 217357 216957 218847 224459
rect 219217 216957 220707 224459
rect 221077 216957 234987 224459
rect 235357 216957 236847 224459
rect 237217 216957 238707 224459
rect 239077 216957 252987 224459
rect 253357 216957 254847 224459
rect 255217 216957 256707 224459
rect 257077 216957 270987 224459
rect 271357 216957 272847 224459
rect 273217 216957 274707 224459
rect 275077 216957 288987 224459
rect 289357 216957 290847 224459
rect 291217 216957 292707 224459
rect 206797 149459 292707 216957
rect 206797 144457 216987 149459
rect 217357 144457 218847 149459
rect 219217 144457 234987 149459
rect 235357 144457 236847 149459
rect 237217 144457 252987 149459
rect 253357 144457 254847 149459
rect 255217 144457 270987 149459
rect 271357 144457 272847 149459
rect 273217 144457 288987 149459
rect 289357 144457 290847 149459
rect 291217 144457 292707 149459
rect 206797 76959 292707 144457
rect 206797 71957 208287 76959
rect 120517 4459 208287 71957
rect 120517 345 126987 4459
rect 127357 345 128847 4459
rect 129217 345 144987 4459
rect 145357 345 146847 4459
rect 147217 345 162987 4459
rect 163357 345 164847 4459
rect 165217 345 180987 4459
rect 181357 345 182847 4459
rect 183217 345 198987 4459
rect 199357 345 200847 4459
rect 201217 345 208287 4459
rect 208657 345 210147 76959
rect 210517 345 212007 76959
rect 212377 345 216987 76959
rect 217357 345 218847 76959
rect 219217 345 220707 76959
rect 221077 345 222567 76959
rect 222937 345 224427 76959
rect 224797 345 226287 76959
rect 226657 345 228147 76959
rect 228517 345 230007 76959
rect 230377 345 234987 76959
rect 235357 345 236847 76959
rect 237217 345 238707 76959
rect 239077 345 240567 76959
rect 240937 345 242427 76959
rect 242797 345 244287 76959
rect 244657 345 246147 76959
rect 246517 345 248007 76959
rect 248377 345 252987 76959
rect 253357 345 254847 76959
rect 255217 345 256707 76959
rect 257077 345 258567 76959
rect 258937 345 260427 76959
rect 260797 345 262287 76959
rect 262657 345 264147 76959
rect 264517 345 266007 76959
rect 266377 345 270987 76959
rect 271357 345 272847 76959
rect 273217 345 274707 76959
rect 275077 345 276567 76959
rect 276937 345 278427 76959
rect 278797 345 280287 76959
rect 280657 345 282147 76959
rect 282517 345 284007 76959
rect 284377 345 288987 76959
rect 289357 345 290847 76959
rect 291217 345 292707 76959
rect 293077 345 294567 297855
rect 294937 345 295330 297855
<< metal5 >>
rect -4243 302917 304235 303227
rect -3763 302437 303755 302747
rect -3283 301957 303275 302267
rect -2803 301477 302795 301787
rect -2323 300997 302315 301307
rect -1843 300517 301835 300827
rect -1363 300037 301355 300347
rect -883 299557 300875 299867
rect -4243 297353 304235 297663
rect -4243 295493 304235 295803
rect -4243 293633 304235 293943
rect -4243 291773 304235 292083
rect -4243 289913 304235 290223
rect -4243 284933 304235 285243
rect -4243 283073 304235 283383
rect -4243 281213 304235 281523
rect -4243 279353 304235 279663
rect -4243 277493 304235 277803
rect -4243 275633 304235 275943
rect -4243 273773 304235 274083
rect -4243 271913 304235 272223
rect -4243 266933 304235 267243
rect -4243 265073 304235 265383
rect -4243 263213 304235 263523
rect -4243 261353 304235 261663
rect -4243 259493 304235 259803
rect -4243 257633 304235 257943
rect -4243 255773 304235 256083
rect -4243 253913 304235 254223
rect -4243 248933 304235 249243
rect -4243 247073 304235 247383
rect -4243 245213 304235 245523
rect -4243 243353 304235 243663
rect -4243 241493 304235 241803
rect -4243 239633 304235 239943
rect -4243 237773 304235 238083
rect -4243 235913 304235 236223
rect -4243 230933 304235 231243
rect -4243 229073 304235 229383
rect -4243 227213 304235 227523
rect -4243 225353 304235 225663
rect -4243 223493 304235 223803
rect -4243 221633 304235 221943
rect -4243 219773 304235 220083
rect -4243 217913 304235 218223
rect -4243 212933 304235 213243
rect -4243 211073 304235 211383
rect -4243 209213 304235 209523
rect -4243 207353 304235 207663
rect -4243 205493 304235 205803
rect -4243 203633 304235 203943
rect -4243 201773 304235 202083
rect -4243 199913 304235 200223
rect -4243 194933 304235 195243
rect -4243 193073 304235 193383
rect -4243 191213 304235 191523
rect -4243 189353 304235 189663
rect -4243 187493 304235 187803
rect -4243 185633 304235 185943
rect -4243 183773 304235 184083
rect -4243 181913 304235 182223
rect -4243 176933 304235 177243
rect -4243 175073 304235 175383
rect -4243 173213 304235 173523
rect -4243 171353 304235 171663
rect -4243 169493 304235 169803
rect -4243 167633 304235 167943
rect -4243 165773 304235 166083
rect -4243 163913 304235 164223
rect -4243 158933 304235 159243
rect -4243 157073 304235 157383
rect -4243 155213 304235 155523
rect -4243 153353 304235 153663
rect -4243 151493 304235 151803
rect -4243 149633 304235 149943
rect -4243 147773 304235 148083
rect -4243 145913 304235 146223
rect -4243 140933 304235 141243
rect -4243 139073 304235 139383
rect -4243 137213 304235 137523
rect -4243 135353 304235 135663
rect -4243 133493 304235 133803
rect -4243 131633 304235 131943
rect -4243 129773 304235 130083
rect -4243 127913 304235 128223
rect -4243 122933 304235 123243
rect -4243 121073 304235 121383
rect -4243 119213 304235 119523
rect -4243 117353 304235 117663
rect -4243 115493 304235 115803
rect -4243 113633 304235 113943
rect -4243 111773 304235 112083
rect -4243 109913 304235 110223
rect -4243 104933 304235 105243
rect -4243 103073 304235 103383
rect -4243 101213 304235 101523
rect -4243 99353 304235 99663
rect -4243 97493 304235 97803
rect -4243 95633 304235 95943
rect -4243 93773 304235 94083
rect -4243 91913 304235 92223
rect -4243 86933 304235 87243
rect -4243 85073 304235 85383
rect -4243 83213 304235 83523
rect -4243 81353 304235 81663
rect -4243 79493 304235 79803
rect -4243 77633 304235 77943
rect -4243 75773 304235 76083
rect -4243 73913 304235 74223
rect -4243 68933 304235 69243
rect -4243 67073 304235 67383
rect -4243 65213 304235 65523
rect -4243 63353 304235 63663
rect -4243 61493 304235 61803
rect -4243 59633 304235 59943
rect -4243 57773 304235 58083
rect -4243 55913 304235 56223
rect -4243 50933 304235 51243
rect -4243 49073 304235 49383
rect -4243 47213 304235 47523
rect -4243 45353 304235 45663
rect -4243 43493 304235 43803
rect -4243 41633 304235 41943
rect -4243 39773 304235 40083
rect -4243 37913 304235 38223
rect -4243 32933 304235 33243
rect -4243 31073 304235 31383
rect -4243 29213 304235 29523
rect -4243 27353 304235 27663
rect -4243 25493 304235 25803
rect -4243 23633 304235 23943
rect -4243 21773 304235 22083
rect -4243 19913 304235 20223
rect -4243 14933 304235 15243
rect -4243 13073 304235 13383
rect -4243 11213 304235 11523
rect -4243 9353 304235 9663
rect -4243 7493 304235 7803
rect -4243 5633 304235 5943
rect -4243 3773 304235 4083
rect -4243 1913 304235 2223
rect -883 13 300875 323
rect -1363 -467 301355 -157
rect -1843 -947 301835 -637
rect -2323 -1427 302315 -1117
rect -2803 -1907 302795 -1597
rect -3283 -2387 303275 -2077
rect -3763 -2867 303755 -2557
rect -4243 -3347 304235 -3037
<< labels >>
rlabel metal3 s 299760 121660 300480 121772 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 228676 299760 228788 300480 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 195524 299760 195636 300480 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 162372 299760 162484 300480 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 129220 299760 129332 300480 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 96068 299760 96180 300480 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 62916 299760 63028 300480 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 29764 299760 29876 300480 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s -480 296828 240 296940 4 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s -480 274652 240 274764 4 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s -480 252476 240 252588 4 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 299760 144284 300480 144396 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s -480 230300 240 230412 4 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s -480 208124 240 208236 4 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s -480 185948 240 186060 4 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s -480 163772 240 163884 4 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s -480 141596 240 141708 4 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s -480 119420 240 119532 4 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s -480 97244 240 97356 4 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s -480 75068 240 75180 4 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s -480 52892 240 53004 4 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 299760 166908 300480 167020 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 299760 189532 300480 189644 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 299760 212156 300480 212268 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 299760 234780 300480 234892 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 299760 257404 300480 257516 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 299760 280028 300480 280140 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 294980 299760 295092 300480 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 261828 299760 261940 300480 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 299760 2884 300480 2996 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 299760 195188 300480 195300 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 299760 217812 300480 217924 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 299760 240436 300480 240548 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 299760 263060 300480 263172 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 299760 285684 300480 285796 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 286692 299760 286804 300480 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 253540 299760 253652 300480 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 220388 299760 220500 300480 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 187236 299760 187348 300480 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 154084 299760 154196 300480 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 299760 19852 300480 19964 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 120932 299760 121044 300480 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 87780 299760 87892 300480 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 54628 299760 54740 300480 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 21476 299760 21588 300480 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s -480 291284 240 291396 4 io_in[24]
port 46 nsew signal input
rlabel metal3 s -480 269108 240 269220 4 io_in[25]
port 47 nsew signal input
rlabel metal3 s -480 246932 240 247044 4 io_in[26]
port 48 nsew signal input
rlabel metal3 s -480 224756 240 224868 4 io_in[27]
port 49 nsew signal input
rlabel metal3 s -480 202580 240 202692 4 io_in[28]
port 50 nsew signal input
rlabel metal3 s -480 180404 240 180516 4 io_in[29]
port 51 nsew signal input
rlabel metal3 s 299760 36820 300480 36932 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s -480 158228 240 158340 4 io_in[30]
port 53 nsew signal input
rlabel metal3 s -480 136052 240 136164 4 io_in[31]
port 54 nsew signal input
rlabel metal3 s -480 113876 240 113988 4 io_in[32]
port 55 nsew signal input
rlabel metal3 s -480 91700 240 91812 4 io_in[33]
port 56 nsew signal input
rlabel metal3 s -480 69524 240 69636 4 io_in[34]
port 57 nsew signal input
rlabel metal3 s -480 47348 240 47460 4 io_in[35]
port 58 nsew signal input
rlabel metal3 s -480 30716 240 30828 4 io_in[36]
port 59 nsew signal input
rlabel metal3 s -480 14084 240 14196 4 io_in[37]
port 60 nsew signal input
rlabel metal3 s 299760 53788 300480 53900 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 299760 70756 300480 70868 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 299760 87724 300480 87836 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 299760 104692 300480 104804 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 299760 127316 300480 127428 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 299760 149940 300480 150052 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 299760 172564 300480 172676 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 299760 14196 300480 14308 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 299760 206500 300480 206612 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 299760 229124 300480 229236 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 299760 251748 300480 251860 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 299760 274372 300480 274484 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 299760 296996 300480 297108 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 270116 299760 270228 300480 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 236964 299760 237076 300480 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 203812 299760 203924 300480 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 170660 299760 170772 300480 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 137508 299760 137620 300480 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 299760 31164 300480 31276 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 104356 299760 104468 300480 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 71204 299760 71316 300480 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 38052 299760 38164 300480 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 4900 299760 5012 300480 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s -480 280196 240 280308 4 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s -480 258020 240 258132 4 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s -480 235844 240 235956 4 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s -480 213668 240 213780 4 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s -480 191492 240 191604 4 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s -480 169316 240 169428 4 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 299760 48132 300480 48244 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s -480 147140 240 147252 4 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s -480 124964 240 125076 4 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s -480 102788 240 102900 4 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s -480 80612 240 80724 4 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s -480 58436 240 58548 4 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s -480 36260 240 36372 4 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s -480 19628 240 19740 4 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s -480 2996 240 3108 4 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 299760 65100 300480 65212 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 299760 82068 300480 82180 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 299760 99036 300480 99148 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 299760 116004 300480 116116 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 299760 138628 300480 138740 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 299760 161252 300480 161364 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 299760 183876 300480 183988 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 299760 8540 300480 8652 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 299760 200844 300480 200956 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 299760 223468 300480 223580 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 299760 246092 300480 246204 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 299760 268716 300480 268828 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 299760 291340 300480 291452 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 278404 299760 278516 300480 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 245252 299760 245364 300480 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 212100 299760 212212 300480 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 178948 299760 179060 300480 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 145796 299760 145908 300480 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 299760 25508 300480 25620 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 112644 299760 112756 300480 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 79492 299760 79604 300480 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 46340 299760 46452 300480 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 13188 299760 13300 300480 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s -480 285740 240 285852 4 io_out[24]
port 122 nsew signal output
rlabel metal3 s -480 263564 240 263676 4 io_out[25]
port 123 nsew signal output
rlabel metal3 s -480 241388 240 241500 4 io_out[26]
port 124 nsew signal output
rlabel metal3 s -480 219212 240 219324 4 io_out[27]
port 125 nsew signal output
rlabel metal3 s -480 197036 240 197148 4 io_out[28]
port 126 nsew signal output
rlabel metal3 s -480 174860 240 174972 4 io_out[29]
port 127 nsew signal output
rlabel metal3 s 299760 42476 300480 42588 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s -480 152684 240 152796 4 io_out[30]
port 129 nsew signal output
rlabel metal3 s -480 130508 240 130620 4 io_out[31]
port 130 nsew signal output
rlabel metal3 s -480 108332 240 108444 4 io_out[32]
port 131 nsew signal output
rlabel metal3 s -480 86156 240 86268 4 io_out[33]
port 132 nsew signal output
rlabel metal3 s -480 63980 240 64092 4 io_out[34]
port 133 nsew signal output
rlabel metal3 s -480 41804 240 41916 4 io_out[35]
port 134 nsew signal output
rlabel metal3 s -480 25172 240 25284 4 io_out[36]
port 135 nsew signal output
rlabel metal3 s -480 8540 240 8652 4 io_out[37]
port 136 nsew signal output
rlabel metal3 s 299760 59444 300480 59556 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 299760 76412 300480 76524 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 299760 93380 300480 93492 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 299760 110348 300480 110460 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 299760 132972 300480 133084 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 299760 155596 300480 155708 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 299760 178220 300480 178332 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 71260 -480 71372 240 8 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 239260 -480 239372 240 8 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 240940 -480 241052 240 8 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 242620 -480 242732 240 8 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 244300 -480 244412 240 8 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 245980 -480 246092 240 8 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 247660 -480 247772 240 8 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 249340 -480 249452 240 8 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 251020 -480 251132 240 8 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 252700 -480 252812 240 8 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 254380 -480 254492 240 8 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 88060 -480 88172 240 8 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 256060 -480 256172 240 8 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 257740 -480 257852 240 8 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 259420 -480 259532 240 8 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 261100 -480 261212 240 8 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 262780 -480 262892 240 8 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 264460 -480 264572 240 8 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 266140 -480 266252 240 8 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 267820 -480 267932 240 8 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 269500 -480 269612 240 8 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 271180 -480 271292 240 8 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 89740 -480 89852 240 8 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 272860 -480 272972 240 8 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 274540 -480 274652 240 8 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 276220 -480 276332 240 8 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 277900 -480 278012 240 8 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 279580 -480 279692 240 8 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 281260 -480 281372 240 8 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 282940 -480 283052 240 8 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 284620 -480 284732 240 8 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 91420 -480 91532 240 8 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 93100 -480 93212 240 8 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 94780 -480 94892 240 8 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 96460 -480 96572 240 8 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 98140 -480 98252 240 8 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 99820 -480 99932 240 8 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 101500 -480 101612 240 8 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 103180 -480 103292 240 8 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 72940 -480 73052 240 8 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 104860 -480 104972 240 8 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 106540 -480 106652 240 8 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 108220 -480 108332 240 8 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 109900 -480 110012 240 8 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 111580 -480 111692 240 8 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 113260 -480 113372 240 8 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 114940 -480 115052 240 8 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 116620 -480 116732 240 8 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 118300 -480 118412 240 8 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 119980 -480 120092 240 8 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 74620 -480 74732 240 8 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 121660 -480 121772 240 8 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 123340 -480 123452 240 8 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 125020 -480 125132 240 8 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 126700 -480 126812 240 8 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 128380 -480 128492 240 8 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 130060 -480 130172 240 8 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 131740 -480 131852 240 8 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 133420 -480 133532 240 8 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 135100 -480 135212 240 8 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 136780 -480 136892 240 8 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 76300 -480 76412 240 8 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 138460 -480 138572 240 8 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 140140 -480 140252 240 8 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 141820 -480 141932 240 8 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 143500 -480 143612 240 8 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 145180 -480 145292 240 8 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 146860 -480 146972 240 8 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 148540 -480 148652 240 8 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 150220 -480 150332 240 8 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 151900 -480 152012 240 8 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 153580 -480 153692 240 8 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 77980 -480 78092 240 8 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 155260 -480 155372 240 8 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 156940 -480 157052 240 8 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 158620 -480 158732 240 8 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 160300 -480 160412 240 8 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 161980 -480 162092 240 8 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 163660 -480 163772 240 8 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 165340 -480 165452 240 8 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 167020 -480 167132 240 8 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 168700 -480 168812 240 8 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 170380 -480 170492 240 8 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 79660 -480 79772 240 8 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 172060 -480 172172 240 8 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 173740 -480 173852 240 8 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 175420 -480 175532 240 8 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 177100 -480 177212 240 8 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 178780 -480 178892 240 8 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 180460 -480 180572 240 8 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 182140 -480 182252 240 8 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 183820 -480 183932 240 8 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 185500 -480 185612 240 8 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 187180 -480 187292 240 8 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 81340 -480 81452 240 8 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 188860 -480 188972 240 8 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 190540 -480 190652 240 8 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 192220 -480 192332 240 8 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 193900 -480 194012 240 8 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 195580 -480 195692 240 8 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 197260 -480 197372 240 8 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 198940 -480 199052 240 8 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 200620 -480 200732 240 8 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 202300 -480 202412 240 8 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 203980 -480 204092 240 8 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 83020 -480 83132 240 8 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 205660 -480 205772 240 8 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 207340 -480 207452 240 8 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 209020 -480 209132 240 8 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 210700 -480 210812 240 8 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 212380 -480 212492 240 8 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 214060 -480 214172 240 8 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 215740 -480 215852 240 8 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 217420 -480 217532 240 8 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 219100 -480 219212 240 8 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 220780 -480 220892 240 8 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 84700 -480 84812 240 8 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 222460 -480 222572 240 8 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 224140 -480 224252 240 8 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 225820 -480 225932 240 8 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 227500 -480 227612 240 8 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 229180 -480 229292 240 8 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 230860 -480 230972 240 8 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 232540 -480 232652 240 8 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 234220 -480 234332 240 8 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 235900 -480 236012 240 8 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 237580 -480 237692 240 8 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 86380 -480 86492 240 8 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 71820 -480 71932 240 8 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 239820 -480 239932 240 8 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 241500 -480 241612 240 8 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 243180 -480 243292 240 8 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 244860 -480 244972 240 8 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 246540 -480 246652 240 8 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 248220 -480 248332 240 8 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 249900 -480 250012 240 8 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 251580 -480 251692 240 8 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 253260 -480 253372 240 8 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 254940 -480 255052 240 8 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 88620 -480 88732 240 8 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 256620 -480 256732 240 8 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 258300 -480 258412 240 8 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 259980 -480 260092 240 8 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 261660 -480 261772 240 8 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 263340 -480 263452 240 8 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 265020 -480 265132 240 8 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 266700 -480 266812 240 8 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 268380 -480 268492 240 8 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 270060 -480 270172 240 8 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 271740 -480 271852 240 8 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 90300 -480 90412 240 8 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 273420 -480 273532 240 8 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 275100 -480 275212 240 8 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 276780 -480 276892 240 8 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 278460 -480 278572 240 8 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 280140 -480 280252 240 8 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 281820 -480 281932 240 8 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 283500 -480 283612 240 8 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 285180 -480 285292 240 8 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 91980 -480 92092 240 8 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 93660 -480 93772 240 8 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 95340 -480 95452 240 8 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 97020 -480 97132 240 8 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 98700 -480 98812 240 8 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 100380 -480 100492 240 8 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 102060 -480 102172 240 8 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 103740 -480 103852 240 8 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 73500 -480 73612 240 8 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 105420 -480 105532 240 8 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 107100 -480 107212 240 8 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 108780 -480 108892 240 8 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 110460 -480 110572 240 8 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 112140 -480 112252 240 8 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 113820 -480 113932 240 8 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 115500 -480 115612 240 8 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 117180 -480 117292 240 8 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 118860 -480 118972 240 8 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 120540 -480 120652 240 8 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 75180 -480 75292 240 8 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 122220 -480 122332 240 8 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 123900 -480 124012 240 8 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 125580 -480 125692 240 8 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 127260 -480 127372 240 8 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 128940 -480 129052 240 8 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 130620 -480 130732 240 8 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 132300 -480 132412 240 8 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 133980 -480 134092 240 8 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 135660 -480 135772 240 8 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 137340 -480 137452 240 8 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 76860 -480 76972 240 8 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 139020 -480 139132 240 8 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 140700 -480 140812 240 8 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 142380 -480 142492 240 8 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 144060 -480 144172 240 8 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 145740 -480 145852 240 8 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 147420 -480 147532 240 8 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 149100 -480 149212 240 8 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 150780 -480 150892 240 8 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 152460 -480 152572 240 8 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 154140 -480 154252 240 8 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 78540 -480 78652 240 8 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 155820 -480 155932 240 8 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 157500 -480 157612 240 8 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 159180 -480 159292 240 8 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 160860 -480 160972 240 8 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 162540 -480 162652 240 8 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 164220 -480 164332 240 8 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 165900 -480 166012 240 8 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 167580 -480 167692 240 8 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 169260 -480 169372 240 8 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 170940 -480 171052 240 8 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 80220 -480 80332 240 8 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 172620 -480 172732 240 8 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 174300 -480 174412 240 8 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 175980 -480 176092 240 8 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 177660 -480 177772 240 8 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 179340 -480 179452 240 8 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 181020 -480 181132 240 8 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 182700 -480 182812 240 8 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 184380 -480 184492 240 8 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 186060 -480 186172 240 8 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 187740 -480 187852 240 8 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 81900 -480 82012 240 8 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 189420 -480 189532 240 8 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 191100 -480 191212 240 8 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 192780 -480 192892 240 8 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 194460 -480 194572 240 8 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 196140 -480 196252 240 8 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 197820 -480 197932 240 8 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 199500 -480 199612 240 8 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 201180 -480 201292 240 8 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 202860 -480 202972 240 8 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 204540 -480 204652 240 8 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 83580 -480 83692 240 8 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 206220 -480 206332 240 8 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 207900 -480 208012 240 8 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 209580 -480 209692 240 8 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 211260 -480 211372 240 8 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 212940 -480 213052 240 8 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 214620 -480 214732 240 8 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 216300 -480 216412 240 8 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 217980 -480 218092 240 8 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 219660 -480 219772 240 8 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 221340 -480 221452 240 8 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 85260 -480 85372 240 8 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 223020 -480 223132 240 8 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 224700 -480 224812 240 8 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 226380 -480 226492 240 8 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 228060 -480 228172 240 8 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 229740 -480 229852 240 8 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 231420 -480 231532 240 8 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 233100 -480 233212 240 8 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 234780 -480 234892 240 8 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 236460 -480 236572 240 8 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 238140 -480 238252 240 8 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 86940 -480 87052 240 8 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 72380 -480 72492 240 8 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 240380 -480 240492 240 8 la_oenb[100]
port 401 nsew signal input
rlabel metal2 s 242060 -480 242172 240 8 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 243740 -480 243852 240 8 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 245420 -480 245532 240 8 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 247100 -480 247212 240 8 la_oenb[104]
port 405 nsew signal input
rlabel metal2 s 248780 -480 248892 240 8 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 250460 -480 250572 240 8 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 252140 -480 252252 240 8 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 253820 -480 253932 240 8 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 255500 -480 255612 240 8 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 89180 -480 89292 240 8 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 257180 -480 257292 240 8 la_oenb[110]
port 412 nsew signal input
rlabel metal2 s 258860 -480 258972 240 8 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 260540 -480 260652 240 8 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 262220 -480 262332 240 8 la_oenb[113]
port 415 nsew signal input
rlabel metal2 s 263900 -480 264012 240 8 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 265580 -480 265692 240 8 la_oenb[115]
port 417 nsew signal input
rlabel metal2 s 267260 -480 267372 240 8 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 268940 -480 269052 240 8 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 270620 -480 270732 240 8 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 272300 -480 272412 240 8 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 90860 -480 90972 240 8 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 273980 -480 274092 240 8 la_oenb[120]
port 423 nsew signal input
rlabel metal2 s 275660 -480 275772 240 8 la_oenb[121]
port 424 nsew signal input
rlabel metal2 s 277340 -480 277452 240 8 la_oenb[122]
port 425 nsew signal input
rlabel metal2 s 279020 -480 279132 240 8 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 280700 -480 280812 240 8 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 282380 -480 282492 240 8 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 284060 -480 284172 240 8 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 285740 -480 285852 240 8 la_oenb[127]
port 430 nsew signal input
rlabel metal2 s 92540 -480 92652 240 8 la_oenb[12]
port 431 nsew signal input
rlabel metal2 s 94220 -480 94332 240 8 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 95900 -480 96012 240 8 la_oenb[14]
port 433 nsew signal input
rlabel metal2 s 97580 -480 97692 240 8 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 99260 -480 99372 240 8 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 100940 -480 101052 240 8 la_oenb[17]
port 436 nsew signal input
rlabel metal2 s 102620 -480 102732 240 8 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 104300 -480 104412 240 8 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 74060 -480 74172 240 8 la_oenb[1]
port 439 nsew signal input
rlabel metal2 s 105980 -480 106092 240 8 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 107660 -480 107772 240 8 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 109340 -480 109452 240 8 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 111020 -480 111132 240 8 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 112700 -480 112812 240 8 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 114380 -480 114492 240 8 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 116060 -480 116172 240 8 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 117740 -480 117852 240 8 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 119420 -480 119532 240 8 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 121100 -480 121212 240 8 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 75740 -480 75852 240 8 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 122780 -480 122892 240 8 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 124460 -480 124572 240 8 la_oenb[31]
port 452 nsew signal input
rlabel metal2 s 126140 -480 126252 240 8 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 127820 -480 127932 240 8 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 129500 -480 129612 240 8 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 131180 -480 131292 240 8 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 132860 -480 132972 240 8 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 134540 -480 134652 240 8 la_oenb[37]
port 458 nsew signal input
rlabel metal2 s 136220 -480 136332 240 8 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 137900 -480 138012 240 8 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 77420 -480 77532 240 8 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 139580 -480 139692 240 8 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 141260 -480 141372 240 8 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 142940 -480 143052 240 8 la_oenb[42]
port 464 nsew signal input
rlabel metal2 s 144620 -480 144732 240 8 la_oenb[43]
port 465 nsew signal input
rlabel metal2 s 146300 -480 146412 240 8 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 147980 -480 148092 240 8 la_oenb[45]
port 467 nsew signal input
rlabel metal2 s 149660 -480 149772 240 8 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 151340 -480 151452 240 8 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 153020 -480 153132 240 8 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 154700 -480 154812 240 8 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 79100 -480 79212 240 8 la_oenb[4]
port 472 nsew signal input
rlabel metal2 s 156380 -480 156492 240 8 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 158060 -480 158172 240 8 la_oenb[51]
port 474 nsew signal input
rlabel metal2 s 159740 -480 159852 240 8 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 161420 -480 161532 240 8 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 163100 -480 163212 240 8 la_oenb[54]
port 477 nsew signal input
rlabel metal2 s 164780 -480 164892 240 8 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 166460 -480 166572 240 8 la_oenb[56]
port 479 nsew signal input
rlabel metal2 s 168140 -480 168252 240 8 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 169820 -480 169932 240 8 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 171500 -480 171612 240 8 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 80780 -480 80892 240 8 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 173180 -480 173292 240 8 la_oenb[60]
port 484 nsew signal input
rlabel metal2 s 174860 -480 174972 240 8 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 176540 -480 176652 240 8 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 178220 -480 178332 240 8 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 179900 -480 180012 240 8 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 181580 -480 181692 240 8 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 183260 -480 183372 240 8 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 184940 -480 185052 240 8 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 186620 -480 186732 240 8 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 188300 -480 188412 240 8 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 82460 -480 82572 240 8 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 189980 -480 190092 240 8 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 191660 -480 191772 240 8 la_oenb[71]
port 496 nsew signal input
rlabel metal2 s 193340 -480 193452 240 8 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 195020 -480 195132 240 8 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 196700 -480 196812 240 8 la_oenb[74]
port 499 nsew signal input
rlabel metal2 s 198380 -480 198492 240 8 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 200060 -480 200172 240 8 la_oenb[76]
port 501 nsew signal input
rlabel metal2 s 201740 -480 201852 240 8 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 203420 -480 203532 240 8 la_oenb[78]
port 503 nsew signal input
rlabel metal2 s 205100 -480 205212 240 8 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 84140 -480 84252 240 8 la_oenb[7]
port 505 nsew signal input
rlabel metal2 s 206780 -480 206892 240 8 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 208460 -480 208572 240 8 la_oenb[81]
port 507 nsew signal input
rlabel metal2 s 210140 -480 210252 240 8 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 211820 -480 211932 240 8 la_oenb[83]
port 509 nsew signal input
rlabel metal2 s 213500 -480 213612 240 8 la_oenb[84]
port 510 nsew signal input
rlabel metal2 s 215180 -480 215292 240 8 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 216860 -480 216972 240 8 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 218540 -480 218652 240 8 la_oenb[87]
port 513 nsew signal input
rlabel metal2 s 220220 -480 220332 240 8 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 221900 -480 222012 240 8 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 85820 -480 85932 240 8 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 223580 -480 223692 240 8 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 225260 -480 225372 240 8 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 226940 -480 227052 240 8 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 228620 -480 228732 240 8 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 230300 -480 230412 240 8 la_oenb[94]
port 521 nsew signal input
rlabel metal2 s 231980 -480 232092 240 8 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 233660 -480 233772 240 8 la_oenb[96]
port 523 nsew signal input
rlabel metal2 s 235340 -480 235452 240 8 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 237020 -480 237132 240 8 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 238700 -480 238812 240 8 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 87500 -480 87612 240 8 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 286300 -480 286412 240 8 user_clock2
port 528 nsew signal input
rlabel metal2 s 286860 -480 286972 240 8 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 287420 -480 287532 240 8 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 287980 -480 288092 240 8 user_irq[2]
port 531 nsew signal output
rlabel metal4 s -883 13 -573 299867 4 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -883 13 300875 323 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -883 299557 300875 299867 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 300565 13 300875 299867 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 1017 -3347 1327 303227 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 19017 -3347 19327 6217 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 19017 26175 19327 76929 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 19017 144487 19327 149429 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 19017 216987 19327 224429 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 37017 -3347 37327 6217 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 37017 26175 37327 76929 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 37017 144487 37327 149429 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 37017 216987 37327 224429 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 55017 -3347 55327 6217 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 55017 26175 55327 76929 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 55017 144487 55327 149429 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 55017 216987 55327 224429 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 73017 -3347 73327 6217 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 73017 26175 73327 76929 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 73017 144487 73327 149429 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 73017 216987 73327 224429 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 91017 -3347 91327 76929 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 91017 144487 91327 149429 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 91017 216987 91327 224429 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 109017 -3347 109327 76929 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 109017 144487 109327 149429 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 109017 216987 109327 224429 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 127017 -3347 127327 4429 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 127017 71987 127327 76929 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 127017 144487 127327 149429 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 127017 216987 127327 224429 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 145017 -3347 145327 4429 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 145017 71987 145327 76929 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 145017 144487 145327 149429 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 145017 216987 145327 224429 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 163017 -3347 163327 4429 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 163017 71987 163327 76929 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 163017 144487 163327 149429 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 163017 216987 163327 224429 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 181017 -3347 181327 4429 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 181017 71987 181327 76929 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 181017 144487 181327 149429 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 181017 216987 181327 224429 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 199017 -3347 199327 4429 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 199017 71987 199327 303227 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 217017 -3347 217327 76929 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 217017 144487 217327 149429 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 217017 216987 217327 224429 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 235017 -3347 235327 76929 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 235017 144487 235327 149429 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 235017 216987 235327 224429 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 253017 -3347 253327 76929 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 253017 144487 253327 149429 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 253017 216987 253327 224429 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 271017 -3347 271327 76929 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 271017 144487 271327 149429 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 271017 216987 271327 224429 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 289017 -3347 289327 76929 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 289017 144487 289327 149429 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 289017 216987 289327 224429 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -4243 1913 304235 2223 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -4243 19913 304235 20223 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -4243 37913 304235 38223 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -4243 55913 304235 56223 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -4243 73913 304235 74223 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -4243 91913 304235 92223 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -4243 109913 304235 110223 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -4243 127913 304235 128223 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -4243 145913 304235 146223 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -4243 163913 304235 164223 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -4243 181913 304235 182223 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -4243 199913 304235 200223 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -4243 217913 304235 218223 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -4243 235913 304235 236223 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -4243 253913 304235 254223 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -4243 271913 304235 272223 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -4243 289913 304235 290223 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s -1843 -947 -1533 300827 4 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -1843 -947 301835 -637 8 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -1843 300517 301835 300827 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 301525 -947 301835 300827 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 4737 -3347 5047 303227 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 22737 -3347 23047 6217 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 22737 26175 23047 76929 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 22737 216987 23047 224429 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 22737 291987 23047 303227 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 40737 -3347 41047 6217 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 40737 26175 41047 76929 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 40737 216987 41047 224429 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 40737 291987 41047 303227 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 58737 -3347 59047 6217 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 58737 26175 59047 76929 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 58737 216987 59047 224429 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 58737 291987 59047 303227 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 76737 -3347 77047 76929 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 76737 216987 77047 224429 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 76737 291987 77047 303227 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 94737 -3347 95047 76929 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 94737 216987 95047 224429 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 94737 291987 95047 303227 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 112737 -3347 113047 76929 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 112737 216987 113047 224429 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 112737 291987 113047 303227 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 130737 216987 131047 224429 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 130737 291987 131047 303227 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 148737 216987 149047 224429 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 148737 291987 149047 303227 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 166737 216987 167047 224429 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 166737 291987 167047 303227 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 184737 216987 185047 224429 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 184737 291987 185047 303227 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 202737 71987 203047 303227 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 220737 -3347 221047 76929 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 220737 216987 221047 224429 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 220737 291987 221047 303227 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 238737 -3347 239047 76929 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 238737 216987 239047 224429 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 238737 291987 239047 303227 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 256737 -3347 257047 76929 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 256737 216987 257047 224429 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 256737 291987 257047 303227 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 274737 -3347 275047 76929 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 274737 216987 275047 224429 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 274737 291987 275047 303227 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 292737 -3347 293047 303227 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4243 5633 304235 5943 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4243 23633 304235 23943 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4243 41633 304235 41943 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4243 59633 304235 59943 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4243 77633 304235 77943 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4243 95633 304235 95943 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4243 113633 304235 113943 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4243 131633 304235 131943 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4243 149633 304235 149943 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4243 167633 304235 167943 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4243 185633 304235 185943 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4243 203633 304235 203943 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4243 221633 304235 221943 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4243 239633 304235 239943 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4243 257633 304235 257943 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4243 275633 304235 275943 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4243 293633 304235 293943 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s -2803 -1907 -2493 301787 4 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -2803 -1907 302795 -1597 8 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -2803 301477 302795 301787 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 302485 -1907 302795 301787 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 8457 -3347 8767 303227 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 26457 26175 26767 76929 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 26457 291987 26767 303227 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 44457 26175 44767 76929 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 44457 291987 44767 303227 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 62457 26175 62767 76929 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 62457 291987 62767 303227 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 80457 -3347 80767 76929 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 80457 291987 80767 303227 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 98457 -3347 98767 303227 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 116457 -3347 116767 76929 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 116457 291987 116767 303227 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 134457 291987 134767 303227 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 152457 291987 152767 303227 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 170457 291987 170767 303227 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 188457 291987 188767 303227 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 206457 71987 206767 303227 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 224457 -3347 224767 76929 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 224457 291987 224767 303227 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 242457 -3347 242767 76929 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 242457 291987 242767 303227 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 260457 -3347 260767 76929 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 260457 291987 260767 303227 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 278457 -3347 278767 76929 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 278457 291987 278767 303227 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 296457 -3347 296767 303227 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -4243 9353 304235 9663 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -4243 27353 304235 27663 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -4243 45353 304235 45663 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -4243 63353 304235 63663 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -4243 81353 304235 81663 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -4243 99353 304235 99663 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -4243 117353 304235 117663 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -4243 135353 304235 135663 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -4243 153353 304235 153663 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -4243 171353 304235 171663 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -4243 189353 304235 189663 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -4243 207353 304235 207663 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -4243 225353 304235 225663 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -4243 243353 304235 243663 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -4243 261353 304235 261663 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -4243 279353 304235 279663 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -4243 297353 304235 297663 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s -3763 -2867 -3453 302747 4 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -3763 -2867 303755 -2557 8 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -3763 302437 303755 302747 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 303445 -2867 303755 302747 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 12177 -3347 12487 76929 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 30177 26175 30487 76929 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 48177 26175 48487 50209 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 48177 52751 48487 76929 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 66177 26175 66487 76929 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 84177 -3347 84487 76929 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 102177 -3347 102487 303227 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 120177 -3347 120487 76929 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 210177 -3347 210487 76929 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 228177 -3347 228487 76929 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 246177 -3347 246487 76929 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 264177 -3347 264487 76929 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 282177 -3347 282487 76929 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -4243 13073 304235 13383 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -4243 31073 304235 31383 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -4243 49073 304235 49383 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -4243 67073 304235 67383 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -4243 85073 304235 85383 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -4243 103073 304235 103383 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -4243 121073 304235 121383 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -4243 139073 304235 139383 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -4243 157073 304235 157383 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -4243 175073 304235 175383 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -4243 193073 304235 193383 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -4243 211073 304235 211383 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -4243 229073 304235 229383 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -4243 247073 304235 247383 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -4243 265073 304235 265383 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -4243 283073 304235 283383 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s -3283 -2387 -2973 302267 4 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -3283 -2387 303275 -2077 8 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -3283 301957 303275 302267 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 302965 -2387 303275 302267 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 10317 -3347 10627 303227 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 28317 26175 28627 76929 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 46317 26175 46627 76929 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 64317 26175 64627 76929 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 82317 -3347 82627 76929 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 100317 -3347 100627 303227 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 118317 -3347 118627 76929 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 208317 -3347 208627 76929 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 226317 -3347 226627 76929 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 244317 -3347 244627 76929 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 262317 -3347 262627 76929 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 280317 -3347 280627 76929 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 298317 -3347 298627 303227 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -4243 11213 304235 11523 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -4243 29213 304235 29523 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -4243 47213 304235 47523 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -4243 65213 304235 65523 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -4243 83213 304235 83523 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -4243 101213 304235 101523 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -4243 119213 304235 119523 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -4243 137213 304235 137523 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -4243 155213 304235 155523 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -4243 173213 304235 173523 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -4243 191213 304235 191523 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -4243 209213 304235 209523 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -4243 227213 304235 227523 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -4243 245213 304235 245523 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -4243 263213 304235 263523 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -4243 281213 304235 281523 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s -4243 -3347 -3933 303227 4 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -4243 -3347 304235 -3037 8 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -4243 302917 304235 303227 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 303925 -3347 304235 303227 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 14037 -3347 14347 76929 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 32037 26175 32347 76929 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 50037 26175 50347 76929 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 68037 26175 68347 76929 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 86037 -3347 86347 76929 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 104037 -3347 104347 303227 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 194037 71987 194347 303227 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 212037 -3347 212347 76929 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 230037 -3347 230347 76929 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 248037 -3347 248347 76929 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 266037 -3347 266347 76929 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 284037 -3347 284347 76929 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -4243 14933 304235 15243 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -4243 32933 304235 33243 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -4243 50933 304235 51243 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -4243 68933 304235 69243 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -4243 86933 304235 87243 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -4243 104933 304235 105243 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -4243 122933 304235 123243 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -4243 140933 304235 141243 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -4243 158933 304235 159243 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -4243 176933 304235 177243 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -4243 194933 304235 195243 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -4243 212933 304235 213243 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -4243 230933 304235 231243 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -4243 248933 304235 249243 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -4243 266933 304235 267243 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -4243 284933 304235 285243 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s -1363 -467 -1053 300347 4 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -1363 -467 301355 -157 8 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -1363 300037 301355 300347 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 301045 -467 301355 300347 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 2877 -3347 3187 303227 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 20877 -3347 21187 6217 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 20877 26175 21187 76929 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 20877 144487 21187 149429 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 20877 216987 21187 224429 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 20877 291987 21187 303227 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 38877 -3347 39187 6217 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 38877 26175 39187 76929 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 38877 144487 39187 149429 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 38877 216987 39187 224429 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 38877 291987 39187 303227 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 56877 -3347 57187 6217 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 56877 26175 57187 76929 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 56877 144487 57187 149429 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 56877 216987 57187 224429 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 56877 291987 57187 303227 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 74877 -3347 75187 76929 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 74877 144487 75187 149429 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 74877 216987 75187 224429 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 74877 291987 75187 303227 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 92877 -3347 93187 76929 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 92877 144487 93187 149429 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 92877 216987 93187 224429 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 92877 291987 93187 303227 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 110877 -3347 111187 76929 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 110877 144487 111187 149429 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 110877 216987 111187 224429 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 110877 291987 111187 303227 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 128877 -3347 129187 4429 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 128877 71987 129187 76929 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 128877 144487 129187 149429 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 128877 216987 129187 224429 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 128877 291987 129187 303227 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 146877 -3347 147187 4429 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 146877 71987 147187 76929 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 146877 144487 147187 149429 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 146877 216987 147187 224429 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 146877 291987 147187 303227 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 164877 -3347 165187 4429 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 164877 71987 165187 76929 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 164877 144487 165187 149429 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 164877 216987 165187 224429 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 164877 291987 165187 303227 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 182877 -3347 183187 4429 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 182877 71987 183187 76929 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 182877 144487 183187 149429 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 182877 216987 183187 224429 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 182877 291987 183187 303227 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 200877 -3347 201187 4429 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 200877 71987 201187 303227 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 218877 -3347 219187 76929 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 218877 144487 219187 149429 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 218877 216987 219187 224429 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 218877 291987 219187 303227 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 236877 -3347 237187 76929 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 236877 144487 237187 149429 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 236877 216987 237187 224429 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 236877 291987 237187 303227 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 254877 -3347 255187 76929 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 254877 144487 255187 149429 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 254877 216987 255187 224429 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 254877 291987 255187 303227 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 272877 -3347 273187 76929 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 272877 144487 273187 149429 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 272877 216987 273187 224429 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 272877 291987 273187 303227 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 290877 -3347 291187 76929 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 290877 144487 291187 149429 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 290877 216987 291187 224429 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 290877 291987 291187 303227 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -4243 3773 304235 4083 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -4243 21773 304235 22083 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -4243 39773 304235 40083 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -4243 57773 304235 58083 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -4243 75773 304235 76083 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -4243 93773 304235 94083 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -4243 111773 304235 112083 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -4243 129773 304235 130083 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -4243 147773 304235 148083 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -4243 165773 304235 166083 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -4243 183773 304235 184083 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -4243 201773 304235 202083 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -4243 219773 304235 220083 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -4243 237773 304235 238083 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -4243 255773 304235 256083 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -4243 273773 304235 274083 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -4243 291773 304235 292083 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s -2323 -1427 -2013 301307 4 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -2323 -1427 302315 -1117 8 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -2323 300997 302315 301307 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 302005 -1427 302315 301307 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 6597 -3347 6907 303227 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 24597 26175 24907 76929 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 24597 291987 24907 303227 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 42597 26175 42907 76929 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 42597 291987 42907 303227 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 60597 26175 60907 76929 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 60597 291987 60907 303227 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 78597 -3347 78907 76929 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 78597 291987 78907 303227 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 96597 -3347 96907 76929 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 96597 291987 96907 303227 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 114597 -3347 114907 76929 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 114597 291987 114907 303227 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 132597 291987 132907 303227 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 150597 291987 150907 303227 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 168597 291987 168907 303227 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 186597 291987 186907 303227 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 204597 71987 204907 303227 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 222597 -3347 222907 76929 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 222597 291987 222907 303227 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 240597 -3347 240907 76929 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 240597 291987 240907 303227 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 258597 -3347 258907 76929 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 258597 291987 258907 303227 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 276597 -3347 276907 76929 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 276597 291987 276907 303227 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 294597 -3347 294907 303227 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -4243 7493 304235 7803 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -4243 25493 304235 25803 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -4243 43493 304235 43803 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -4243 61493 304235 61803 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -4243 79493 304235 79803 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -4243 97493 304235 97803 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -4243 115493 304235 115803 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -4243 133493 304235 133803 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -4243 151493 304235 151803 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -4243 169493 304235 169803 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -4243 187493 304235 187803 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -4243 205493 304235 205803 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -4243 223493 304235 223803 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -4243 241493 304235 241803 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -4243 259493 304235 259803 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -4243 277493 304235 277803 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -4243 295493 304235 295803 6 vssd2
port 539 nsew ground bidirectional
rlabel metal2 s 11900 -480 12012 240 8 wb_clk_i
port 540 nsew signal input
rlabel metal2 s 12460 -480 12572 240 8 wb_rst_i
port 541 nsew signal input
rlabel metal2 s 13020 -480 13132 240 8 wbs_ack_o
port 542 nsew signal output
rlabel metal2 s 15260 -480 15372 240 8 wbs_adr_i[0]
port 543 nsew signal input
rlabel metal2 s 34300 -480 34412 240 8 wbs_adr_i[10]
port 544 nsew signal input
rlabel metal2 s 35980 -480 36092 240 8 wbs_adr_i[11]
port 545 nsew signal input
rlabel metal2 s 37660 -480 37772 240 8 wbs_adr_i[12]
port 546 nsew signal input
rlabel metal2 s 39340 -480 39452 240 8 wbs_adr_i[13]
port 547 nsew signal input
rlabel metal2 s 41020 -480 41132 240 8 wbs_adr_i[14]
port 548 nsew signal input
rlabel metal2 s 42700 -480 42812 240 8 wbs_adr_i[15]
port 549 nsew signal input
rlabel metal2 s 44380 -480 44492 240 8 wbs_adr_i[16]
port 550 nsew signal input
rlabel metal2 s 46060 -480 46172 240 8 wbs_adr_i[17]
port 551 nsew signal input
rlabel metal2 s 47740 -480 47852 240 8 wbs_adr_i[18]
port 552 nsew signal input
rlabel metal2 s 49420 -480 49532 240 8 wbs_adr_i[19]
port 553 nsew signal input
rlabel metal2 s 17500 -480 17612 240 8 wbs_adr_i[1]
port 554 nsew signal input
rlabel metal2 s 51100 -480 51212 240 8 wbs_adr_i[20]
port 555 nsew signal input
rlabel metal2 s 52780 -480 52892 240 8 wbs_adr_i[21]
port 556 nsew signal input
rlabel metal2 s 54460 -480 54572 240 8 wbs_adr_i[22]
port 557 nsew signal input
rlabel metal2 s 56140 -480 56252 240 8 wbs_adr_i[23]
port 558 nsew signal input
rlabel metal2 s 57820 -480 57932 240 8 wbs_adr_i[24]
port 559 nsew signal input
rlabel metal2 s 59500 -480 59612 240 8 wbs_adr_i[25]
port 560 nsew signal input
rlabel metal2 s 61180 -480 61292 240 8 wbs_adr_i[26]
port 561 nsew signal input
rlabel metal2 s 62860 -480 62972 240 8 wbs_adr_i[27]
port 562 nsew signal input
rlabel metal2 s 64540 -480 64652 240 8 wbs_adr_i[28]
port 563 nsew signal input
rlabel metal2 s 66220 -480 66332 240 8 wbs_adr_i[29]
port 564 nsew signal input
rlabel metal2 s 19740 -480 19852 240 8 wbs_adr_i[2]
port 565 nsew signal input
rlabel metal2 s 67900 -480 68012 240 8 wbs_adr_i[30]
port 566 nsew signal input
rlabel metal2 s 69580 -480 69692 240 8 wbs_adr_i[31]
port 567 nsew signal input
rlabel metal2 s 21980 -480 22092 240 8 wbs_adr_i[3]
port 568 nsew signal input
rlabel metal2 s 24220 -480 24332 240 8 wbs_adr_i[4]
port 569 nsew signal input
rlabel metal2 s 25900 -480 26012 240 8 wbs_adr_i[5]
port 570 nsew signal input
rlabel metal2 s 27580 -480 27692 240 8 wbs_adr_i[6]
port 571 nsew signal input
rlabel metal2 s 29260 -480 29372 240 8 wbs_adr_i[7]
port 572 nsew signal input
rlabel metal2 s 30940 -480 31052 240 8 wbs_adr_i[8]
port 573 nsew signal input
rlabel metal2 s 32620 -480 32732 240 8 wbs_adr_i[9]
port 574 nsew signal input
rlabel metal2 s 13580 -480 13692 240 8 wbs_cyc_i
port 575 nsew signal input
rlabel metal2 s 15820 -480 15932 240 8 wbs_dat_i[0]
port 576 nsew signal input
rlabel metal2 s 34860 -480 34972 240 8 wbs_dat_i[10]
port 577 nsew signal input
rlabel metal2 s 36540 -480 36652 240 8 wbs_dat_i[11]
port 578 nsew signal input
rlabel metal2 s 38220 -480 38332 240 8 wbs_dat_i[12]
port 579 nsew signal input
rlabel metal2 s 39900 -480 40012 240 8 wbs_dat_i[13]
port 580 nsew signal input
rlabel metal2 s 41580 -480 41692 240 8 wbs_dat_i[14]
port 581 nsew signal input
rlabel metal2 s 43260 -480 43372 240 8 wbs_dat_i[15]
port 582 nsew signal input
rlabel metal2 s 44940 -480 45052 240 8 wbs_dat_i[16]
port 583 nsew signal input
rlabel metal2 s 46620 -480 46732 240 8 wbs_dat_i[17]
port 584 nsew signal input
rlabel metal2 s 48300 -480 48412 240 8 wbs_dat_i[18]
port 585 nsew signal input
rlabel metal2 s 49980 -480 50092 240 8 wbs_dat_i[19]
port 586 nsew signal input
rlabel metal2 s 18060 -480 18172 240 8 wbs_dat_i[1]
port 587 nsew signal input
rlabel metal2 s 51660 -480 51772 240 8 wbs_dat_i[20]
port 588 nsew signal input
rlabel metal2 s 53340 -480 53452 240 8 wbs_dat_i[21]
port 589 nsew signal input
rlabel metal2 s 55020 -480 55132 240 8 wbs_dat_i[22]
port 590 nsew signal input
rlabel metal2 s 56700 -480 56812 240 8 wbs_dat_i[23]
port 591 nsew signal input
rlabel metal2 s 58380 -480 58492 240 8 wbs_dat_i[24]
port 592 nsew signal input
rlabel metal2 s 60060 -480 60172 240 8 wbs_dat_i[25]
port 593 nsew signal input
rlabel metal2 s 61740 -480 61852 240 8 wbs_dat_i[26]
port 594 nsew signal input
rlabel metal2 s 63420 -480 63532 240 8 wbs_dat_i[27]
port 595 nsew signal input
rlabel metal2 s 65100 -480 65212 240 8 wbs_dat_i[28]
port 596 nsew signal input
rlabel metal2 s 66780 -480 66892 240 8 wbs_dat_i[29]
port 597 nsew signal input
rlabel metal2 s 20300 -480 20412 240 8 wbs_dat_i[2]
port 598 nsew signal input
rlabel metal2 s 68460 -480 68572 240 8 wbs_dat_i[30]
port 599 nsew signal input
rlabel metal2 s 70140 -480 70252 240 8 wbs_dat_i[31]
port 600 nsew signal input
rlabel metal2 s 22540 -480 22652 240 8 wbs_dat_i[3]
port 601 nsew signal input
rlabel metal2 s 24780 -480 24892 240 8 wbs_dat_i[4]
port 602 nsew signal input
rlabel metal2 s 26460 -480 26572 240 8 wbs_dat_i[5]
port 603 nsew signal input
rlabel metal2 s 28140 -480 28252 240 8 wbs_dat_i[6]
port 604 nsew signal input
rlabel metal2 s 29820 -480 29932 240 8 wbs_dat_i[7]
port 605 nsew signal input
rlabel metal2 s 31500 -480 31612 240 8 wbs_dat_i[8]
port 606 nsew signal input
rlabel metal2 s 33180 -480 33292 240 8 wbs_dat_i[9]
port 607 nsew signal input
rlabel metal2 s 16380 -480 16492 240 8 wbs_dat_o[0]
port 608 nsew signal output
rlabel metal2 s 35420 -480 35532 240 8 wbs_dat_o[10]
port 609 nsew signal output
rlabel metal2 s 37100 -480 37212 240 8 wbs_dat_o[11]
port 610 nsew signal output
rlabel metal2 s 38780 -480 38892 240 8 wbs_dat_o[12]
port 611 nsew signal output
rlabel metal2 s 40460 -480 40572 240 8 wbs_dat_o[13]
port 612 nsew signal output
rlabel metal2 s 42140 -480 42252 240 8 wbs_dat_o[14]
port 613 nsew signal output
rlabel metal2 s 43820 -480 43932 240 8 wbs_dat_o[15]
port 614 nsew signal output
rlabel metal2 s 45500 -480 45612 240 8 wbs_dat_o[16]
port 615 nsew signal output
rlabel metal2 s 47180 -480 47292 240 8 wbs_dat_o[17]
port 616 nsew signal output
rlabel metal2 s 48860 -480 48972 240 8 wbs_dat_o[18]
port 617 nsew signal output
rlabel metal2 s 50540 -480 50652 240 8 wbs_dat_o[19]
port 618 nsew signal output
rlabel metal2 s 18620 -480 18732 240 8 wbs_dat_o[1]
port 619 nsew signal output
rlabel metal2 s 52220 -480 52332 240 8 wbs_dat_o[20]
port 620 nsew signal output
rlabel metal2 s 53900 -480 54012 240 8 wbs_dat_o[21]
port 621 nsew signal output
rlabel metal2 s 55580 -480 55692 240 8 wbs_dat_o[22]
port 622 nsew signal output
rlabel metal2 s 57260 -480 57372 240 8 wbs_dat_o[23]
port 623 nsew signal output
rlabel metal2 s 58940 -480 59052 240 8 wbs_dat_o[24]
port 624 nsew signal output
rlabel metal2 s 60620 -480 60732 240 8 wbs_dat_o[25]
port 625 nsew signal output
rlabel metal2 s 62300 -480 62412 240 8 wbs_dat_o[26]
port 626 nsew signal output
rlabel metal2 s 63980 -480 64092 240 8 wbs_dat_o[27]
port 627 nsew signal output
rlabel metal2 s 65660 -480 65772 240 8 wbs_dat_o[28]
port 628 nsew signal output
rlabel metal2 s 67340 -480 67452 240 8 wbs_dat_o[29]
port 629 nsew signal output
rlabel metal2 s 20860 -480 20972 240 8 wbs_dat_o[2]
port 630 nsew signal output
rlabel metal2 s 69020 -480 69132 240 8 wbs_dat_o[30]
port 631 nsew signal output
rlabel metal2 s 70700 -480 70812 240 8 wbs_dat_o[31]
port 632 nsew signal output
rlabel metal2 s 23100 -480 23212 240 8 wbs_dat_o[3]
port 633 nsew signal output
rlabel metal2 s 25340 -480 25452 240 8 wbs_dat_o[4]
port 634 nsew signal output
rlabel metal2 s 27020 -480 27132 240 8 wbs_dat_o[5]
port 635 nsew signal output
rlabel metal2 s 28700 -480 28812 240 8 wbs_dat_o[6]
port 636 nsew signal output
rlabel metal2 s 30380 -480 30492 240 8 wbs_dat_o[7]
port 637 nsew signal output
rlabel metal2 s 32060 -480 32172 240 8 wbs_dat_o[8]
port 638 nsew signal output
rlabel metal2 s 33740 -480 33852 240 8 wbs_dat_o[9]
port 639 nsew signal output
rlabel metal2 s 16940 -480 17052 240 8 wbs_sel_i[0]
port 640 nsew signal input
rlabel metal2 s 19180 -480 19292 240 8 wbs_sel_i[1]
port 641 nsew signal input
rlabel metal2 s 21420 -480 21532 240 8 wbs_sel_i[2]
port 642 nsew signal input
rlabel metal2 s 23660 -480 23772 240 8 wbs_sel_i[3]
port 643 nsew signal input
rlabel metal2 s 14140 -480 14252 240 8 wbs_stb_i
port 644 nsew signal input
rlabel metal2 s 14700 -480 14812 240 8 wbs_we_i
port 645 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 300000 300000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 26724796
string GDS_FILE /home/jasteve4/Documents/MicroMotorController/openlane/user_project_wrapper/runs/22_12_05_15_21/results/signoff/user_project_wrapper.magic.gds
string GDS_START 23184140
<< end >>


magic
tech gf180mcuC
magscale 1 10
timestamp 1670279885
<< metal1 >>
rect 1344 46282 48608 46316
rect 1344 46230 2058 46282
rect 2110 46230 2162 46282
rect 2214 46230 2266 46282
rect 2318 46230 2370 46282
rect 2422 46230 2474 46282
rect 2526 46230 2578 46282
rect 2630 46230 38058 46282
rect 38110 46230 38162 46282
rect 38214 46230 38266 46282
rect 38318 46230 38370 46282
rect 38422 46230 38474 46282
rect 38526 46230 38578 46282
rect 38630 46230 48608 46282
rect 1344 46196 48608 46230
rect 1822 46114 1874 46126
rect 1822 46050 1874 46062
rect 46050 45950 46062 46002
rect 46114 45950 46126 46002
rect 45042 45838 45054 45890
rect 45106 45838 45118 45890
rect 46834 45838 46846 45890
rect 46898 45838 46910 45890
rect 47730 45726 47742 45778
rect 47794 45726 47806 45778
rect 44158 45666 44210 45678
rect 44158 45602 44210 45614
rect 1344 45498 48608 45532
rect 1344 45446 5778 45498
rect 5830 45446 5882 45498
rect 5934 45446 5986 45498
rect 6038 45446 6090 45498
rect 6142 45446 6194 45498
rect 6246 45446 6298 45498
rect 6350 45446 41778 45498
rect 41830 45446 41882 45498
rect 41934 45446 41986 45498
rect 42038 45446 42090 45498
rect 42142 45446 42194 45498
rect 42246 45446 42298 45498
rect 42350 45446 48608 45498
rect 1344 45412 48608 45446
rect 45838 45330 45890 45342
rect 45838 45266 45890 45278
rect 46834 45054 46846 45106
rect 46898 45054 46910 45106
rect 46398 44994 46450 45006
rect 47842 44942 47854 44994
rect 47906 44942 47918 44994
rect 46398 44930 46450 44942
rect 1344 44714 48608 44748
rect 1344 44662 2058 44714
rect 2110 44662 2162 44714
rect 2214 44662 2266 44714
rect 2318 44662 2370 44714
rect 2422 44662 2474 44714
rect 2526 44662 2578 44714
rect 2630 44662 38058 44714
rect 38110 44662 38162 44714
rect 38214 44662 38266 44714
rect 38318 44662 38370 44714
rect 38422 44662 38474 44714
rect 38526 44662 38578 44714
rect 38630 44662 48608 44714
rect 1344 44628 48608 44662
rect 46286 44322 46338 44334
rect 46834 44270 46846 44322
rect 46898 44270 46910 44322
rect 46286 44258 46338 44270
rect 47730 44158 47742 44210
rect 47794 44158 47806 44210
rect 1344 43930 48608 43964
rect 1344 43878 5778 43930
rect 5830 43878 5882 43930
rect 5934 43878 5986 43930
rect 6038 43878 6090 43930
rect 6142 43878 6194 43930
rect 6246 43878 6298 43930
rect 6350 43878 41778 43930
rect 41830 43878 41882 43930
rect 41934 43878 41986 43930
rect 42038 43878 42090 43930
rect 42142 43878 42194 43930
rect 42246 43878 42298 43930
rect 42350 43878 48608 43930
rect 1344 43844 48608 43878
rect 1344 43146 48608 43180
rect 1344 43094 2058 43146
rect 2110 43094 2162 43146
rect 2214 43094 2266 43146
rect 2318 43094 2370 43146
rect 2422 43094 2474 43146
rect 2526 43094 2578 43146
rect 2630 43094 38058 43146
rect 38110 43094 38162 43146
rect 38214 43094 38266 43146
rect 38318 43094 38370 43146
rect 38422 43094 38474 43146
rect 38526 43094 38578 43146
rect 38630 43094 48608 43146
rect 1344 43060 48608 43094
rect 46834 42702 46846 42754
rect 46898 42702 46910 42754
rect 47730 42590 47742 42642
rect 47794 42590 47806 42642
rect 46286 42530 46338 42542
rect 46286 42466 46338 42478
rect 1344 42362 48608 42396
rect 1344 42310 5778 42362
rect 5830 42310 5882 42362
rect 5934 42310 5986 42362
rect 6038 42310 6090 42362
rect 6142 42310 6194 42362
rect 6246 42310 6298 42362
rect 6350 42310 41778 42362
rect 41830 42310 41882 42362
rect 41934 42310 41986 42362
rect 42038 42310 42090 42362
rect 42142 42310 42194 42362
rect 42246 42310 42298 42362
rect 42350 42310 48608 42362
rect 1344 42276 48608 42310
rect 1344 41578 48608 41612
rect 1344 41526 2058 41578
rect 2110 41526 2162 41578
rect 2214 41526 2266 41578
rect 2318 41526 2370 41578
rect 2422 41526 2474 41578
rect 2526 41526 2578 41578
rect 2630 41526 38058 41578
rect 38110 41526 38162 41578
rect 38214 41526 38266 41578
rect 38318 41526 38370 41578
rect 38422 41526 38474 41578
rect 38526 41526 38578 41578
rect 38630 41526 48608 41578
rect 1344 41492 48608 41526
rect 3042 41134 3054 41186
rect 3106 41134 3118 41186
rect 46834 41134 46846 41186
rect 46898 41134 46910 41186
rect 2146 41022 2158 41074
rect 2210 41022 2222 41074
rect 47730 41022 47742 41074
rect 47794 41022 47806 41074
rect 3502 40962 3554 40974
rect 3502 40898 3554 40910
rect 46286 40962 46338 40974
rect 46286 40898 46338 40910
rect 1344 40794 48608 40828
rect 1344 40742 5778 40794
rect 5830 40742 5882 40794
rect 5934 40742 5986 40794
rect 6038 40742 6090 40794
rect 6142 40742 6194 40794
rect 6246 40742 6298 40794
rect 6350 40742 41778 40794
rect 41830 40742 41882 40794
rect 41934 40742 41986 40794
rect 42038 40742 42090 40794
rect 42142 40742 42194 40794
rect 42246 40742 42298 40794
rect 42350 40742 48608 40794
rect 1344 40708 48608 40742
rect 1344 40010 48608 40044
rect 1344 39958 2058 40010
rect 2110 39958 2162 40010
rect 2214 39958 2266 40010
rect 2318 39958 2370 40010
rect 2422 39958 2474 40010
rect 2526 39958 2578 40010
rect 2630 39958 38058 40010
rect 38110 39958 38162 40010
rect 38214 39958 38266 40010
rect 38318 39958 38370 40010
rect 38422 39958 38474 40010
rect 38526 39958 38578 40010
rect 38630 39958 48608 40010
rect 1344 39924 48608 39958
rect 46834 39566 46846 39618
rect 46898 39566 46910 39618
rect 47730 39454 47742 39506
rect 47794 39454 47806 39506
rect 46286 39394 46338 39406
rect 46286 39330 46338 39342
rect 1344 39226 48608 39260
rect 1344 39174 5778 39226
rect 5830 39174 5882 39226
rect 5934 39174 5986 39226
rect 6038 39174 6090 39226
rect 6142 39174 6194 39226
rect 6246 39174 6298 39226
rect 6350 39174 41778 39226
rect 41830 39174 41882 39226
rect 41934 39174 41986 39226
rect 42038 39174 42090 39226
rect 42142 39174 42194 39226
rect 42246 39174 42298 39226
rect 42350 39174 48608 39226
rect 1344 39140 48608 39174
rect 46834 38782 46846 38834
rect 46898 38782 46910 38834
rect 46398 38722 46450 38734
rect 47842 38670 47854 38722
rect 47906 38670 47918 38722
rect 46398 38658 46450 38670
rect 1344 38442 48608 38476
rect 1344 38390 2058 38442
rect 2110 38390 2162 38442
rect 2214 38390 2266 38442
rect 2318 38390 2370 38442
rect 2422 38390 2474 38442
rect 2526 38390 2578 38442
rect 2630 38390 38058 38442
rect 38110 38390 38162 38442
rect 38214 38390 38266 38442
rect 38318 38390 38370 38442
rect 38422 38390 38474 38442
rect 38526 38390 38578 38442
rect 38630 38390 48608 38442
rect 1344 38356 48608 38390
rect 1344 37658 48608 37692
rect 1344 37606 5778 37658
rect 5830 37606 5882 37658
rect 5934 37606 5986 37658
rect 6038 37606 6090 37658
rect 6142 37606 6194 37658
rect 6246 37606 6298 37658
rect 6350 37606 41778 37658
rect 41830 37606 41882 37658
rect 41934 37606 41986 37658
rect 42038 37606 42090 37658
rect 42142 37606 42194 37658
rect 42246 37606 42298 37658
rect 42350 37606 48608 37658
rect 1344 37572 48608 37606
rect 46834 37214 46846 37266
rect 46898 37214 46910 37266
rect 46398 37154 46450 37166
rect 47842 37102 47854 37154
rect 47906 37102 47918 37154
rect 46398 37090 46450 37102
rect 1344 36874 48608 36908
rect 1344 36822 2058 36874
rect 2110 36822 2162 36874
rect 2214 36822 2266 36874
rect 2318 36822 2370 36874
rect 2422 36822 2474 36874
rect 2526 36822 2578 36874
rect 2630 36822 38058 36874
rect 38110 36822 38162 36874
rect 38214 36822 38266 36874
rect 38318 36822 38370 36874
rect 38422 36822 38474 36874
rect 38526 36822 38578 36874
rect 38630 36822 48608 36874
rect 1344 36788 48608 36822
rect 17950 36370 18002 36382
rect 17950 36306 18002 36318
rect 18286 36370 18338 36382
rect 18286 36306 18338 36318
rect 17390 36258 17442 36270
rect 17390 36194 17442 36206
rect 1344 36090 48608 36124
rect 1344 36038 5778 36090
rect 5830 36038 5882 36090
rect 5934 36038 5986 36090
rect 6038 36038 6090 36090
rect 6142 36038 6194 36090
rect 6246 36038 6298 36090
rect 6350 36038 41778 36090
rect 41830 36038 41882 36090
rect 41934 36038 41986 36090
rect 42038 36038 42090 36090
rect 42142 36038 42194 36090
rect 42246 36038 42298 36090
rect 42350 36038 48608 36090
rect 1344 36004 48608 36038
rect 46398 35698 46450 35710
rect 46946 35646 46958 35698
rect 47010 35646 47022 35698
rect 46398 35634 46450 35646
rect 47842 35534 47854 35586
rect 47906 35534 47918 35586
rect 1344 35306 48608 35340
rect 1344 35254 2058 35306
rect 2110 35254 2162 35306
rect 2214 35254 2266 35306
rect 2318 35254 2370 35306
rect 2422 35254 2474 35306
rect 2526 35254 2578 35306
rect 2630 35254 38058 35306
rect 38110 35254 38162 35306
rect 38214 35254 38266 35306
rect 38318 35254 38370 35306
rect 38422 35254 38474 35306
rect 38526 35254 38578 35306
rect 38630 35254 48608 35306
rect 1344 35220 48608 35254
rect 1822 34690 1874 34702
rect 1822 34626 1874 34638
rect 1344 34522 48608 34556
rect 1344 34470 5778 34522
rect 5830 34470 5882 34522
rect 5934 34470 5986 34522
rect 6038 34470 6090 34522
rect 6142 34470 6194 34522
rect 6246 34470 6298 34522
rect 6350 34470 41778 34522
rect 41830 34470 41882 34522
rect 41934 34470 41986 34522
rect 42038 34470 42090 34522
rect 42142 34470 42194 34522
rect 42246 34470 42298 34522
rect 42350 34470 48608 34522
rect 1344 34436 48608 34470
rect 46946 34078 46958 34130
rect 47010 34078 47022 34130
rect 46398 34018 46450 34030
rect 46834 34015 46846 34018
rect 46398 33954 46450 33966
rect 46625 33969 46846 34015
rect 46274 33854 46286 33906
rect 46338 33903 46350 33906
rect 46625 33903 46671 33969
rect 46834 33966 46846 33969
rect 46898 33966 46910 34018
rect 47842 33966 47854 34018
rect 47906 33966 47918 34018
rect 46338 33857 46671 33903
rect 46338 33854 46350 33857
rect 1344 33738 48608 33772
rect 1344 33686 2058 33738
rect 2110 33686 2162 33738
rect 2214 33686 2266 33738
rect 2318 33686 2370 33738
rect 2422 33686 2474 33738
rect 2526 33686 2578 33738
rect 2630 33686 38058 33738
rect 38110 33686 38162 33738
rect 38214 33686 38266 33738
rect 38318 33686 38370 33738
rect 38422 33686 38474 33738
rect 38526 33686 38578 33738
rect 38630 33686 48608 33738
rect 1344 33652 48608 33686
rect 1344 32954 48608 32988
rect 1344 32902 5778 32954
rect 5830 32902 5882 32954
rect 5934 32902 5986 32954
rect 6038 32902 6090 32954
rect 6142 32902 6194 32954
rect 6246 32902 6298 32954
rect 6350 32902 41778 32954
rect 41830 32902 41882 32954
rect 41934 32902 41986 32954
rect 42038 32902 42090 32954
rect 42142 32902 42194 32954
rect 42246 32902 42298 32954
rect 42350 32902 48608 32954
rect 1344 32868 48608 32902
rect 46834 32510 46846 32562
rect 46898 32510 46910 32562
rect 46398 32450 46450 32462
rect 47842 32398 47854 32450
rect 47906 32398 47918 32450
rect 46398 32386 46450 32398
rect 1344 32170 48608 32204
rect 1344 32118 2058 32170
rect 2110 32118 2162 32170
rect 2214 32118 2266 32170
rect 2318 32118 2370 32170
rect 2422 32118 2474 32170
rect 2526 32118 2578 32170
rect 2630 32118 38058 32170
rect 38110 32118 38162 32170
rect 38214 32118 38266 32170
rect 38318 32118 38370 32170
rect 38422 32118 38474 32170
rect 38526 32118 38578 32170
rect 38630 32118 48608 32170
rect 1344 32084 48608 32118
rect 1344 31386 48608 31420
rect 1344 31334 5778 31386
rect 5830 31334 5882 31386
rect 5934 31334 5986 31386
rect 6038 31334 6090 31386
rect 6142 31334 6194 31386
rect 6246 31334 6298 31386
rect 6350 31334 41778 31386
rect 41830 31334 41882 31386
rect 41934 31334 41986 31386
rect 42038 31334 42090 31386
rect 42142 31334 42194 31386
rect 42246 31334 42298 31386
rect 42350 31334 48608 31386
rect 1344 31300 48608 31334
rect 46398 30994 46450 31006
rect 46946 30942 46958 30994
rect 47010 30942 47022 30994
rect 46398 30930 46450 30942
rect 46498 30830 46510 30882
rect 46562 30879 46574 30882
rect 46834 30879 46846 30882
rect 46562 30833 46846 30879
rect 46562 30830 46574 30833
rect 46834 30830 46846 30833
rect 46898 30830 46910 30882
rect 47842 30830 47854 30882
rect 47906 30830 47918 30882
rect 1344 30602 48608 30636
rect 1344 30550 2058 30602
rect 2110 30550 2162 30602
rect 2214 30550 2266 30602
rect 2318 30550 2370 30602
rect 2422 30550 2474 30602
rect 2526 30550 2578 30602
rect 2630 30550 38058 30602
rect 38110 30550 38162 30602
rect 38214 30550 38266 30602
rect 38318 30550 38370 30602
rect 38422 30550 38474 30602
rect 38526 30550 38578 30602
rect 38630 30550 48608 30602
rect 1344 30516 48608 30550
rect 1344 29818 48608 29852
rect 1344 29766 5778 29818
rect 5830 29766 5882 29818
rect 5934 29766 5986 29818
rect 6038 29766 6090 29818
rect 6142 29766 6194 29818
rect 6246 29766 6298 29818
rect 6350 29766 41778 29818
rect 41830 29766 41882 29818
rect 41934 29766 41986 29818
rect 42038 29766 42090 29818
rect 42142 29766 42194 29818
rect 42246 29766 42298 29818
rect 42350 29766 48608 29818
rect 1344 29732 48608 29766
rect 38994 29486 39006 29538
rect 39058 29486 39070 29538
rect 38334 29426 38386 29438
rect 38770 29374 38782 29426
rect 38834 29374 38846 29426
rect 46834 29374 46846 29426
rect 46898 29374 46910 29426
rect 38334 29362 38386 29374
rect 36878 29314 36930 29326
rect 36878 29250 36930 29262
rect 37326 29314 37378 29326
rect 37326 29250 37378 29262
rect 39678 29314 39730 29326
rect 39678 29250 39730 29262
rect 46398 29314 46450 29326
rect 47842 29262 47854 29314
rect 47906 29262 47918 29314
rect 46398 29250 46450 29262
rect 37998 29202 38050 29214
rect 37998 29138 38050 29150
rect 1344 29034 48608 29068
rect 1344 28982 2058 29034
rect 2110 28982 2162 29034
rect 2214 28982 2266 29034
rect 2318 28982 2370 29034
rect 2422 28982 2474 29034
rect 2526 28982 2578 29034
rect 2630 28982 38058 29034
rect 38110 28982 38162 29034
rect 38214 28982 38266 29034
rect 38318 28982 38370 29034
rect 38422 28982 38474 29034
rect 38526 28982 38578 29034
rect 38630 28982 48608 29034
rect 1344 28948 48608 28982
rect 39666 28814 39678 28866
rect 39730 28863 39742 28866
rect 40226 28863 40238 28866
rect 39730 28817 40238 28863
rect 39730 28814 39742 28817
rect 40226 28814 40238 28817
rect 40290 28814 40302 28866
rect 36766 28754 36818 28766
rect 36766 28690 36818 28702
rect 38334 28754 38386 28766
rect 47842 28702 47854 28754
rect 47906 28702 47918 28754
rect 38334 28690 38386 28702
rect 37998 28642 38050 28654
rect 37998 28578 38050 28590
rect 46286 28642 46338 28654
rect 46834 28590 46846 28642
rect 46898 28590 46910 28642
rect 46286 28578 46338 28590
rect 1822 28530 1874 28542
rect 40126 28530 40178 28542
rect 38546 28478 38558 28530
rect 38610 28478 38622 28530
rect 38882 28478 38894 28530
rect 38946 28478 38958 28530
rect 1822 28466 1874 28478
rect 40126 28466 40178 28478
rect 2158 28418 2210 28430
rect 2158 28354 2210 28366
rect 39678 28418 39730 28430
rect 39678 28354 39730 28366
rect 1344 28250 48608 28284
rect 1344 28198 5778 28250
rect 5830 28198 5882 28250
rect 5934 28198 5986 28250
rect 6038 28198 6090 28250
rect 6142 28198 6194 28250
rect 6246 28198 6298 28250
rect 6350 28198 41778 28250
rect 41830 28198 41882 28250
rect 41934 28198 41986 28250
rect 42038 28198 42090 28250
rect 42142 28198 42194 28250
rect 42246 28198 42298 28250
rect 42350 28198 48608 28250
rect 1344 28164 48608 28198
rect 1822 28082 1874 28094
rect 1822 28018 1874 28030
rect 36654 28082 36706 28094
rect 36654 28018 36706 28030
rect 38210 27918 38222 27970
rect 38274 27918 38286 27970
rect 37662 27858 37714 27870
rect 39118 27858 39170 27870
rect 38098 27806 38110 27858
rect 38162 27806 38174 27858
rect 37662 27794 37714 27806
rect 39118 27794 39170 27806
rect 39678 27858 39730 27870
rect 39678 27794 39730 27806
rect 36206 27746 36258 27758
rect 36206 27682 36258 27694
rect 37326 27634 37378 27646
rect 37326 27570 37378 27582
rect 1344 27466 48608 27500
rect 1344 27414 2058 27466
rect 2110 27414 2162 27466
rect 2214 27414 2266 27466
rect 2318 27414 2370 27466
rect 2422 27414 2474 27466
rect 2526 27414 2578 27466
rect 2630 27414 38058 27466
rect 38110 27414 38162 27466
rect 38214 27414 38266 27466
rect 38318 27414 38370 27466
rect 38422 27414 38474 27466
rect 38526 27414 38578 27466
rect 38630 27414 48608 27466
rect 1344 27380 48608 27414
rect 38782 27186 38834 27198
rect 38782 27122 38834 27134
rect 46834 27022 46846 27074
rect 46898 27022 46910 27074
rect 39678 26962 39730 26974
rect 39678 26898 39730 26910
rect 46286 26962 46338 26974
rect 47730 26910 47742 26962
rect 47794 26910 47806 26962
rect 46286 26898 46338 26910
rect 40238 26850 40290 26862
rect 40238 26786 40290 26798
rect 1344 26682 48608 26716
rect 1344 26630 5778 26682
rect 5830 26630 5882 26682
rect 5934 26630 5986 26682
rect 6038 26630 6090 26682
rect 6142 26630 6194 26682
rect 6246 26630 6298 26682
rect 6350 26630 41778 26682
rect 41830 26630 41882 26682
rect 41934 26630 41986 26682
rect 42038 26630 42090 26682
rect 42142 26630 42194 26682
rect 42246 26630 42298 26682
rect 42350 26630 48608 26682
rect 1344 26596 48608 26630
rect 39106 26350 39118 26402
rect 39170 26350 39182 26402
rect 39330 26238 39342 26290
rect 39394 26238 39406 26290
rect 37102 26178 37154 26190
rect 37102 26114 37154 26126
rect 37550 26178 37602 26190
rect 37550 26114 37602 26126
rect 38558 26178 38610 26190
rect 38558 26114 38610 26126
rect 38222 26066 38274 26078
rect 38222 26002 38274 26014
rect 1344 25898 48608 25932
rect 1344 25846 2058 25898
rect 2110 25846 2162 25898
rect 2214 25846 2266 25898
rect 2318 25846 2370 25898
rect 2422 25846 2474 25898
rect 2526 25846 2578 25898
rect 2630 25846 38058 25898
rect 38110 25846 38162 25898
rect 38214 25846 38266 25898
rect 38318 25846 38370 25898
rect 38422 25846 38474 25898
rect 38526 25846 38578 25898
rect 38630 25846 48608 25898
rect 1344 25812 48608 25846
rect 40338 25566 40350 25618
rect 40402 25566 40414 25618
rect 46946 25454 46958 25506
rect 47010 25454 47022 25506
rect 47730 25342 47742 25394
rect 47794 25342 47806 25394
rect 40798 25282 40850 25294
rect 40798 25218 40850 25230
rect 46286 25282 46338 25294
rect 46286 25218 46338 25230
rect 1344 25114 48608 25148
rect 1344 25062 5778 25114
rect 5830 25062 5882 25114
rect 5934 25062 5986 25114
rect 6038 25062 6090 25114
rect 6142 25062 6194 25114
rect 6246 25062 6298 25114
rect 6350 25062 41778 25114
rect 41830 25062 41882 25114
rect 41934 25062 41986 25114
rect 42038 25062 42090 25114
rect 42142 25062 42194 25114
rect 42246 25062 42298 25114
rect 42350 25062 48608 25114
rect 1344 25028 48608 25062
rect 39106 24782 39118 24834
rect 39170 24782 39182 24834
rect 38446 24722 38498 24734
rect 39218 24670 39230 24722
rect 39282 24670 39294 24722
rect 38446 24658 38498 24670
rect 36990 24610 37042 24622
rect 36990 24546 37042 24558
rect 37438 24610 37490 24622
rect 37438 24546 37490 24558
rect 38110 24498 38162 24510
rect 38110 24434 38162 24446
rect 1344 24330 48608 24364
rect 1344 24278 2058 24330
rect 2110 24278 2162 24330
rect 2214 24278 2266 24330
rect 2318 24278 2370 24330
rect 2422 24278 2474 24330
rect 2526 24278 2578 24330
rect 2630 24278 38058 24330
rect 38110 24278 38162 24330
rect 38214 24278 38266 24330
rect 38318 24278 38370 24330
rect 38422 24278 38474 24330
rect 38526 24278 38578 24330
rect 38630 24278 48608 24330
rect 1344 24244 48608 24278
rect 39678 24050 39730 24062
rect 39678 23986 39730 23998
rect 38334 23938 38386 23950
rect 39106 23886 39118 23938
rect 39170 23886 39182 23938
rect 40786 23886 40798 23938
rect 40850 23886 40862 23938
rect 46834 23886 46846 23938
rect 46898 23886 46910 23938
rect 38334 23874 38386 23886
rect 40350 23826 40402 23838
rect 38994 23774 39006 23826
rect 39058 23774 39070 23826
rect 47730 23774 47742 23826
rect 47794 23774 47806 23826
rect 40350 23762 40402 23774
rect 36766 23714 36818 23726
rect 36766 23650 36818 23662
rect 37998 23714 38050 23726
rect 37998 23650 38050 23662
rect 46286 23714 46338 23726
rect 46286 23650 46338 23662
rect 1344 23546 48608 23580
rect 1344 23494 5778 23546
rect 5830 23494 5882 23546
rect 5934 23494 5986 23546
rect 6038 23494 6090 23546
rect 6142 23494 6194 23546
rect 6246 23494 6298 23546
rect 6350 23494 41778 23546
rect 41830 23494 41882 23546
rect 41934 23494 41986 23546
rect 42038 23494 42090 23546
rect 42142 23494 42194 23546
rect 42246 23494 42298 23546
rect 42350 23494 48608 23546
rect 1344 23460 48608 23494
rect 38994 23214 39006 23266
rect 39058 23214 39070 23266
rect 39106 23102 39118 23154
rect 39170 23102 39182 23154
rect 36878 23042 36930 23054
rect 36878 22978 36930 22990
rect 37326 23042 37378 23054
rect 37326 22978 37378 22990
rect 37998 22930 38050 22942
rect 37998 22866 38050 22878
rect 38334 22930 38386 22942
rect 38334 22866 38386 22878
rect 1344 22762 48608 22796
rect 1344 22710 2058 22762
rect 2110 22710 2162 22762
rect 2214 22710 2266 22762
rect 2318 22710 2370 22762
rect 2422 22710 2474 22762
rect 2526 22710 2578 22762
rect 2630 22710 38058 22762
rect 38110 22710 38162 22762
rect 38214 22710 38266 22762
rect 38318 22710 38370 22762
rect 38422 22710 38474 22762
rect 38526 22710 38578 22762
rect 38630 22710 48608 22762
rect 1344 22676 48608 22710
rect 46834 22318 46846 22370
rect 46898 22318 46910 22370
rect 28366 22258 28418 22270
rect 28366 22194 28418 22206
rect 38110 22258 38162 22270
rect 38110 22194 38162 22206
rect 38670 22258 38722 22270
rect 47730 22206 47742 22258
rect 47794 22206 47806 22258
rect 38670 22194 38722 22206
rect 1822 22146 1874 22158
rect 1822 22082 1874 22094
rect 28030 22146 28082 22158
rect 28030 22082 28082 22094
rect 38222 22146 38274 22158
rect 38222 22082 38274 22094
rect 46286 22146 46338 22158
rect 46286 22082 46338 22094
rect 1344 21978 48608 22012
rect 1344 21926 5778 21978
rect 5830 21926 5882 21978
rect 5934 21926 5986 21978
rect 6038 21926 6090 21978
rect 6142 21926 6194 21978
rect 6246 21926 6298 21978
rect 6350 21926 41778 21978
rect 41830 21926 41882 21978
rect 41934 21926 41986 21978
rect 42038 21926 42090 21978
rect 42142 21926 42194 21978
rect 42246 21926 42298 21978
rect 42350 21926 48608 21978
rect 1344 21892 48608 21926
rect 38434 21646 38446 21698
rect 38498 21646 38510 21698
rect 38658 21534 38670 21586
rect 38722 21534 38734 21586
rect 36430 21474 36482 21486
rect 36430 21410 36482 21422
rect 36878 21474 36930 21486
rect 36878 21410 36930 21422
rect 37550 21362 37602 21374
rect 37550 21298 37602 21310
rect 37886 21362 37938 21374
rect 37886 21298 37938 21310
rect 1344 21194 48608 21228
rect 1344 21142 2058 21194
rect 2110 21142 2162 21194
rect 2214 21142 2266 21194
rect 2318 21142 2370 21194
rect 2422 21142 2474 21194
rect 2526 21142 2578 21194
rect 2630 21142 38058 21194
rect 38110 21142 38162 21194
rect 38214 21142 38266 21194
rect 38318 21142 38370 21194
rect 38422 21142 38474 21194
rect 38526 21142 38578 21194
rect 38630 21142 48608 21194
rect 1344 21108 48608 21142
rect 29822 21026 29874 21038
rect 29822 20962 29874 20974
rect 37998 21026 38050 21038
rect 37998 20962 38050 20974
rect 31502 20914 31554 20926
rect 31502 20850 31554 20862
rect 36766 20914 36818 20926
rect 36766 20850 36818 20862
rect 30158 20802 30210 20814
rect 30930 20750 30942 20802
rect 30994 20750 31006 20802
rect 38770 20750 38782 20802
rect 38834 20750 38846 20802
rect 46834 20750 46846 20802
rect 46898 20750 46910 20802
rect 30158 20738 30210 20750
rect 33518 20690 33570 20702
rect 39454 20690 39506 20702
rect 30818 20638 30830 20690
rect 30882 20638 30894 20690
rect 38658 20638 38670 20690
rect 38722 20638 38734 20690
rect 33518 20626 33570 20638
rect 39454 20626 39506 20638
rect 39902 20690 39954 20702
rect 39902 20626 39954 20638
rect 40014 20690 40066 20702
rect 40014 20626 40066 20638
rect 40462 20690 40514 20702
rect 40462 20626 40514 20638
rect 40798 20690 40850 20702
rect 47730 20638 47742 20690
rect 47794 20638 47806 20690
rect 40798 20626 40850 20638
rect 28814 20578 28866 20590
rect 28814 20514 28866 20526
rect 33182 20578 33234 20590
rect 33182 20514 33234 20526
rect 36318 20578 36370 20590
rect 36318 20514 36370 20526
rect 37662 20578 37714 20590
rect 37662 20514 37714 20526
rect 39678 20578 39730 20590
rect 39678 20514 39730 20526
rect 46286 20578 46338 20590
rect 46286 20514 46338 20526
rect 1344 20410 48608 20444
rect 1344 20358 5778 20410
rect 5830 20358 5882 20410
rect 5934 20358 5986 20410
rect 6038 20358 6090 20410
rect 6142 20358 6194 20410
rect 6246 20358 6298 20410
rect 6350 20358 41778 20410
rect 41830 20358 41882 20410
rect 41934 20358 41986 20410
rect 42038 20358 42090 20410
rect 42142 20358 42194 20410
rect 42246 20358 42298 20410
rect 42350 20358 48608 20410
rect 1344 20324 48608 20358
rect 33630 20242 33682 20254
rect 33630 20178 33682 20190
rect 29374 20130 29426 20142
rect 29374 20066 29426 20078
rect 32286 20130 32338 20142
rect 32286 20066 32338 20078
rect 34526 20130 34578 20142
rect 37986 20078 37998 20130
rect 38050 20078 38062 20130
rect 34526 20066 34578 20078
rect 32622 20018 32674 20030
rect 32622 19954 32674 19966
rect 33966 20018 34018 20030
rect 37438 20018 37490 20030
rect 34738 19966 34750 20018
rect 34802 19966 34814 20018
rect 38210 19966 38222 20018
rect 38274 19966 38286 20018
rect 33966 19954 34018 19966
rect 37438 19954 37490 19966
rect 35982 19906 36034 19918
rect 35982 19842 36034 19854
rect 36430 19906 36482 19918
rect 36430 19842 36482 19854
rect 39118 19906 39170 19918
rect 39118 19842 39170 19854
rect 37102 19794 37154 19806
rect 37102 19730 37154 19742
rect 1344 19626 48608 19660
rect 1344 19574 2058 19626
rect 2110 19574 2162 19626
rect 2214 19574 2266 19626
rect 2318 19574 2370 19626
rect 2422 19574 2474 19626
rect 2526 19574 2578 19626
rect 2630 19574 38058 19626
rect 38110 19574 38162 19626
rect 38214 19574 38266 19626
rect 38318 19574 38370 19626
rect 38422 19574 38474 19626
rect 38526 19574 38578 19626
rect 38630 19574 48608 19626
rect 1344 19540 48608 19574
rect 34302 19458 34354 19470
rect 34302 19394 34354 19406
rect 37998 19458 38050 19470
rect 37998 19394 38050 19406
rect 36766 19346 36818 19358
rect 36766 19282 36818 19294
rect 38658 19182 38670 19234
rect 38722 19182 38734 19234
rect 46834 19182 46846 19234
rect 46898 19182 46910 19234
rect 31278 19122 31330 19134
rect 31278 19058 31330 19070
rect 34190 19122 34242 19134
rect 34190 19058 34242 19070
rect 37662 19122 37714 19134
rect 38770 19070 38782 19122
rect 38834 19070 38846 19122
rect 47730 19070 47742 19122
rect 47794 19070 47806 19122
rect 37662 19058 37714 19070
rect 30942 19010 30994 19022
rect 30942 18946 30994 18958
rect 33742 19010 33794 19022
rect 33742 18946 33794 18958
rect 34302 19010 34354 19022
rect 34302 18946 34354 18958
rect 34862 19010 34914 19022
rect 34862 18946 34914 18958
rect 35758 19010 35810 19022
rect 35758 18946 35810 18958
rect 36206 19010 36258 19022
rect 36206 18946 36258 18958
rect 46286 19010 46338 19022
rect 46286 18946 46338 18958
rect 1344 18842 48608 18876
rect 1344 18790 5778 18842
rect 5830 18790 5882 18842
rect 5934 18790 5986 18842
rect 6038 18790 6090 18842
rect 6142 18790 6194 18842
rect 6246 18790 6298 18842
rect 6350 18790 41778 18842
rect 41830 18790 41882 18842
rect 41934 18790 41986 18842
rect 42038 18790 42090 18842
rect 42142 18790 42194 18842
rect 42246 18790 42298 18842
rect 42350 18790 48608 18842
rect 1344 18756 48608 18790
rect 30046 18674 30098 18686
rect 30046 18610 30098 18622
rect 29150 18562 29202 18574
rect 29150 18498 29202 18510
rect 29486 18562 29538 18574
rect 29486 18498 29538 18510
rect 30942 18562 30994 18574
rect 30942 18498 30994 18510
rect 31278 18562 31330 18574
rect 31278 18498 31330 18510
rect 31838 18562 31890 18574
rect 31838 18498 31890 18510
rect 32174 18562 32226 18574
rect 32174 18498 32226 18510
rect 35422 18562 35474 18574
rect 37314 18510 37326 18562
rect 37378 18510 37390 18562
rect 35422 18498 35474 18510
rect 34862 18450 34914 18462
rect 36766 18450 36818 18462
rect 38110 18450 38162 18462
rect 35634 18398 35646 18450
rect 35698 18398 35710 18450
rect 37538 18398 37550 18450
rect 37602 18398 37614 18450
rect 34862 18386 34914 18398
rect 36766 18386 36818 18398
rect 38110 18386 38162 18398
rect 38558 18450 38610 18462
rect 46834 18398 46846 18450
rect 46898 18398 46910 18450
rect 38558 18386 38610 18398
rect 36430 18338 36482 18350
rect 36430 18274 36482 18286
rect 46398 18338 46450 18350
rect 47842 18286 47854 18338
rect 47906 18286 47918 18338
rect 46398 18274 46450 18286
rect 1344 18058 48608 18092
rect 1344 18006 2058 18058
rect 2110 18006 2162 18058
rect 2214 18006 2266 18058
rect 2318 18006 2370 18058
rect 2422 18006 2474 18058
rect 2526 18006 2578 18058
rect 2630 18006 38058 18058
rect 38110 18006 38162 18058
rect 38214 18006 38266 18058
rect 38318 18006 38370 18058
rect 38422 18006 38474 18058
rect 38526 18006 38578 18058
rect 38630 18006 48608 18058
rect 1344 17972 48608 18006
rect 35534 17890 35586 17902
rect 35534 17826 35586 17838
rect 30382 17778 30434 17790
rect 30382 17714 30434 17726
rect 32062 17778 32114 17790
rect 32062 17714 32114 17726
rect 38334 17778 38386 17790
rect 38334 17714 38386 17726
rect 31614 17666 31666 17678
rect 35870 17666 35922 17678
rect 29698 17614 29710 17666
rect 29762 17614 29774 17666
rect 34738 17614 34750 17666
rect 34802 17614 34814 17666
rect 36642 17614 36654 17666
rect 36706 17614 36718 17666
rect 31614 17602 31666 17614
rect 35870 17602 35922 17614
rect 37886 17554 37938 17566
rect 36418 17502 36430 17554
rect 36482 17502 36494 17554
rect 37886 17490 37938 17502
rect 29934 17442 29986 17454
rect 29934 17378 29986 17390
rect 31278 17442 31330 17454
rect 31278 17378 31330 17390
rect 33966 17442 34018 17454
rect 33966 17378 34018 17390
rect 34526 17442 34578 17454
rect 34526 17378 34578 17390
rect 37550 17442 37602 17454
rect 37550 17378 37602 17390
rect 1344 17274 48608 17308
rect 1344 17222 5778 17274
rect 5830 17222 5882 17274
rect 5934 17222 5986 17274
rect 6038 17222 6090 17274
rect 6142 17222 6194 17274
rect 6246 17222 6298 17274
rect 6350 17222 41778 17274
rect 41830 17222 41882 17274
rect 41934 17222 41986 17274
rect 42038 17222 42090 17274
rect 42142 17222 42194 17274
rect 42246 17222 42298 17274
rect 42350 17222 48608 17274
rect 1344 17188 48608 17222
rect 32062 17106 32114 17118
rect 32062 17042 32114 17054
rect 35422 17106 35474 17118
rect 35422 17042 35474 17054
rect 37326 17106 37378 17118
rect 37326 17042 37378 17054
rect 39118 17106 39170 17118
rect 39118 17042 39170 17054
rect 31166 16994 31218 17006
rect 31166 16930 31218 16942
rect 31502 16994 31554 17006
rect 41582 16994 41634 17006
rect 36306 16942 36318 16994
rect 36370 16942 36382 16994
rect 38210 16942 38222 16994
rect 38274 16942 38286 16994
rect 31502 16930 31554 16942
rect 41582 16930 41634 16942
rect 41918 16994 41970 17006
rect 41918 16930 41970 16942
rect 35758 16882 35810 16894
rect 46398 16882 46450 16894
rect 36530 16830 36542 16882
rect 36594 16830 36606 16882
rect 38322 16830 38334 16882
rect 38386 16830 38398 16882
rect 39330 16830 39342 16882
rect 39394 16830 39406 16882
rect 46834 16830 46846 16882
rect 46898 16830 46910 16882
rect 47730 16830 47742 16882
rect 47794 16830 47806 16882
rect 35758 16818 35810 16830
rect 46398 16818 46450 16830
rect 34302 16770 34354 16782
rect 34302 16706 34354 16718
rect 34750 16770 34802 16782
rect 34750 16706 34802 16718
rect 37662 16658 37714 16670
rect 37662 16594 37714 16606
rect 1344 16490 48608 16524
rect 1344 16438 2058 16490
rect 2110 16438 2162 16490
rect 2214 16438 2266 16490
rect 2318 16438 2370 16490
rect 2422 16438 2474 16490
rect 2526 16438 2578 16490
rect 2630 16438 38058 16490
rect 38110 16438 38162 16490
rect 38214 16438 38266 16490
rect 38318 16438 38370 16490
rect 38422 16438 38474 16490
rect 38526 16438 38578 16490
rect 38630 16438 48608 16490
rect 1344 16404 48608 16438
rect 35086 16322 35138 16334
rect 37426 16270 37438 16322
rect 37490 16319 37502 16322
rect 38322 16319 38334 16322
rect 37490 16273 38334 16319
rect 37490 16270 37502 16273
rect 38322 16270 38334 16273
rect 38386 16270 38398 16322
rect 35086 16258 35138 16270
rect 27918 16210 27970 16222
rect 27918 16146 27970 16158
rect 31838 16210 31890 16222
rect 31838 16146 31890 16158
rect 35646 16210 35698 16222
rect 35646 16146 35698 16158
rect 37998 16210 38050 16222
rect 37998 16146 38050 16158
rect 38334 16210 38386 16222
rect 38334 16146 38386 16158
rect 38894 16210 38946 16222
rect 38894 16146 38946 16158
rect 27470 16098 27522 16110
rect 27470 16034 27522 16046
rect 30494 16098 30546 16110
rect 30494 16034 30546 16046
rect 32846 16098 32898 16110
rect 32846 16034 32898 16046
rect 34750 16098 34802 16110
rect 36418 16046 36430 16098
rect 36482 16046 36494 16098
rect 40786 16046 40798 16098
rect 40850 16046 40862 16098
rect 34750 16034 34802 16046
rect 1822 15986 1874 15998
rect 1822 15922 1874 15934
rect 31390 15986 31442 15998
rect 40014 15986 40066 15998
rect 34178 15934 34190 15986
rect 34242 15934 34254 15986
rect 34402 15934 34414 15986
rect 34466 15934 34478 15986
rect 31390 15922 31442 15934
rect 40014 15922 40066 15934
rect 2158 15874 2210 15886
rect 2158 15810 2210 15822
rect 27134 15874 27186 15886
rect 27134 15810 27186 15822
rect 30158 15874 30210 15886
rect 30158 15810 30210 15822
rect 31054 15874 31106 15886
rect 31054 15810 31106 15822
rect 33294 15874 33346 15886
rect 33294 15810 33346 15822
rect 36206 15874 36258 15886
rect 36206 15810 36258 15822
rect 37438 15874 37490 15886
rect 37438 15810 37490 15822
rect 39678 15874 39730 15886
rect 39678 15810 39730 15822
rect 40574 15874 40626 15886
rect 40574 15810 40626 15822
rect 1344 15706 48608 15740
rect 1344 15654 5778 15706
rect 5830 15654 5882 15706
rect 5934 15654 5986 15706
rect 6038 15654 6090 15706
rect 6142 15654 6194 15706
rect 6246 15654 6298 15706
rect 6350 15654 41778 15706
rect 41830 15654 41882 15706
rect 41934 15654 41986 15706
rect 42038 15654 42090 15706
rect 42142 15654 42194 15706
rect 42246 15654 42298 15706
rect 42350 15654 48608 15706
rect 1344 15620 48608 15654
rect 1822 15538 1874 15550
rect 1822 15474 1874 15486
rect 30046 15538 30098 15550
rect 30046 15474 30098 15486
rect 30830 15538 30882 15550
rect 30830 15474 30882 15486
rect 33518 15538 33570 15550
rect 33518 15474 33570 15486
rect 35310 15538 35362 15550
rect 35310 15474 35362 15486
rect 36094 15538 36146 15550
rect 36094 15474 36146 15486
rect 39118 15538 39170 15550
rect 39118 15474 39170 15486
rect 29150 15426 29202 15438
rect 29150 15362 29202 15374
rect 29486 15426 29538 15438
rect 34290 15374 34302 15426
rect 34354 15374 34366 15426
rect 34738 15374 34750 15426
rect 34802 15374 34814 15426
rect 36978 15374 36990 15426
rect 37042 15374 37054 15426
rect 38210 15374 38222 15426
rect 38274 15374 38286 15426
rect 29486 15362 29538 15374
rect 34974 15314 35026 15326
rect 38782 15314 38834 15326
rect 36866 15262 36878 15314
rect 36930 15262 36942 15314
rect 37986 15262 37998 15314
rect 38050 15262 38062 15314
rect 34974 15250 35026 15262
rect 38782 15250 38834 15262
rect 40014 15314 40066 15326
rect 40014 15250 40066 15262
rect 40574 15314 40626 15326
rect 40574 15250 40626 15262
rect 41470 15314 41522 15326
rect 41470 15250 41522 15262
rect 46286 15314 46338 15326
rect 46834 15262 46846 15314
rect 46898 15262 46910 15314
rect 46286 15250 46338 15262
rect 47842 15150 47854 15202
rect 47906 15150 47918 15202
rect 36430 15090 36482 15102
rect 36430 15026 36482 15038
rect 1344 14922 48608 14956
rect 1344 14870 2058 14922
rect 2110 14870 2162 14922
rect 2214 14870 2266 14922
rect 2318 14870 2370 14922
rect 2422 14870 2474 14922
rect 2526 14870 2578 14922
rect 2630 14870 38058 14922
rect 38110 14870 38162 14922
rect 38214 14870 38266 14922
rect 38318 14870 38370 14922
rect 38422 14870 38474 14922
rect 38526 14870 38578 14922
rect 38630 14870 48608 14922
rect 1344 14836 48608 14870
rect 34526 14754 34578 14766
rect 34526 14690 34578 14702
rect 34862 14754 34914 14766
rect 34862 14690 34914 14702
rect 38782 14754 38834 14766
rect 38782 14690 38834 14702
rect 33294 14642 33346 14654
rect 33294 14578 33346 14590
rect 33742 14642 33794 14654
rect 33742 14578 33794 14590
rect 36766 14642 36818 14654
rect 36766 14578 36818 14590
rect 38446 14642 38498 14654
rect 38446 14578 38498 14590
rect 35634 14478 35646 14530
rect 35698 14478 35710 14530
rect 39890 14478 39902 14530
rect 39954 14478 39966 14530
rect 40574 14418 40626 14430
rect 35522 14366 35534 14418
rect 35586 14366 35598 14418
rect 37874 14366 37886 14418
rect 37938 14366 37950 14418
rect 38098 14366 38110 14418
rect 38162 14366 38174 14418
rect 40574 14354 40626 14366
rect 36206 14306 36258 14318
rect 36206 14242 36258 14254
rect 39678 14306 39730 14318
rect 39678 14242 39730 14254
rect 41134 14306 41186 14318
rect 41134 14242 41186 14254
rect 1344 14138 48608 14172
rect 1344 14086 5778 14138
rect 5830 14086 5882 14138
rect 5934 14086 5986 14138
rect 6038 14086 6090 14138
rect 6142 14086 6194 14138
rect 6246 14086 6298 14138
rect 6350 14086 41778 14138
rect 41830 14086 41882 14138
rect 41934 14086 41986 14138
rect 42038 14086 42090 14138
rect 42142 14086 42194 14138
rect 42246 14086 42298 14138
rect 42350 14086 48608 14138
rect 1344 14052 48608 14086
rect 36094 13970 36146 13982
rect 36094 13906 36146 13918
rect 38222 13970 38274 13982
rect 38222 13906 38274 13918
rect 39006 13970 39058 13982
rect 39006 13906 39058 13918
rect 37314 13806 37326 13858
rect 37378 13806 37390 13858
rect 37650 13806 37662 13858
rect 37714 13806 37726 13858
rect 40114 13806 40126 13858
rect 40178 13806 40190 13858
rect 37886 13746 37938 13758
rect 40686 13746 40738 13758
rect 40002 13694 40014 13746
rect 40066 13694 40078 13746
rect 37886 13682 37938 13694
rect 40686 13682 40738 13694
rect 46286 13746 46338 13758
rect 46834 13694 46846 13746
rect 46898 13694 46910 13746
rect 46286 13682 46338 13694
rect 34078 13634 34130 13646
rect 34078 13570 34130 13582
rect 36430 13634 36482 13646
rect 47842 13582 47854 13634
rect 47906 13582 47918 13634
rect 36430 13570 36482 13582
rect 39342 13522 39394 13534
rect 39342 13458 39394 13470
rect 1344 13354 48608 13388
rect 1344 13302 2058 13354
rect 2110 13302 2162 13354
rect 2214 13302 2266 13354
rect 2318 13302 2370 13354
rect 2422 13302 2474 13354
rect 2526 13302 2578 13354
rect 2630 13302 38058 13354
rect 38110 13302 38162 13354
rect 38214 13302 38266 13354
rect 38318 13302 38370 13354
rect 38422 13302 38474 13354
rect 38526 13302 38578 13354
rect 38630 13302 48608 13354
rect 1344 13268 48608 13302
rect 38558 13074 38610 13086
rect 19058 13022 19070 13074
rect 19122 13022 19134 13074
rect 30370 13022 30382 13074
rect 30434 13022 30446 13074
rect 32498 13022 32510 13074
rect 32562 13022 32574 13074
rect 38558 13010 38610 13022
rect 16146 12910 16158 12962
rect 16210 12910 16222 12962
rect 29586 12910 29598 12962
rect 29650 12910 29662 12962
rect 41458 12910 41470 12962
rect 41522 12910 41534 12962
rect 19630 12850 19682 12862
rect 16930 12798 16942 12850
rect 16994 12798 17006 12850
rect 19630 12786 19682 12798
rect 40798 12850 40850 12862
rect 40798 12786 40850 12798
rect 41918 12850 41970 12862
rect 41918 12786 41970 12798
rect 15598 12738 15650 12750
rect 15598 12674 15650 12686
rect 32958 12738 33010 12750
rect 32958 12674 33010 12686
rect 36654 12738 36706 12750
rect 36654 12674 36706 12686
rect 37438 12738 37490 12750
rect 37438 12674 37490 12686
rect 40462 12738 40514 12750
rect 40462 12674 40514 12686
rect 1344 12570 48608 12604
rect 1344 12518 5778 12570
rect 5830 12518 5882 12570
rect 5934 12518 5986 12570
rect 6038 12518 6090 12570
rect 6142 12518 6194 12570
rect 6246 12518 6298 12570
rect 6350 12518 41778 12570
rect 41830 12518 41882 12570
rect 41934 12518 41986 12570
rect 42038 12518 42090 12570
rect 42142 12518 42194 12570
rect 42246 12518 42298 12570
rect 42350 12518 48608 12570
rect 1344 12484 48608 12518
rect 20750 12402 20802 12414
rect 20750 12338 20802 12350
rect 32734 12402 32786 12414
rect 32734 12338 32786 12350
rect 40462 12290 40514 12302
rect 43374 12290 43426 12302
rect 29250 12238 29262 12290
rect 29314 12238 29326 12290
rect 35970 12238 35982 12290
rect 36034 12238 36046 12290
rect 42578 12238 42590 12290
rect 42642 12238 42654 12290
rect 40462 12226 40514 12238
rect 43374 12226 43426 12238
rect 46286 12290 46338 12302
rect 46286 12226 46338 12238
rect 40798 12178 40850 12190
rect 28466 12126 28478 12178
rect 28530 12126 28542 12178
rect 35298 12126 35310 12178
rect 35362 12126 35374 12178
rect 40798 12114 40850 12126
rect 42030 12178 42082 12190
rect 42690 12126 42702 12178
rect 42754 12126 42766 12178
rect 46834 12126 46846 12178
rect 46898 12126 46910 12178
rect 42030 12114 42082 12126
rect 27918 12066 27970 12078
rect 31838 12066 31890 12078
rect 31378 12014 31390 12066
rect 31442 12014 31454 12066
rect 27918 12002 27970 12014
rect 31838 12002 31890 12014
rect 34638 12066 34690 12078
rect 41694 12066 41746 12078
rect 38098 12014 38110 12066
rect 38162 12014 38174 12066
rect 47842 12014 47854 12066
rect 47906 12014 47918 12066
rect 34638 12002 34690 12014
rect 41694 12002 41746 12014
rect 1344 11786 48608 11820
rect 1344 11734 2058 11786
rect 2110 11734 2162 11786
rect 2214 11734 2266 11786
rect 2318 11734 2370 11786
rect 2422 11734 2474 11786
rect 2526 11734 2578 11786
rect 2630 11734 38058 11786
rect 38110 11734 38162 11786
rect 38214 11734 38266 11786
rect 38318 11734 38370 11786
rect 38422 11734 38474 11786
rect 38526 11734 38578 11786
rect 38630 11734 48608 11786
rect 1344 11700 48608 11734
rect 28590 11506 28642 11518
rect 36542 11506 36594 11518
rect 41134 11506 41186 11518
rect 18386 11454 18398 11506
rect 18450 11454 18462 11506
rect 20514 11454 20526 11506
rect 20578 11454 20590 11506
rect 21634 11454 21646 11506
rect 21698 11454 21710 11506
rect 23762 11454 23774 11506
rect 23826 11454 23838 11506
rect 25890 11454 25902 11506
rect 25954 11454 25966 11506
rect 28018 11454 28030 11506
rect 28082 11454 28094 11506
rect 30370 11454 30382 11506
rect 30434 11454 30446 11506
rect 32498 11454 32510 11506
rect 32562 11454 32574 11506
rect 33842 11454 33854 11506
rect 33906 11454 33918 11506
rect 35970 11454 35982 11506
rect 36034 11454 36046 11506
rect 38322 11454 38334 11506
rect 38386 11454 38398 11506
rect 40450 11454 40462 11506
rect 40514 11454 40526 11506
rect 28590 11442 28642 11454
rect 36542 11442 36594 11454
rect 41134 11442 41186 11454
rect 41806 11394 41858 11406
rect 17602 11342 17614 11394
rect 17666 11342 17678 11394
rect 24546 11342 24558 11394
rect 24610 11342 24622 11394
rect 25106 11342 25118 11394
rect 25170 11342 25182 11394
rect 29586 11342 29598 11394
rect 29650 11342 29662 11394
rect 33170 11342 33182 11394
rect 33234 11342 33246 11394
rect 37538 11342 37550 11394
rect 37602 11342 37614 11394
rect 43138 11342 43150 11394
rect 43202 11342 43214 11394
rect 41806 11330 41858 11342
rect 42366 11282 42418 11294
rect 42366 11218 42418 11230
rect 17054 11170 17106 11182
rect 17054 11106 17106 11118
rect 42926 11170 42978 11182
rect 42926 11106 42978 11118
rect 1344 11002 48608 11036
rect 1344 10950 5778 11002
rect 5830 10950 5882 11002
rect 5934 10950 5986 11002
rect 6038 10950 6090 11002
rect 6142 10950 6194 11002
rect 6246 10950 6298 11002
rect 6350 10950 41778 11002
rect 41830 10950 41882 11002
rect 41934 10950 41986 11002
rect 42038 10950 42090 11002
rect 42142 10950 42194 11002
rect 42246 10950 42298 11002
rect 42350 10950 48608 11002
rect 1344 10916 48608 10950
rect 2830 10834 2882 10846
rect 2830 10770 2882 10782
rect 22878 10834 22930 10846
rect 22878 10770 22930 10782
rect 24782 10834 24834 10846
rect 24782 10770 24834 10782
rect 32734 10834 32786 10846
rect 32734 10770 32786 10782
rect 37214 10834 37266 10846
rect 37214 10770 37266 10782
rect 37662 10834 37714 10846
rect 37662 10770 37714 10782
rect 41694 10834 41746 10846
rect 41694 10770 41746 10782
rect 17614 10722 17666 10734
rect 4162 10670 4174 10722
rect 4226 10670 4238 10722
rect 14802 10670 14814 10722
rect 14866 10670 14878 10722
rect 20290 10670 20302 10722
rect 20354 10670 20366 10722
rect 28242 10670 28254 10722
rect 28306 10670 28318 10722
rect 34626 10670 34638 10722
rect 34690 10670 34702 10722
rect 42578 10670 42590 10722
rect 42642 10670 42654 10722
rect 17614 10658 17666 10670
rect 3490 10558 3502 10610
rect 3554 10558 3566 10610
rect 14018 10558 14030 10610
rect 14082 10558 14094 10610
rect 19506 10558 19518 10610
rect 19570 10558 19582 10610
rect 27458 10558 27470 10610
rect 27522 10558 27534 10610
rect 33954 10558 33966 10610
rect 34018 10558 34030 10610
rect 42690 10558 42702 10610
rect 42754 10558 42766 10610
rect 46834 10558 46846 10610
rect 46898 10558 46910 10610
rect 6750 10498 6802 10510
rect 6290 10446 6302 10498
rect 6354 10446 6366 10498
rect 6750 10434 6802 10446
rect 13470 10498 13522 10510
rect 18958 10498 19010 10510
rect 30830 10498 30882 10510
rect 40798 10498 40850 10510
rect 16930 10446 16942 10498
rect 16994 10446 17006 10498
rect 22418 10446 22430 10498
rect 22482 10446 22494 10498
rect 30370 10446 30382 10498
rect 30434 10446 30446 10498
rect 36754 10446 36766 10498
rect 36818 10446 36830 10498
rect 13470 10434 13522 10446
rect 18958 10434 19010 10446
rect 30830 10434 30882 10446
rect 40798 10434 40850 10446
rect 42030 10498 42082 10510
rect 42030 10434 42082 10446
rect 46286 10498 46338 10510
rect 47842 10446 47854 10498
rect 47906 10446 47918 10498
rect 46286 10434 46338 10446
rect 1344 10218 48608 10252
rect 1344 10166 2058 10218
rect 2110 10166 2162 10218
rect 2214 10166 2266 10218
rect 2318 10166 2370 10218
rect 2422 10166 2474 10218
rect 2526 10166 2578 10218
rect 2630 10166 38058 10218
rect 38110 10166 38162 10218
rect 38214 10166 38266 10218
rect 38318 10166 38370 10218
rect 38422 10166 38474 10218
rect 38526 10166 38578 10218
rect 38630 10166 48608 10218
rect 1344 10132 48608 10166
rect 16046 9938 16098 9950
rect 32958 9938 33010 9950
rect 4946 9886 4958 9938
rect 5010 9886 5022 9938
rect 19506 9886 19518 9938
rect 19570 9886 19582 9938
rect 30370 9886 30382 9938
rect 30434 9886 30446 9938
rect 32498 9886 32510 9938
rect 32562 9886 32574 9938
rect 16046 9874 16098 9886
rect 32958 9874 33010 9886
rect 33518 9938 33570 9950
rect 33518 9874 33570 9886
rect 2146 9774 2158 9826
rect 2210 9774 2222 9826
rect 16594 9774 16606 9826
rect 16658 9774 16670 9826
rect 29586 9774 29598 9826
rect 29650 9774 29662 9826
rect 20078 9714 20130 9726
rect 2818 9662 2830 9714
rect 2882 9662 2894 9714
rect 17378 9662 17390 9714
rect 17442 9662 17454 9714
rect 20078 9650 20130 9662
rect 42478 9714 42530 9726
rect 42478 9650 42530 9662
rect 5630 9602 5682 9614
rect 5630 9538 5682 9550
rect 41246 9602 41298 9614
rect 41246 9538 41298 9550
rect 42142 9602 42194 9614
rect 42142 9538 42194 9550
rect 1344 9434 48608 9468
rect 1344 9382 5778 9434
rect 5830 9382 5882 9434
rect 5934 9382 5986 9434
rect 6038 9382 6090 9434
rect 6142 9382 6194 9434
rect 6246 9382 6298 9434
rect 6350 9382 41778 9434
rect 41830 9382 41882 9434
rect 41934 9382 41986 9434
rect 42038 9382 42090 9434
rect 42142 9382 42194 9434
rect 42246 9382 42298 9434
rect 42350 9382 48608 9434
rect 1344 9348 48608 9382
rect 1822 9266 1874 9278
rect 1822 9202 1874 9214
rect 2942 9266 2994 9278
rect 2942 9202 2994 9214
rect 33518 9266 33570 9278
rect 33518 9202 33570 9214
rect 33966 9266 34018 9278
rect 33966 9202 34018 9214
rect 35198 9266 35250 9278
rect 35198 9202 35250 9214
rect 4274 9102 4286 9154
rect 4338 9102 4350 9154
rect 36530 9102 36542 9154
rect 36594 9102 36606 9154
rect 19182 9042 19234 9054
rect 46398 9042 46450 9054
rect 3602 8990 3614 9042
rect 3666 8990 3678 9042
rect 16706 8990 16718 9042
rect 16770 8990 16782 9042
rect 19618 8990 19630 9042
rect 19682 8990 19694 9042
rect 29922 8990 29934 9042
rect 29986 8990 29998 9042
rect 35746 8990 35758 9042
rect 35810 8990 35822 9042
rect 46834 8990 46846 9042
rect 46898 8990 46910 9042
rect 19182 8978 19234 8990
rect 46398 8978 46450 8990
rect 6862 8930 6914 8942
rect 6402 8878 6414 8930
rect 6466 8878 6478 8930
rect 6862 8866 6914 8878
rect 8990 8930 9042 8942
rect 17726 8930 17778 8942
rect 11778 8878 11790 8930
rect 11842 8878 11854 8930
rect 23426 8878 23438 8930
rect 23490 8878 23502 8930
rect 30706 8878 30718 8930
rect 30770 8878 30782 8930
rect 32834 8878 32846 8930
rect 32898 8878 32910 8930
rect 38658 8878 38670 8930
rect 38722 8878 38734 8930
rect 47842 8878 47854 8930
rect 47906 8878 47918 8930
rect 8990 8866 9042 8878
rect 17726 8866 17778 8878
rect 1344 8650 48608 8684
rect 1344 8598 2058 8650
rect 2110 8598 2162 8650
rect 2214 8598 2266 8650
rect 2318 8598 2370 8650
rect 2422 8598 2474 8650
rect 2526 8598 2578 8650
rect 2630 8598 38058 8650
rect 38110 8598 38162 8650
rect 38214 8598 38266 8650
rect 38318 8598 38370 8650
rect 38422 8598 38474 8650
rect 38526 8598 38578 8650
rect 38630 8598 48608 8650
rect 1344 8564 48608 8598
rect 41134 8370 41186 8382
rect 2034 8318 2046 8370
rect 2098 8318 2110 8370
rect 4162 8318 4174 8370
rect 4226 8318 4238 8370
rect 6514 8318 6526 8370
rect 6578 8318 6590 8370
rect 8642 8318 8654 8370
rect 8706 8318 8718 8370
rect 12898 8318 12910 8370
rect 12962 8318 12974 8370
rect 19954 8318 19966 8370
rect 20018 8318 20030 8370
rect 41134 8306 41186 8318
rect 42590 8370 42642 8382
rect 42590 8306 42642 8318
rect 42926 8370 42978 8382
rect 42926 8306 42978 8318
rect 4946 8206 4958 8258
rect 5010 8206 5022 8258
rect 5730 8206 5742 8258
rect 5794 8206 5806 8258
rect 9986 8206 9998 8258
rect 10050 8206 10062 8258
rect 17042 8206 17054 8258
rect 17106 8206 17118 8258
rect 42018 8206 42030 8258
rect 42082 8206 42094 8258
rect 46834 8206 46846 8258
rect 46898 8206 46910 8258
rect 9550 8146 9602 8158
rect 40686 8146 40738 8158
rect 10770 8094 10782 8146
rect 10834 8094 10846 8146
rect 17826 8094 17838 8146
rect 17890 8094 17902 8146
rect 41906 8094 41918 8146
rect 41970 8094 41982 8146
rect 47730 8094 47742 8146
rect 47794 8094 47806 8146
rect 9550 8082 9602 8094
rect 40686 8082 40738 8094
rect 13582 8034 13634 8046
rect 13582 7970 13634 7982
rect 16494 8034 16546 8046
rect 16494 7970 16546 7982
rect 20526 8034 20578 8046
rect 20526 7970 20578 7982
rect 46286 8034 46338 8046
rect 46286 7970 46338 7982
rect 1344 7866 48608 7900
rect 1344 7814 5778 7866
rect 5830 7814 5882 7866
rect 5934 7814 5986 7866
rect 6038 7814 6090 7866
rect 6142 7814 6194 7866
rect 6246 7814 6298 7866
rect 6350 7814 41778 7866
rect 41830 7814 41882 7866
rect 41934 7814 41986 7866
rect 42038 7814 42090 7866
rect 42142 7814 42194 7866
rect 42246 7814 42298 7866
rect 42350 7814 48608 7866
rect 1344 7780 48608 7814
rect 9662 7698 9714 7710
rect 9662 7634 9714 7646
rect 17614 7698 17666 7710
rect 17614 7634 17666 7646
rect 39006 7698 39058 7710
rect 39006 7634 39058 7646
rect 40798 7698 40850 7710
rect 40798 7634 40850 7646
rect 41470 7698 41522 7710
rect 41470 7634 41522 7646
rect 6850 7534 6862 7586
rect 6914 7534 6926 7586
rect 30818 7534 30830 7586
rect 30882 7534 30894 7586
rect 36418 7534 36430 7586
rect 36482 7534 36494 7586
rect 26238 7474 26290 7486
rect 6178 7422 6190 7474
rect 6242 7422 6254 7474
rect 16706 7422 16718 7474
rect 16770 7422 16782 7474
rect 28242 7422 28254 7474
rect 28306 7422 28318 7474
rect 35634 7422 35646 7474
rect 35698 7422 35710 7474
rect 26238 7410 26290 7422
rect 5182 7362 5234 7374
rect 35198 7362 35250 7374
rect 41918 7362 41970 7374
rect 8978 7310 8990 7362
rect 9042 7310 9054 7362
rect 11778 7310 11790 7362
rect 11842 7310 11854 7362
rect 38546 7310 38558 7362
rect 38610 7310 38622 7362
rect 5182 7298 5234 7310
rect 35198 7298 35250 7310
rect 41918 7298 41970 7310
rect 42814 7362 42866 7374
rect 42814 7298 42866 7310
rect 43262 7362 43314 7374
rect 43262 7298 43314 7310
rect 43710 7362 43762 7374
rect 43710 7298 43762 7310
rect 43934 7250 43986 7262
rect 44258 7198 44270 7250
rect 44322 7198 44334 7250
rect 43934 7186 43986 7198
rect 1344 7082 48608 7116
rect 1344 7030 2058 7082
rect 2110 7030 2162 7082
rect 2214 7030 2266 7082
rect 2318 7030 2370 7082
rect 2422 7030 2474 7082
rect 2526 7030 2578 7082
rect 2630 7030 38058 7082
rect 38110 7030 38162 7082
rect 38214 7030 38266 7082
rect 38318 7030 38370 7082
rect 38422 7030 38474 7082
rect 38526 7030 38578 7082
rect 38630 7030 48608 7082
rect 1344 6996 48608 7030
rect 42254 6914 42306 6926
rect 42254 6850 42306 6862
rect 17390 6802 17442 6814
rect 37550 6802 37602 6814
rect 16594 6750 16606 6802
rect 16658 6750 16670 6802
rect 20850 6750 20862 6802
rect 20914 6750 20926 6802
rect 28802 6750 28814 6802
rect 28866 6750 28878 6802
rect 17390 6738 17442 6750
rect 37550 6738 37602 6750
rect 13022 6690 13074 6702
rect 40350 6690 40402 6702
rect 13794 6638 13806 6690
rect 13858 6638 13870 6690
rect 14466 6638 14478 6690
rect 14530 6638 14542 6690
rect 17938 6638 17950 6690
rect 18002 6638 18014 6690
rect 26002 6638 26014 6690
rect 26066 6638 26078 6690
rect 13022 6626 13074 6638
rect 40350 6626 40402 6638
rect 40686 6690 40738 6702
rect 42590 6690 42642 6702
rect 46286 6690 46338 6702
rect 41570 6638 41582 6690
rect 41634 6638 41646 6690
rect 43474 6638 43486 6690
rect 43538 6638 43550 6690
rect 46834 6638 46846 6690
rect 46898 6638 46910 6690
rect 40686 6626 40738 6638
rect 42590 6626 42642 6638
rect 46286 6626 46338 6638
rect 21646 6578 21698 6590
rect 29598 6578 29650 6590
rect 18722 6526 18734 6578
rect 18786 6526 18798 6578
rect 26674 6526 26686 6578
rect 26738 6526 26750 6578
rect 21646 6514 21698 6526
rect 29598 6514 29650 6526
rect 38110 6578 38162 6590
rect 38110 6514 38162 6526
rect 38558 6578 38610 6590
rect 39778 6526 39790 6578
rect 39842 6526 39854 6578
rect 40114 6526 40126 6578
rect 40178 6526 40190 6578
rect 41682 6526 41694 6578
rect 41746 6526 41758 6578
rect 47730 6526 47742 6578
rect 47794 6526 47806 6578
rect 38558 6514 38610 6526
rect 12462 6466 12514 6478
rect 12462 6402 12514 6414
rect 29934 6466 29986 6478
rect 29934 6402 29986 6414
rect 38894 6466 38946 6478
rect 38894 6402 38946 6414
rect 43262 6466 43314 6478
rect 43262 6402 43314 6414
rect 1344 6298 48608 6332
rect 1344 6246 5778 6298
rect 5830 6246 5882 6298
rect 5934 6246 5986 6298
rect 6038 6246 6090 6298
rect 6142 6246 6194 6298
rect 6246 6246 6298 6298
rect 6350 6246 41778 6298
rect 41830 6246 41882 6298
rect 41934 6246 41986 6298
rect 42038 6246 42090 6298
rect 42142 6246 42194 6298
rect 42246 6246 42298 6298
rect 42350 6246 48608 6298
rect 1344 6212 48608 6246
rect 15934 6130 15986 6142
rect 15934 6066 15986 6078
rect 16382 6130 16434 6142
rect 16382 6066 16434 6078
rect 43486 6018 43538 6030
rect 13346 5966 13358 6018
rect 13410 5966 13422 6018
rect 36194 5966 36206 6018
rect 36258 5966 36270 6018
rect 39330 5966 39342 6018
rect 39394 5966 39406 6018
rect 39666 5966 39678 6018
rect 39730 5966 39742 6018
rect 41906 5966 41918 6018
rect 41970 5966 41982 6018
rect 43486 5954 43538 5966
rect 44382 6018 44434 6030
rect 44382 5954 44434 5966
rect 29038 5906 29090 5918
rect 42478 5906 42530 5918
rect 12674 5854 12686 5906
rect 12738 5854 12750 5906
rect 25778 5854 25790 5906
rect 25842 5854 25854 5906
rect 26450 5854 26462 5906
rect 26514 5854 26526 5906
rect 35410 5854 35422 5906
rect 35474 5854 35486 5906
rect 41682 5854 41694 5906
rect 41746 5854 41758 5906
rect 29038 5842 29090 5854
rect 42478 5842 42530 5854
rect 42814 5906 42866 5918
rect 43698 5854 43710 5906
rect 43762 5854 43774 5906
rect 44594 5854 44606 5906
rect 44658 5854 44670 5906
rect 42814 5842 42866 5854
rect 29486 5794 29538 5806
rect 15474 5742 15486 5794
rect 15538 5742 15550 5794
rect 28578 5742 28590 5794
rect 28642 5742 28654 5794
rect 29486 5730 29538 5742
rect 34862 5794 34914 5806
rect 40798 5794 40850 5806
rect 38322 5742 38334 5794
rect 38386 5742 38398 5794
rect 34862 5730 34914 5742
rect 40798 5730 40850 5742
rect 39902 5682 39954 5694
rect 39902 5618 39954 5630
rect 40238 5682 40290 5694
rect 40238 5618 40290 5630
rect 1344 5514 48608 5548
rect 1344 5462 2058 5514
rect 2110 5462 2162 5514
rect 2214 5462 2266 5514
rect 2318 5462 2370 5514
rect 2422 5462 2474 5514
rect 2526 5462 2578 5514
rect 2630 5462 38058 5514
rect 38110 5462 38162 5514
rect 38214 5462 38266 5514
rect 38318 5462 38370 5514
rect 38422 5462 38474 5514
rect 38526 5462 38578 5514
rect 38630 5462 48608 5514
rect 1344 5428 48608 5462
rect 42254 5346 42306 5358
rect 16482 5294 16494 5346
rect 16546 5343 16558 5346
rect 17154 5343 17166 5346
rect 16546 5297 17166 5343
rect 16546 5294 16558 5297
rect 17154 5294 17166 5297
rect 17218 5294 17230 5346
rect 42254 5282 42306 5294
rect 16494 5234 16546 5246
rect 16494 5170 16546 5182
rect 16942 5234 16994 5246
rect 28702 5234 28754 5246
rect 33070 5234 33122 5246
rect 18162 5182 18174 5234
rect 18226 5182 18238 5234
rect 20290 5182 20302 5234
rect 20354 5182 20366 5234
rect 32498 5182 32510 5234
rect 32562 5182 32574 5234
rect 36754 5182 36766 5234
rect 36818 5182 36830 5234
rect 38322 5182 38334 5234
rect 38386 5182 38398 5234
rect 40450 5182 40462 5234
rect 40514 5182 40526 5234
rect 47842 5182 47854 5234
rect 47906 5182 47918 5234
rect 16942 5170 16994 5182
rect 28702 5170 28754 5182
rect 33070 5170 33122 5182
rect 41918 5122 41970 5134
rect 17378 5070 17390 5122
rect 17442 5070 17454 5122
rect 24434 5070 24446 5122
rect 24498 5070 24510 5122
rect 29698 5070 29710 5122
rect 29762 5070 29774 5122
rect 30370 5070 30382 5122
rect 30434 5070 30446 5122
rect 33842 5070 33854 5122
rect 33906 5070 33918 5122
rect 37538 5070 37550 5122
rect 37602 5070 37614 5122
rect 41918 5058 41970 5070
rect 43710 5122 43762 5134
rect 43710 5058 43762 5070
rect 46398 5122 46450 5134
rect 46834 5070 46846 5122
rect 46898 5070 46910 5122
rect 46398 5058 46450 5070
rect 43262 5010 43314 5022
rect 28018 4958 28030 5010
rect 28082 4958 28094 5010
rect 34626 4958 34638 5010
rect 34690 4958 34702 5010
rect 41346 4958 41358 5010
rect 41410 4958 41422 5010
rect 41682 4958 41694 5010
rect 41746 4958 41758 5010
rect 43262 4946 43314 4958
rect 42926 4898 42978 4910
rect 42926 4834 42978 4846
rect 1344 4730 48608 4764
rect 1344 4678 5778 4730
rect 5830 4678 5882 4730
rect 5934 4678 5986 4730
rect 6038 4678 6090 4730
rect 6142 4678 6194 4730
rect 6246 4678 6298 4730
rect 6350 4678 41778 4730
rect 41830 4678 41882 4730
rect 41934 4678 41986 4730
rect 42038 4678 42090 4730
rect 42142 4678 42194 4730
rect 42246 4678 42298 4730
rect 42350 4678 48608 4730
rect 1344 4644 48608 4678
rect 24222 4562 24274 4574
rect 24222 4498 24274 4510
rect 29262 4562 29314 4574
rect 29262 4498 29314 4510
rect 29710 4562 29762 4574
rect 29710 4498 29762 4510
rect 33518 4562 33570 4574
rect 33518 4498 33570 4510
rect 34078 4562 34130 4574
rect 34078 4498 34130 4510
rect 38110 4562 38162 4574
rect 38894 4562 38946 4574
rect 38434 4510 38446 4562
rect 38498 4510 38510 4562
rect 38110 4498 38162 4510
rect 38894 4498 38946 4510
rect 40686 4562 40738 4574
rect 40686 4498 40738 4510
rect 41582 4562 41634 4574
rect 41582 4498 41634 4510
rect 42702 4562 42754 4574
rect 42702 4498 42754 4510
rect 47182 4562 47234 4574
rect 47182 4498 47234 4510
rect 47742 4562 47794 4574
rect 47742 4498 47794 4510
rect 40126 4450 40178 4462
rect 22530 4398 22542 4450
rect 22594 4398 22606 4450
rect 26450 4398 26462 4450
rect 26514 4398 26526 4450
rect 48066 4398 48078 4450
rect 48130 4398 48142 4450
rect 40126 4386 40178 4398
rect 23774 4338 23826 4350
rect 41918 4338 41970 4350
rect 23314 4286 23326 4338
rect 23378 4286 23390 4338
rect 25778 4286 25790 4338
rect 25842 4286 25854 4338
rect 34626 4286 34638 4338
rect 34690 4286 34702 4338
rect 23774 4274 23826 4286
rect 41918 4274 41970 4286
rect 1822 4226 1874 4238
rect 20402 4174 20414 4226
rect 20466 4174 20478 4226
rect 28578 4174 28590 4226
rect 28642 4174 28654 4226
rect 35410 4174 35422 4226
rect 35474 4174 35486 4226
rect 37538 4174 37550 4226
rect 37602 4174 37614 4226
rect 1822 4162 1874 4174
rect 1344 3946 48608 3980
rect 1344 3894 2058 3946
rect 2110 3894 2162 3946
rect 2214 3894 2266 3946
rect 2318 3894 2370 3946
rect 2422 3894 2474 3946
rect 2526 3894 2578 3946
rect 2630 3894 38058 3946
rect 38110 3894 38162 3946
rect 38214 3894 38266 3946
rect 38318 3894 38370 3946
rect 38422 3894 38474 3946
rect 38526 3894 38578 3946
rect 38630 3894 48608 3946
rect 1344 3860 48608 3894
rect 29026 3726 29038 3778
rect 29090 3775 29102 3778
rect 30034 3775 30046 3778
rect 29090 3729 30046 3775
rect 29090 3726 29102 3729
rect 30034 3726 30046 3729
rect 30098 3726 30110 3778
rect 29262 3666 29314 3678
rect 28466 3614 28478 3666
rect 28530 3614 28542 3666
rect 29262 3602 29314 3614
rect 30158 3666 30210 3678
rect 30158 3602 30210 3614
rect 37326 3666 37378 3678
rect 37326 3602 37378 3614
rect 37886 3666 37938 3678
rect 37886 3602 37938 3614
rect 1822 3554 1874 3566
rect 46398 3554 46450 3566
rect 25666 3502 25678 3554
rect 25730 3502 25742 3554
rect 46834 3502 46846 3554
rect 46898 3502 46910 3554
rect 1822 3490 1874 3502
rect 46398 3490 46450 3502
rect 29710 3442 29762 3454
rect 26338 3390 26350 3442
rect 26402 3390 26414 3442
rect 47730 3390 47742 3442
rect 47794 3390 47806 3442
rect 29710 3378 29762 3390
rect 2158 3330 2210 3342
rect 2158 3266 2210 3278
rect 8654 3330 8706 3342
rect 8654 3266 8706 3278
rect 14142 3330 14194 3342
rect 14142 3266 14194 3278
rect 19630 3330 19682 3342
rect 19630 3266 19682 3278
rect 24558 3330 24610 3342
rect 24558 3266 24610 3278
rect 1344 3162 48608 3196
rect 1344 3110 5778 3162
rect 5830 3110 5882 3162
rect 5934 3110 5986 3162
rect 6038 3110 6090 3162
rect 6142 3110 6194 3162
rect 6246 3110 6298 3162
rect 6350 3110 41778 3162
rect 41830 3110 41882 3162
rect 41934 3110 41986 3162
rect 42038 3110 42090 3162
rect 42142 3110 42194 3162
rect 42246 3110 42298 3162
rect 42350 3110 48608 3162
rect 1344 3076 48608 3110
<< via1 >>
rect 2058 46230 2110 46282
rect 2162 46230 2214 46282
rect 2266 46230 2318 46282
rect 2370 46230 2422 46282
rect 2474 46230 2526 46282
rect 2578 46230 2630 46282
rect 38058 46230 38110 46282
rect 38162 46230 38214 46282
rect 38266 46230 38318 46282
rect 38370 46230 38422 46282
rect 38474 46230 38526 46282
rect 38578 46230 38630 46282
rect 1822 46062 1874 46114
rect 46062 45950 46114 46002
rect 45054 45838 45106 45890
rect 46846 45838 46898 45890
rect 47742 45726 47794 45778
rect 44158 45614 44210 45666
rect 5778 45446 5830 45498
rect 5882 45446 5934 45498
rect 5986 45446 6038 45498
rect 6090 45446 6142 45498
rect 6194 45446 6246 45498
rect 6298 45446 6350 45498
rect 41778 45446 41830 45498
rect 41882 45446 41934 45498
rect 41986 45446 42038 45498
rect 42090 45446 42142 45498
rect 42194 45446 42246 45498
rect 42298 45446 42350 45498
rect 45838 45278 45890 45330
rect 46846 45054 46898 45106
rect 46398 44942 46450 44994
rect 47854 44942 47906 44994
rect 2058 44662 2110 44714
rect 2162 44662 2214 44714
rect 2266 44662 2318 44714
rect 2370 44662 2422 44714
rect 2474 44662 2526 44714
rect 2578 44662 2630 44714
rect 38058 44662 38110 44714
rect 38162 44662 38214 44714
rect 38266 44662 38318 44714
rect 38370 44662 38422 44714
rect 38474 44662 38526 44714
rect 38578 44662 38630 44714
rect 46286 44270 46338 44322
rect 46846 44270 46898 44322
rect 47742 44158 47794 44210
rect 5778 43878 5830 43930
rect 5882 43878 5934 43930
rect 5986 43878 6038 43930
rect 6090 43878 6142 43930
rect 6194 43878 6246 43930
rect 6298 43878 6350 43930
rect 41778 43878 41830 43930
rect 41882 43878 41934 43930
rect 41986 43878 42038 43930
rect 42090 43878 42142 43930
rect 42194 43878 42246 43930
rect 42298 43878 42350 43930
rect 2058 43094 2110 43146
rect 2162 43094 2214 43146
rect 2266 43094 2318 43146
rect 2370 43094 2422 43146
rect 2474 43094 2526 43146
rect 2578 43094 2630 43146
rect 38058 43094 38110 43146
rect 38162 43094 38214 43146
rect 38266 43094 38318 43146
rect 38370 43094 38422 43146
rect 38474 43094 38526 43146
rect 38578 43094 38630 43146
rect 46846 42702 46898 42754
rect 47742 42590 47794 42642
rect 46286 42478 46338 42530
rect 5778 42310 5830 42362
rect 5882 42310 5934 42362
rect 5986 42310 6038 42362
rect 6090 42310 6142 42362
rect 6194 42310 6246 42362
rect 6298 42310 6350 42362
rect 41778 42310 41830 42362
rect 41882 42310 41934 42362
rect 41986 42310 42038 42362
rect 42090 42310 42142 42362
rect 42194 42310 42246 42362
rect 42298 42310 42350 42362
rect 2058 41526 2110 41578
rect 2162 41526 2214 41578
rect 2266 41526 2318 41578
rect 2370 41526 2422 41578
rect 2474 41526 2526 41578
rect 2578 41526 2630 41578
rect 38058 41526 38110 41578
rect 38162 41526 38214 41578
rect 38266 41526 38318 41578
rect 38370 41526 38422 41578
rect 38474 41526 38526 41578
rect 38578 41526 38630 41578
rect 3054 41134 3106 41186
rect 46846 41134 46898 41186
rect 2158 41022 2210 41074
rect 47742 41022 47794 41074
rect 3502 40910 3554 40962
rect 46286 40910 46338 40962
rect 5778 40742 5830 40794
rect 5882 40742 5934 40794
rect 5986 40742 6038 40794
rect 6090 40742 6142 40794
rect 6194 40742 6246 40794
rect 6298 40742 6350 40794
rect 41778 40742 41830 40794
rect 41882 40742 41934 40794
rect 41986 40742 42038 40794
rect 42090 40742 42142 40794
rect 42194 40742 42246 40794
rect 42298 40742 42350 40794
rect 2058 39958 2110 40010
rect 2162 39958 2214 40010
rect 2266 39958 2318 40010
rect 2370 39958 2422 40010
rect 2474 39958 2526 40010
rect 2578 39958 2630 40010
rect 38058 39958 38110 40010
rect 38162 39958 38214 40010
rect 38266 39958 38318 40010
rect 38370 39958 38422 40010
rect 38474 39958 38526 40010
rect 38578 39958 38630 40010
rect 46846 39566 46898 39618
rect 47742 39454 47794 39506
rect 46286 39342 46338 39394
rect 5778 39174 5830 39226
rect 5882 39174 5934 39226
rect 5986 39174 6038 39226
rect 6090 39174 6142 39226
rect 6194 39174 6246 39226
rect 6298 39174 6350 39226
rect 41778 39174 41830 39226
rect 41882 39174 41934 39226
rect 41986 39174 42038 39226
rect 42090 39174 42142 39226
rect 42194 39174 42246 39226
rect 42298 39174 42350 39226
rect 46846 38782 46898 38834
rect 46398 38670 46450 38722
rect 47854 38670 47906 38722
rect 2058 38390 2110 38442
rect 2162 38390 2214 38442
rect 2266 38390 2318 38442
rect 2370 38390 2422 38442
rect 2474 38390 2526 38442
rect 2578 38390 2630 38442
rect 38058 38390 38110 38442
rect 38162 38390 38214 38442
rect 38266 38390 38318 38442
rect 38370 38390 38422 38442
rect 38474 38390 38526 38442
rect 38578 38390 38630 38442
rect 5778 37606 5830 37658
rect 5882 37606 5934 37658
rect 5986 37606 6038 37658
rect 6090 37606 6142 37658
rect 6194 37606 6246 37658
rect 6298 37606 6350 37658
rect 41778 37606 41830 37658
rect 41882 37606 41934 37658
rect 41986 37606 42038 37658
rect 42090 37606 42142 37658
rect 42194 37606 42246 37658
rect 42298 37606 42350 37658
rect 46846 37214 46898 37266
rect 46398 37102 46450 37154
rect 47854 37102 47906 37154
rect 2058 36822 2110 36874
rect 2162 36822 2214 36874
rect 2266 36822 2318 36874
rect 2370 36822 2422 36874
rect 2474 36822 2526 36874
rect 2578 36822 2630 36874
rect 38058 36822 38110 36874
rect 38162 36822 38214 36874
rect 38266 36822 38318 36874
rect 38370 36822 38422 36874
rect 38474 36822 38526 36874
rect 38578 36822 38630 36874
rect 17950 36318 18002 36370
rect 18286 36318 18338 36370
rect 17390 36206 17442 36258
rect 5778 36038 5830 36090
rect 5882 36038 5934 36090
rect 5986 36038 6038 36090
rect 6090 36038 6142 36090
rect 6194 36038 6246 36090
rect 6298 36038 6350 36090
rect 41778 36038 41830 36090
rect 41882 36038 41934 36090
rect 41986 36038 42038 36090
rect 42090 36038 42142 36090
rect 42194 36038 42246 36090
rect 42298 36038 42350 36090
rect 46398 35646 46450 35698
rect 46958 35646 47010 35698
rect 47854 35534 47906 35586
rect 2058 35254 2110 35306
rect 2162 35254 2214 35306
rect 2266 35254 2318 35306
rect 2370 35254 2422 35306
rect 2474 35254 2526 35306
rect 2578 35254 2630 35306
rect 38058 35254 38110 35306
rect 38162 35254 38214 35306
rect 38266 35254 38318 35306
rect 38370 35254 38422 35306
rect 38474 35254 38526 35306
rect 38578 35254 38630 35306
rect 1822 34638 1874 34690
rect 5778 34470 5830 34522
rect 5882 34470 5934 34522
rect 5986 34470 6038 34522
rect 6090 34470 6142 34522
rect 6194 34470 6246 34522
rect 6298 34470 6350 34522
rect 41778 34470 41830 34522
rect 41882 34470 41934 34522
rect 41986 34470 42038 34522
rect 42090 34470 42142 34522
rect 42194 34470 42246 34522
rect 42298 34470 42350 34522
rect 46958 34078 47010 34130
rect 46398 33966 46450 34018
rect 46286 33854 46338 33906
rect 46846 33966 46898 34018
rect 47854 33966 47906 34018
rect 2058 33686 2110 33738
rect 2162 33686 2214 33738
rect 2266 33686 2318 33738
rect 2370 33686 2422 33738
rect 2474 33686 2526 33738
rect 2578 33686 2630 33738
rect 38058 33686 38110 33738
rect 38162 33686 38214 33738
rect 38266 33686 38318 33738
rect 38370 33686 38422 33738
rect 38474 33686 38526 33738
rect 38578 33686 38630 33738
rect 5778 32902 5830 32954
rect 5882 32902 5934 32954
rect 5986 32902 6038 32954
rect 6090 32902 6142 32954
rect 6194 32902 6246 32954
rect 6298 32902 6350 32954
rect 41778 32902 41830 32954
rect 41882 32902 41934 32954
rect 41986 32902 42038 32954
rect 42090 32902 42142 32954
rect 42194 32902 42246 32954
rect 42298 32902 42350 32954
rect 46846 32510 46898 32562
rect 46398 32398 46450 32450
rect 47854 32398 47906 32450
rect 2058 32118 2110 32170
rect 2162 32118 2214 32170
rect 2266 32118 2318 32170
rect 2370 32118 2422 32170
rect 2474 32118 2526 32170
rect 2578 32118 2630 32170
rect 38058 32118 38110 32170
rect 38162 32118 38214 32170
rect 38266 32118 38318 32170
rect 38370 32118 38422 32170
rect 38474 32118 38526 32170
rect 38578 32118 38630 32170
rect 5778 31334 5830 31386
rect 5882 31334 5934 31386
rect 5986 31334 6038 31386
rect 6090 31334 6142 31386
rect 6194 31334 6246 31386
rect 6298 31334 6350 31386
rect 41778 31334 41830 31386
rect 41882 31334 41934 31386
rect 41986 31334 42038 31386
rect 42090 31334 42142 31386
rect 42194 31334 42246 31386
rect 42298 31334 42350 31386
rect 46398 30942 46450 30994
rect 46958 30942 47010 30994
rect 46510 30830 46562 30882
rect 46846 30830 46898 30882
rect 47854 30830 47906 30882
rect 2058 30550 2110 30602
rect 2162 30550 2214 30602
rect 2266 30550 2318 30602
rect 2370 30550 2422 30602
rect 2474 30550 2526 30602
rect 2578 30550 2630 30602
rect 38058 30550 38110 30602
rect 38162 30550 38214 30602
rect 38266 30550 38318 30602
rect 38370 30550 38422 30602
rect 38474 30550 38526 30602
rect 38578 30550 38630 30602
rect 5778 29766 5830 29818
rect 5882 29766 5934 29818
rect 5986 29766 6038 29818
rect 6090 29766 6142 29818
rect 6194 29766 6246 29818
rect 6298 29766 6350 29818
rect 41778 29766 41830 29818
rect 41882 29766 41934 29818
rect 41986 29766 42038 29818
rect 42090 29766 42142 29818
rect 42194 29766 42246 29818
rect 42298 29766 42350 29818
rect 39006 29486 39058 29538
rect 38334 29374 38386 29426
rect 38782 29374 38834 29426
rect 46846 29374 46898 29426
rect 36878 29262 36930 29314
rect 37326 29262 37378 29314
rect 39678 29262 39730 29314
rect 46398 29262 46450 29314
rect 47854 29262 47906 29314
rect 37998 29150 38050 29202
rect 2058 28982 2110 29034
rect 2162 28982 2214 29034
rect 2266 28982 2318 29034
rect 2370 28982 2422 29034
rect 2474 28982 2526 29034
rect 2578 28982 2630 29034
rect 38058 28982 38110 29034
rect 38162 28982 38214 29034
rect 38266 28982 38318 29034
rect 38370 28982 38422 29034
rect 38474 28982 38526 29034
rect 38578 28982 38630 29034
rect 39678 28814 39730 28866
rect 40238 28814 40290 28866
rect 36766 28702 36818 28754
rect 38334 28702 38386 28754
rect 47854 28702 47906 28754
rect 37998 28590 38050 28642
rect 46286 28590 46338 28642
rect 46846 28590 46898 28642
rect 1822 28478 1874 28530
rect 38558 28478 38610 28530
rect 38894 28478 38946 28530
rect 40126 28478 40178 28530
rect 2158 28366 2210 28418
rect 39678 28366 39730 28418
rect 5778 28198 5830 28250
rect 5882 28198 5934 28250
rect 5986 28198 6038 28250
rect 6090 28198 6142 28250
rect 6194 28198 6246 28250
rect 6298 28198 6350 28250
rect 41778 28198 41830 28250
rect 41882 28198 41934 28250
rect 41986 28198 42038 28250
rect 42090 28198 42142 28250
rect 42194 28198 42246 28250
rect 42298 28198 42350 28250
rect 1822 28030 1874 28082
rect 36654 28030 36706 28082
rect 38222 27918 38274 27970
rect 37662 27806 37714 27858
rect 38110 27806 38162 27858
rect 39118 27806 39170 27858
rect 39678 27806 39730 27858
rect 36206 27694 36258 27746
rect 37326 27582 37378 27634
rect 2058 27414 2110 27466
rect 2162 27414 2214 27466
rect 2266 27414 2318 27466
rect 2370 27414 2422 27466
rect 2474 27414 2526 27466
rect 2578 27414 2630 27466
rect 38058 27414 38110 27466
rect 38162 27414 38214 27466
rect 38266 27414 38318 27466
rect 38370 27414 38422 27466
rect 38474 27414 38526 27466
rect 38578 27414 38630 27466
rect 38782 27134 38834 27186
rect 46846 27022 46898 27074
rect 39678 26910 39730 26962
rect 46286 26910 46338 26962
rect 47742 26910 47794 26962
rect 40238 26798 40290 26850
rect 5778 26630 5830 26682
rect 5882 26630 5934 26682
rect 5986 26630 6038 26682
rect 6090 26630 6142 26682
rect 6194 26630 6246 26682
rect 6298 26630 6350 26682
rect 41778 26630 41830 26682
rect 41882 26630 41934 26682
rect 41986 26630 42038 26682
rect 42090 26630 42142 26682
rect 42194 26630 42246 26682
rect 42298 26630 42350 26682
rect 39118 26350 39170 26402
rect 39342 26238 39394 26290
rect 37102 26126 37154 26178
rect 37550 26126 37602 26178
rect 38558 26126 38610 26178
rect 38222 26014 38274 26066
rect 2058 25846 2110 25898
rect 2162 25846 2214 25898
rect 2266 25846 2318 25898
rect 2370 25846 2422 25898
rect 2474 25846 2526 25898
rect 2578 25846 2630 25898
rect 38058 25846 38110 25898
rect 38162 25846 38214 25898
rect 38266 25846 38318 25898
rect 38370 25846 38422 25898
rect 38474 25846 38526 25898
rect 38578 25846 38630 25898
rect 40350 25566 40402 25618
rect 46958 25454 47010 25506
rect 47742 25342 47794 25394
rect 40798 25230 40850 25282
rect 46286 25230 46338 25282
rect 5778 25062 5830 25114
rect 5882 25062 5934 25114
rect 5986 25062 6038 25114
rect 6090 25062 6142 25114
rect 6194 25062 6246 25114
rect 6298 25062 6350 25114
rect 41778 25062 41830 25114
rect 41882 25062 41934 25114
rect 41986 25062 42038 25114
rect 42090 25062 42142 25114
rect 42194 25062 42246 25114
rect 42298 25062 42350 25114
rect 39118 24782 39170 24834
rect 38446 24670 38498 24722
rect 39230 24670 39282 24722
rect 36990 24558 37042 24610
rect 37438 24558 37490 24610
rect 38110 24446 38162 24498
rect 2058 24278 2110 24330
rect 2162 24278 2214 24330
rect 2266 24278 2318 24330
rect 2370 24278 2422 24330
rect 2474 24278 2526 24330
rect 2578 24278 2630 24330
rect 38058 24278 38110 24330
rect 38162 24278 38214 24330
rect 38266 24278 38318 24330
rect 38370 24278 38422 24330
rect 38474 24278 38526 24330
rect 38578 24278 38630 24330
rect 39678 23998 39730 24050
rect 38334 23886 38386 23938
rect 39118 23886 39170 23938
rect 40798 23886 40850 23938
rect 46846 23886 46898 23938
rect 39006 23774 39058 23826
rect 40350 23774 40402 23826
rect 47742 23774 47794 23826
rect 36766 23662 36818 23714
rect 37998 23662 38050 23714
rect 46286 23662 46338 23714
rect 5778 23494 5830 23546
rect 5882 23494 5934 23546
rect 5986 23494 6038 23546
rect 6090 23494 6142 23546
rect 6194 23494 6246 23546
rect 6298 23494 6350 23546
rect 41778 23494 41830 23546
rect 41882 23494 41934 23546
rect 41986 23494 42038 23546
rect 42090 23494 42142 23546
rect 42194 23494 42246 23546
rect 42298 23494 42350 23546
rect 39006 23214 39058 23266
rect 39118 23102 39170 23154
rect 36878 22990 36930 23042
rect 37326 22990 37378 23042
rect 37998 22878 38050 22930
rect 38334 22878 38386 22930
rect 2058 22710 2110 22762
rect 2162 22710 2214 22762
rect 2266 22710 2318 22762
rect 2370 22710 2422 22762
rect 2474 22710 2526 22762
rect 2578 22710 2630 22762
rect 38058 22710 38110 22762
rect 38162 22710 38214 22762
rect 38266 22710 38318 22762
rect 38370 22710 38422 22762
rect 38474 22710 38526 22762
rect 38578 22710 38630 22762
rect 46846 22318 46898 22370
rect 28366 22206 28418 22258
rect 38110 22206 38162 22258
rect 38670 22206 38722 22258
rect 47742 22206 47794 22258
rect 1822 22094 1874 22146
rect 28030 22094 28082 22146
rect 38222 22094 38274 22146
rect 46286 22094 46338 22146
rect 5778 21926 5830 21978
rect 5882 21926 5934 21978
rect 5986 21926 6038 21978
rect 6090 21926 6142 21978
rect 6194 21926 6246 21978
rect 6298 21926 6350 21978
rect 41778 21926 41830 21978
rect 41882 21926 41934 21978
rect 41986 21926 42038 21978
rect 42090 21926 42142 21978
rect 42194 21926 42246 21978
rect 42298 21926 42350 21978
rect 38446 21646 38498 21698
rect 38670 21534 38722 21586
rect 36430 21422 36482 21474
rect 36878 21422 36930 21474
rect 37550 21310 37602 21362
rect 37886 21310 37938 21362
rect 2058 21142 2110 21194
rect 2162 21142 2214 21194
rect 2266 21142 2318 21194
rect 2370 21142 2422 21194
rect 2474 21142 2526 21194
rect 2578 21142 2630 21194
rect 38058 21142 38110 21194
rect 38162 21142 38214 21194
rect 38266 21142 38318 21194
rect 38370 21142 38422 21194
rect 38474 21142 38526 21194
rect 38578 21142 38630 21194
rect 29822 20974 29874 21026
rect 37998 20974 38050 21026
rect 31502 20862 31554 20914
rect 36766 20862 36818 20914
rect 30158 20750 30210 20802
rect 30942 20750 30994 20802
rect 38782 20750 38834 20802
rect 46846 20750 46898 20802
rect 30830 20638 30882 20690
rect 33518 20638 33570 20690
rect 38670 20638 38722 20690
rect 39454 20638 39506 20690
rect 39902 20638 39954 20690
rect 40014 20638 40066 20690
rect 40462 20638 40514 20690
rect 40798 20638 40850 20690
rect 47742 20638 47794 20690
rect 28814 20526 28866 20578
rect 33182 20526 33234 20578
rect 36318 20526 36370 20578
rect 37662 20526 37714 20578
rect 39678 20526 39730 20578
rect 46286 20526 46338 20578
rect 5778 20358 5830 20410
rect 5882 20358 5934 20410
rect 5986 20358 6038 20410
rect 6090 20358 6142 20410
rect 6194 20358 6246 20410
rect 6298 20358 6350 20410
rect 41778 20358 41830 20410
rect 41882 20358 41934 20410
rect 41986 20358 42038 20410
rect 42090 20358 42142 20410
rect 42194 20358 42246 20410
rect 42298 20358 42350 20410
rect 33630 20190 33682 20242
rect 29374 20078 29426 20130
rect 32286 20078 32338 20130
rect 34526 20078 34578 20130
rect 37998 20078 38050 20130
rect 32622 19966 32674 20018
rect 33966 19966 34018 20018
rect 34750 19966 34802 20018
rect 37438 19966 37490 20018
rect 38222 19966 38274 20018
rect 35982 19854 36034 19906
rect 36430 19854 36482 19906
rect 39118 19854 39170 19906
rect 37102 19742 37154 19794
rect 2058 19574 2110 19626
rect 2162 19574 2214 19626
rect 2266 19574 2318 19626
rect 2370 19574 2422 19626
rect 2474 19574 2526 19626
rect 2578 19574 2630 19626
rect 38058 19574 38110 19626
rect 38162 19574 38214 19626
rect 38266 19574 38318 19626
rect 38370 19574 38422 19626
rect 38474 19574 38526 19626
rect 38578 19574 38630 19626
rect 34302 19406 34354 19458
rect 37998 19406 38050 19458
rect 36766 19294 36818 19346
rect 38670 19182 38722 19234
rect 46846 19182 46898 19234
rect 31278 19070 31330 19122
rect 34190 19070 34242 19122
rect 37662 19070 37714 19122
rect 38782 19070 38834 19122
rect 47742 19070 47794 19122
rect 30942 18958 30994 19010
rect 33742 18958 33794 19010
rect 34302 18958 34354 19010
rect 34862 18958 34914 19010
rect 35758 18958 35810 19010
rect 36206 18958 36258 19010
rect 46286 18958 46338 19010
rect 5778 18790 5830 18842
rect 5882 18790 5934 18842
rect 5986 18790 6038 18842
rect 6090 18790 6142 18842
rect 6194 18790 6246 18842
rect 6298 18790 6350 18842
rect 41778 18790 41830 18842
rect 41882 18790 41934 18842
rect 41986 18790 42038 18842
rect 42090 18790 42142 18842
rect 42194 18790 42246 18842
rect 42298 18790 42350 18842
rect 30046 18622 30098 18674
rect 29150 18510 29202 18562
rect 29486 18510 29538 18562
rect 30942 18510 30994 18562
rect 31278 18510 31330 18562
rect 31838 18510 31890 18562
rect 32174 18510 32226 18562
rect 35422 18510 35474 18562
rect 37326 18510 37378 18562
rect 34862 18398 34914 18450
rect 35646 18398 35698 18450
rect 36766 18398 36818 18450
rect 37550 18398 37602 18450
rect 38110 18398 38162 18450
rect 38558 18398 38610 18450
rect 46846 18398 46898 18450
rect 36430 18286 36482 18338
rect 46398 18286 46450 18338
rect 47854 18286 47906 18338
rect 2058 18006 2110 18058
rect 2162 18006 2214 18058
rect 2266 18006 2318 18058
rect 2370 18006 2422 18058
rect 2474 18006 2526 18058
rect 2578 18006 2630 18058
rect 38058 18006 38110 18058
rect 38162 18006 38214 18058
rect 38266 18006 38318 18058
rect 38370 18006 38422 18058
rect 38474 18006 38526 18058
rect 38578 18006 38630 18058
rect 35534 17838 35586 17890
rect 30382 17726 30434 17778
rect 32062 17726 32114 17778
rect 38334 17726 38386 17778
rect 29710 17614 29762 17666
rect 31614 17614 31666 17666
rect 34750 17614 34802 17666
rect 35870 17614 35922 17666
rect 36654 17614 36706 17666
rect 36430 17502 36482 17554
rect 37886 17502 37938 17554
rect 29934 17390 29986 17442
rect 31278 17390 31330 17442
rect 33966 17390 34018 17442
rect 34526 17390 34578 17442
rect 37550 17390 37602 17442
rect 5778 17222 5830 17274
rect 5882 17222 5934 17274
rect 5986 17222 6038 17274
rect 6090 17222 6142 17274
rect 6194 17222 6246 17274
rect 6298 17222 6350 17274
rect 41778 17222 41830 17274
rect 41882 17222 41934 17274
rect 41986 17222 42038 17274
rect 42090 17222 42142 17274
rect 42194 17222 42246 17274
rect 42298 17222 42350 17274
rect 32062 17054 32114 17106
rect 35422 17054 35474 17106
rect 37326 17054 37378 17106
rect 39118 17054 39170 17106
rect 31166 16942 31218 16994
rect 31502 16942 31554 16994
rect 36318 16942 36370 16994
rect 38222 16942 38274 16994
rect 41582 16942 41634 16994
rect 41918 16942 41970 16994
rect 35758 16830 35810 16882
rect 36542 16830 36594 16882
rect 38334 16830 38386 16882
rect 39342 16830 39394 16882
rect 46398 16830 46450 16882
rect 46846 16830 46898 16882
rect 47742 16830 47794 16882
rect 34302 16718 34354 16770
rect 34750 16718 34802 16770
rect 37662 16606 37714 16658
rect 2058 16438 2110 16490
rect 2162 16438 2214 16490
rect 2266 16438 2318 16490
rect 2370 16438 2422 16490
rect 2474 16438 2526 16490
rect 2578 16438 2630 16490
rect 38058 16438 38110 16490
rect 38162 16438 38214 16490
rect 38266 16438 38318 16490
rect 38370 16438 38422 16490
rect 38474 16438 38526 16490
rect 38578 16438 38630 16490
rect 35086 16270 35138 16322
rect 37438 16270 37490 16322
rect 38334 16270 38386 16322
rect 27918 16158 27970 16210
rect 31838 16158 31890 16210
rect 35646 16158 35698 16210
rect 37998 16158 38050 16210
rect 38334 16158 38386 16210
rect 38894 16158 38946 16210
rect 27470 16046 27522 16098
rect 30494 16046 30546 16098
rect 32846 16046 32898 16098
rect 34750 16046 34802 16098
rect 36430 16046 36482 16098
rect 40798 16046 40850 16098
rect 1822 15934 1874 15986
rect 31390 15934 31442 15986
rect 34190 15934 34242 15986
rect 34414 15934 34466 15986
rect 40014 15934 40066 15986
rect 2158 15822 2210 15874
rect 27134 15822 27186 15874
rect 30158 15822 30210 15874
rect 31054 15822 31106 15874
rect 33294 15822 33346 15874
rect 36206 15822 36258 15874
rect 37438 15822 37490 15874
rect 39678 15822 39730 15874
rect 40574 15822 40626 15874
rect 5778 15654 5830 15706
rect 5882 15654 5934 15706
rect 5986 15654 6038 15706
rect 6090 15654 6142 15706
rect 6194 15654 6246 15706
rect 6298 15654 6350 15706
rect 41778 15654 41830 15706
rect 41882 15654 41934 15706
rect 41986 15654 42038 15706
rect 42090 15654 42142 15706
rect 42194 15654 42246 15706
rect 42298 15654 42350 15706
rect 1822 15486 1874 15538
rect 30046 15486 30098 15538
rect 30830 15486 30882 15538
rect 33518 15486 33570 15538
rect 35310 15486 35362 15538
rect 36094 15486 36146 15538
rect 39118 15486 39170 15538
rect 29150 15374 29202 15426
rect 29486 15374 29538 15426
rect 34302 15374 34354 15426
rect 34750 15374 34802 15426
rect 36990 15374 37042 15426
rect 38222 15374 38274 15426
rect 34974 15262 35026 15314
rect 36878 15262 36930 15314
rect 37998 15262 38050 15314
rect 38782 15262 38834 15314
rect 40014 15262 40066 15314
rect 40574 15262 40626 15314
rect 41470 15262 41522 15314
rect 46286 15262 46338 15314
rect 46846 15262 46898 15314
rect 47854 15150 47906 15202
rect 36430 15038 36482 15090
rect 2058 14870 2110 14922
rect 2162 14870 2214 14922
rect 2266 14870 2318 14922
rect 2370 14870 2422 14922
rect 2474 14870 2526 14922
rect 2578 14870 2630 14922
rect 38058 14870 38110 14922
rect 38162 14870 38214 14922
rect 38266 14870 38318 14922
rect 38370 14870 38422 14922
rect 38474 14870 38526 14922
rect 38578 14870 38630 14922
rect 34526 14702 34578 14754
rect 34862 14702 34914 14754
rect 38782 14702 38834 14754
rect 33294 14590 33346 14642
rect 33742 14590 33794 14642
rect 36766 14590 36818 14642
rect 38446 14590 38498 14642
rect 35646 14478 35698 14530
rect 39902 14478 39954 14530
rect 35534 14366 35586 14418
rect 37886 14366 37938 14418
rect 38110 14366 38162 14418
rect 40574 14366 40626 14418
rect 36206 14254 36258 14306
rect 39678 14254 39730 14306
rect 41134 14254 41186 14306
rect 5778 14086 5830 14138
rect 5882 14086 5934 14138
rect 5986 14086 6038 14138
rect 6090 14086 6142 14138
rect 6194 14086 6246 14138
rect 6298 14086 6350 14138
rect 41778 14086 41830 14138
rect 41882 14086 41934 14138
rect 41986 14086 42038 14138
rect 42090 14086 42142 14138
rect 42194 14086 42246 14138
rect 42298 14086 42350 14138
rect 36094 13918 36146 13970
rect 38222 13918 38274 13970
rect 39006 13918 39058 13970
rect 37326 13806 37378 13858
rect 37662 13806 37714 13858
rect 40126 13806 40178 13858
rect 37886 13694 37938 13746
rect 40014 13694 40066 13746
rect 40686 13694 40738 13746
rect 46286 13694 46338 13746
rect 46846 13694 46898 13746
rect 34078 13582 34130 13634
rect 36430 13582 36482 13634
rect 47854 13582 47906 13634
rect 39342 13470 39394 13522
rect 2058 13302 2110 13354
rect 2162 13302 2214 13354
rect 2266 13302 2318 13354
rect 2370 13302 2422 13354
rect 2474 13302 2526 13354
rect 2578 13302 2630 13354
rect 38058 13302 38110 13354
rect 38162 13302 38214 13354
rect 38266 13302 38318 13354
rect 38370 13302 38422 13354
rect 38474 13302 38526 13354
rect 38578 13302 38630 13354
rect 19070 13022 19122 13074
rect 30382 13022 30434 13074
rect 32510 13022 32562 13074
rect 38558 13022 38610 13074
rect 16158 12910 16210 12962
rect 29598 12910 29650 12962
rect 41470 12910 41522 12962
rect 16942 12798 16994 12850
rect 19630 12798 19682 12850
rect 40798 12798 40850 12850
rect 41918 12798 41970 12850
rect 15598 12686 15650 12738
rect 32958 12686 33010 12738
rect 36654 12686 36706 12738
rect 37438 12686 37490 12738
rect 40462 12686 40514 12738
rect 5778 12518 5830 12570
rect 5882 12518 5934 12570
rect 5986 12518 6038 12570
rect 6090 12518 6142 12570
rect 6194 12518 6246 12570
rect 6298 12518 6350 12570
rect 41778 12518 41830 12570
rect 41882 12518 41934 12570
rect 41986 12518 42038 12570
rect 42090 12518 42142 12570
rect 42194 12518 42246 12570
rect 42298 12518 42350 12570
rect 20750 12350 20802 12402
rect 32734 12350 32786 12402
rect 29262 12238 29314 12290
rect 35982 12238 36034 12290
rect 40462 12238 40514 12290
rect 42590 12238 42642 12290
rect 43374 12238 43426 12290
rect 46286 12238 46338 12290
rect 28478 12126 28530 12178
rect 35310 12126 35362 12178
rect 40798 12126 40850 12178
rect 42030 12126 42082 12178
rect 42702 12126 42754 12178
rect 46846 12126 46898 12178
rect 27918 12014 27970 12066
rect 31390 12014 31442 12066
rect 31838 12014 31890 12066
rect 34638 12014 34690 12066
rect 38110 12014 38162 12066
rect 41694 12014 41746 12066
rect 47854 12014 47906 12066
rect 2058 11734 2110 11786
rect 2162 11734 2214 11786
rect 2266 11734 2318 11786
rect 2370 11734 2422 11786
rect 2474 11734 2526 11786
rect 2578 11734 2630 11786
rect 38058 11734 38110 11786
rect 38162 11734 38214 11786
rect 38266 11734 38318 11786
rect 38370 11734 38422 11786
rect 38474 11734 38526 11786
rect 38578 11734 38630 11786
rect 18398 11454 18450 11506
rect 20526 11454 20578 11506
rect 21646 11454 21698 11506
rect 23774 11454 23826 11506
rect 25902 11454 25954 11506
rect 28030 11454 28082 11506
rect 28590 11454 28642 11506
rect 30382 11454 30434 11506
rect 32510 11454 32562 11506
rect 33854 11454 33906 11506
rect 35982 11454 36034 11506
rect 36542 11454 36594 11506
rect 38334 11454 38386 11506
rect 40462 11454 40514 11506
rect 41134 11454 41186 11506
rect 17614 11342 17666 11394
rect 24558 11342 24610 11394
rect 25118 11342 25170 11394
rect 29598 11342 29650 11394
rect 33182 11342 33234 11394
rect 37550 11342 37602 11394
rect 41806 11342 41858 11394
rect 43150 11342 43202 11394
rect 42366 11230 42418 11282
rect 17054 11118 17106 11170
rect 42926 11118 42978 11170
rect 5778 10950 5830 11002
rect 5882 10950 5934 11002
rect 5986 10950 6038 11002
rect 6090 10950 6142 11002
rect 6194 10950 6246 11002
rect 6298 10950 6350 11002
rect 41778 10950 41830 11002
rect 41882 10950 41934 11002
rect 41986 10950 42038 11002
rect 42090 10950 42142 11002
rect 42194 10950 42246 11002
rect 42298 10950 42350 11002
rect 2830 10782 2882 10834
rect 22878 10782 22930 10834
rect 24782 10782 24834 10834
rect 32734 10782 32786 10834
rect 37214 10782 37266 10834
rect 37662 10782 37714 10834
rect 41694 10782 41746 10834
rect 4174 10670 4226 10722
rect 14814 10670 14866 10722
rect 17614 10670 17666 10722
rect 20302 10670 20354 10722
rect 28254 10670 28306 10722
rect 34638 10670 34690 10722
rect 42590 10670 42642 10722
rect 3502 10558 3554 10610
rect 14030 10558 14082 10610
rect 19518 10558 19570 10610
rect 27470 10558 27522 10610
rect 33966 10558 34018 10610
rect 42702 10558 42754 10610
rect 46846 10558 46898 10610
rect 6302 10446 6354 10498
rect 6750 10446 6802 10498
rect 13470 10446 13522 10498
rect 16942 10446 16994 10498
rect 18958 10446 19010 10498
rect 22430 10446 22482 10498
rect 30382 10446 30434 10498
rect 30830 10446 30882 10498
rect 36766 10446 36818 10498
rect 40798 10446 40850 10498
rect 42030 10446 42082 10498
rect 46286 10446 46338 10498
rect 47854 10446 47906 10498
rect 2058 10166 2110 10218
rect 2162 10166 2214 10218
rect 2266 10166 2318 10218
rect 2370 10166 2422 10218
rect 2474 10166 2526 10218
rect 2578 10166 2630 10218
rect 38058 10166 38110 10218
rect 38162 10166 38214 10218
rect 38266 10166 38318 10218
rect 38370 10166 38422 10218
rect 38474 10166 38526 10218
rect 38578 10166 38630 10218
rect 4958 9886 5010 9938
rect 16046 9886 16098 9938
rect 19518 9886 19570 9938
rect 30382 9886 30434 9938
rect 32510 9886 32562 9938
rect 32958 9886 33010 9938
rect 33518 9886 33570 9938
rect 2158 9774 2210 9826
rect 16606 9774 16658 9826
rect 29598 9774 29650 9826
rect 2830 9662 2882 9714
rect 17390 9662 17442 9714
rect 20078 9662 20130 9714
rect 42478 9662 42530 9714
rect 5630 9550 5682 9602
rect 41246 9550 41298 9602
rect 42142 9550 42194 9602
rect 5778 9382 5830 9434
rect 5882 9382 5934 9434
rect 5986 9382 6038 9434
rect 6090 9382 6142 9434
rect 6194 9382 6246 9434
rect 6298 9382 6350 9434
rect 41778 9382 41830 9434
rect 41882 9382 41934 9434
rect 41986 9382 42038 9434
rect 42090 9382 42142 9434
rect 42194 9382 42246 9434
rect 42298 9382 42350 9434
rect 1822 9214 1874 9266
rect 2942 9214 2994 9266
rect 33518 9214 33570 9266
rect 33966 9214 34018 9266
rect 35198 9214 35250 9266
rect 4286 9102 4338 9154
rect 36542 9102 36594 9154
rect 3614 8990 3666 9042
rect 16718 8990 16770 9042
rect 19182 8990 19234 9042
rect 19630 8990 19682 9042
rect 29934 8990 29986 9042
rect 35758 8990 35810 9042
rect 46398 8990 46450 9042
rect 46846 8990 46898 9042
rect 6414 8878 6466 8930
rect 6862 8878 6914 8930
rect 8990 8878 9042 8930
rect 11790 8878 11842 8930
rect 17726 8878 17778 8930
rect 23438 8878 23490 8930
rect 30718 8878 30770 8930
rect 32846 8878 32898 8930
rect 38670 8878 38722 8930
rect 47854 8878 47906 8930
rect 2058 8598 2110 8650
rect 2162 8598 2214 8650
rect 2266 8598 2318 8650
rect 2370 8598 2422 8650
rect 2474 8598 2526 8650
rect 2578 8598 2630 8650
rect 38058 8598 38110 8650
rect 38162 8598 38214 8650
rect 38266 8598 38318 8650
rect 38370 8598 38422 8650
rect 38474 8598 38526 8650
rect 38578 8598 38630 8650
rect 2046 8318 2098 8370
rect 4174 8318 4226 8370
rect 6526 8318 6578 8370
rect 8654 8318 8706 8370
rect 12910 8318 12962 8370
rect 19966 8318 20018 8370
rect 41134 8318 41186 8370
rect 42590 8318 42642 8370
rect 42926 8318 42978 8370
rect 4958 8206 5010 8258
rect 5742 8206 5794 8258
rect 9998 8206 10050 8258
rect 17054 8206 17106 8258
rect 42030 8206 42082 8258
rect 46846 8206 46898 8258
rect 9550 8094 9602 8146
rect 10782 8094 10834 8146
rect 17838 8094 17890 8146
rect 40686 8094 40738 8146
rect 41918 8094 41970 8146
rect 47742 8094 47794 8146
rect 13582 7982 13634 8034
rect 16494 7982 16546 8034
rect 20526 7982 20578 8034
rect 46286 7982 46338 8034
rect 5778 7814 5830 7866
rect 5882 7814 5934 7866
rect 5986 7814 6038 7866
rect 6090 7814 6142 7866
rect 6194 7814 6246 7866
rect 6298 7814 6350 7866
rect 41778 7814 41830 7866
rect 41882 7814 41934 7866
rect 41986 7814 42038 7866
rect 42090 7814 42142 7866
rect 42194 7814 42246 7866
rect 42298 7814 42350 7866
rect 9662 7646 9714 7698
rect 17614 7646 17666 7698
rect 39006 7646 39058 7698
rect 40798 7646 40850 7698
rect 41470 7646 41522 7698
rect 6862 7534 6914 7586
rect 30830 7534 30882 7586
rect 36430 7534 36482 7586
rect 6190 7422 6242 7474
rect 16718 7422 16770 7474
rect 26238 7422 26290 7474
rect 28254 7422 28306 7474
rect 35646 7422 35698 7474
rect 5182 7310 5234 7362
rect 8990 7310 9042 7362
rect 11790 7310 11842 7362
rect 35198 7310 35250 7362
rect 38558 7310 38610 7362
rect 41918 7310 41970 7362
rect 42814 7310 42866 7362
rect 43262 7310 43314 7362
rect 43710 7310 43762 7362
rect 43934 7198 43986 7250
rect 44270 7198 44322 7250
rect 2058 7030 2110 7082
rect 2162 7030 2214 7082
rect 2266 7030 2318 7082
rect 2370 7030 2422 7082
rect 2474 7030 2526 7082
rect 2578 7030 2630 7082
rect 38058 7030 38110 7082
rect 38162 7030 38214 7082
rect 38266 7030 38318 7082
rect 38370 7030 38422 7082
rect 38474 7030 38526 7082
rect 38578 7030 38630 7082
rect 42254 6862 42306 6914
rect 16606 6750 16658 6802
rect 17390 6750 17442 6802
rect 20862 6750 20914 6802
rect 28814 6750 28866 6802
rect 37550 6750 37602 6802
rect 13022 6638 13074 6690
rect 13806 6638 13858 6690
rect 14478 6638 14530 6690
rect 17950 6638 18002 6690
rect 26014 6638 26066 6690
rect 40350 6638 40402 6690
rect 40686 6638 40738 6690
rect 41582 6638 41634 6690
rect 42590 6638 42642 6690
rect 43486 6638 43538 6690
rect 46286 6638 46338 6690
rect 46846 6638 46898 6690
rect 18734 6526 18786 6578
rect 21646 6526 21698 6578
rect 26686 6526 26738 6578
rect 29598 6526 29650 6578
rect 38110 6526 38162 6578
rect 38558 6526 38610 6578
rect 39790 6526 39842 6578
rect 40126 6526 40178 6578
rect 41694 6526 41746 6578
rect 47742 6526 47794 6578
rect 12462 6414 12514 6466
rect 29934 6414 29986 6466
rect 38894 6414 38946 6466
rect 43262 6414 43314 6466
rect 5778 6246 5830 6298
rect 5882 6246 5934 6298
rect 5986 6246 6038 6298
rect 6090 6246 6142 6298
rect 6194 6246 6246 6298
rect 6298 6246 6350 6298
rect 41778 6246 41830 6298
rect 41882 6246 41934 6298
rect 41986 6246 42038 6298
rect 42090 6246 42142 6298
rect 42194 6246 42246 6298
rect 42298 6246 42350 6298
rect 15934 6078 15986 6130
rect 16382 6078 16434 6130
rect 13358 5966 13410 6018
rect 36206 5966 36258 6018
rect 39342 5966 39394 6018
rect 39678 5966 39730 6018
rect 41918 5966 41970 6018
rect 43486 5966 43538 6018
rect 44382 5966 44434 6018
rect 12686 5854 12738 5906
rect 25790 5854 25842 5906
rect 26462 5854 26514 5906
rect 29038 5854 29090 5906
rect 35422 5854 35474 5906
rect 41694 5854 41746 5906
rect 42478 5854 42530 5906
rect 42814 5854 42866 5906
rect 43710 5854 43762 5906
rect 44606 5854 44658 5906
rect 15486 5742 15538 5794
rect 28590 5742 28642 5794
rect 29486 5742 29538 5794
rect 34862 5742 34914 5794
rect 38334 5742 38386 5794
rect 40798 5742 40850 5794
rect 39902 5630 39954 5682
rect 40238 5630 40290 5682
rect 2058 5462 2110 5514
rect 2162 5462 2214 5514
rect 2266 5462 2318 5514
rect 2370 5462 2422 5514
rect 2474 5462 2526 5514
rect 2578 5462 2630 5514
rect 38058 5462 38110 5514
rect 38162 5462 38214 5514
rect 38266 5462 38318 5514
rect 38370 5462 38422 5514
rect 38474 5462 38526 5514
rect 38578 5462 38630 5514
rect 16494 5294 16546 5346
rect 17166 5294 17218 5346
rect 42254 5294 42306 5346
rect 16494 5182 16546 5234
rect 16942 5182 16994 5234
rect 18174 5182 18226 5234
rect 20302 5182 20354 5234
rect 28702 5182 28754 5234
rect 32510 5182 32562 5234
rect 33070 5182 33122 5234
rect 36766 5182 36818 5234
rect 38334 5182 38386 5234
rect 40462 5182 40514 5234
rect 47854 5182 47906 5234
rect 17390 5070 17442 5122
rect 24446 5070 24498 5122
rect 29710 5070 29762 5122
rect 30382 5070 30434 5122
rect 33854 5070 33906 5122
rect 37550 5070 37602 5122
rect 41918 5070 41970 5122
rect 43710 5070 43762 5122
rect 46398 5070 46450 5122
rect 46846 5070 46898 5122
rect 28030 4958 28082 5010
rect 34638 4958 34690 5010
rect 41358 4958 41410 5010
rect 41694 4958 41746 5010
rect 43262 4958 43314 5010
rect 42926 4846 42978 4898
rect 5778 4678 5830 4730
rect 5882 4678 5934 4730
rect 5986 4678 6038 4730
rect 6090 4678 6142 4730
rect 6194 4678 6246 4730
rect 6298 4678 6350 4730
rect 41778 4678 41830 4730
rect 41882 4678 41934 4730
rect 41986 4678 42038 4730
rect 42090 4678 42142 4730
rect 42194 4678 42246 4730
rect 42298 4678 42350 4730
rect 24222 4510 24274 4562
rect 29262 4510 29314 4562
rect 29710 4510 29762 4562
rect 33518 4510 33570 4562
rect 34078 4510 34130 4562
rect 38110 4510 38162 4562
rect 38446 4510 38498 4562
rect 38894 4510 38946 4562
rect 40686 4510 40738 4562
rect 41582 4510 41634 4562
rect 42702 4510 42754 4562
rect 47182 4510 47234 4562
rect 47742 4510 47794 4562
rect 22542 4398 22594 4450
rect 26462 4398 26514 4450
rect 40126 4398 40178 4450
rect 48078 4398 48130 4450
rect 23326 4286 23378 4338
rect 23774 4286 23826 4338
rect 25790 4286 25842 4338
rect 34638 4286 34690 4338
rect 41918 4286 41970 4338
rect 1822 4174 1874 4226
rect 20414 4174 20466 4226
rect 28590 4174 28642 4226
rect 35422 4174 35474 4226
rect 37550 4174 37602 4226
rect 2058 3894 2110 3946
rect 2162 3894 2214 3946
rect 2266 3894 2318 3946
rect 2370 3894 2422 3946
rect 2474 3894 2526 3946
rect 2578 3894 2630 3946
rect 38058 3894 38110 3946
rect 38162 3894 38214 3946
rect 38266 3894 38318 3946
rect 38370 3894 38422 3946
rect 38474 3894 38526 3946
rect 38578 3894 38630 3946
rect 29038 3726 29090 3778
rect 30046 3726 30098 3778
rect 28478 3614 28530 3666
rect 29262 3614 29314 3666
rect 30158 3614 30210 3666
rect 37326 3614 37378 3666
rect 37886 3614 37938 3666
rect 1822 3502 1874 3554
rect 25678 3502 25730 3554
rect 46398 3502 46450 3554
rect 46846 3502 46898 3554
rect 26350 3390 26402 3442
rect 29710 3390 29762 3442
rect 47742 3390 47794 3442
rect 2158 3278 2210 3330
rect 8654 3278 8706 3330
rect 14142 3278 14194 3330
rect 19630 3278 19682 3330
rect 24558 3278 24610 3330
rect 5778 3110 5830 3162
rect 5882 3110 5934 3162
rect 5986 3110 6038 3162
rect 6090 3110 6142 3162
rect 6194 3110 6246 3162
rect 6298 3110 6350 3162
rect 41778 3110 41830 3162
rect 41882 3110 41934 3162
rect 41986 3110 42038 3162
rect 42090 3110 42142 3162
rect 42194 3110 42246 3162
rect 42298 3110 42350 3162
<< metal2 >>
rect 46060 48244 46116 48254
rect 1820 46452 1876 46462
rect 1820 46114 1876 46396
rect 2056 46284 2632 46294
rect 2112 46228 2160 46284
rect 2216 46228 2264 46284
rect 2320 46228 2368 46284
rect 2424 46228 2472 46284
rect 2528 46228 2576 46284
rect 2056 46218 2632 46228
rect 38056 46284 38632 46294
rect 38112 46228 38160 46284
rect 38216 46228 38264 46284
rect 38320 46228 38368 46284
rect 38424 46228 38472 46284
rect 38528 46228 38576 46284
rect 38056 46218 38632 46228
rect 1820 46062 1822 46114
rect 1874 46062 1876 46114
rect 1820 46050 1876 46062
rect 46060 46002 46116 48188
rect 46060 45950 46062 46002
rect 46114 45950 46116 46002
rect 46060 45938 46116 45950
rect 47852 46788 47908 46798
rect 45052 45890 45108 45902
rect 46844 45892 46900 45902
rect 45052 45838 45054 45890
rect 45106 45838 45108 45890
rect 44156 45668 44212 45678
rect 45052 45668 45108 45838
rect 44156 45666 45108 45668
rect 44156 45614 44158 45666
rect 44210 45614 45108 45666
rect 44156 45612 45108 45614
rect 46172 45890 46900 45892
rect 46172 45838 46846 45890
rect 46898 45838 46900 45890
rect 46172 45836 46900 45838
rect 5776 45500 6352 45510
rect 5832 45444 5880 45500
rect 5936 45444 5984 45500
rect 6040 45444 6088 45500
rect 6144 45444 6192 45500
rect 6248 45444 6296 45500
rect 5776 45434 6352 45444
rect 41776 45500 42352 45510
rect 41832 45444 41880 45500
rect 41936 45444 41984 45500
rect 42040 45444 42088 45500
rect 42144 45444 42192 45500
rect 42248 45444 42296 45500
rect 41776 45434 42352 45444
rect 2056 44716 2632 44726
rect 2112 44660 2160 44716
rect 2216 44660 2264 44716
rect 2320 44660 2368 44716
rect 2424 44660 2472 44716
rect 2528 44660 2576 44716
rect 2056 44650 2632 44660
rect 38056 44716 38632 44726
rect 38112 44660 38160 44716
rect 38216 44660 38264 44716
rect 38320 44660 38368 44716
rect 38424 44660 38472 44716
rect 38528 44660 38576 44716
rect 38056 44650 38632 44660
rect 5776 43932 6352 43942
rect 5832 43876 5880 43932
rect 5936 43876 5984 43932
rect 6040 43876 6088 43932
rect 6144 43876 6192 43932
rect 6248 43876 6296 43932
rect 5776 43866 6352 43876
rect 41776 43932 42352 43942
rect 41832 43876 41880 43932
rect 41936 43876 41984 43932
rect 42040 43876 42088 43932
rect 42144 43876 42192 43932
rect 42248 43876 42296 43932
rect 41776 43866 42352 43876
rect 2056 43148 2632 43158
rect 2112 43092 2160 43148
rect 2216 43092 2264 43148
rect 2320 43092 2368 43148
rect 2424 43092 2472 43148
rect 2528 43092 2576 43148
rect 2056 43082 2632 43092
rect 38056 43148 38632 43158
rect 38112 43092 38160 43148
rect 38216 43092 38264 43148
rect 38320 43092 38368 43148
rect 38424 43092 38472 43148
rect 38528 43092 38576 43148
rect 38056 43082 38632 43092
rect 5776 42364 6352 42374
rect 5832 42308 5880 42364
rect 5936 42308 5984 42364
rect 6040 42308 6088 42364
rect 6144 42308 6192 42364
rect 6248 42308 6296 42364
rect 5776 42298 6352 42308
rect 41776 42364 42352 42374
rect 41832 42308 41880 42364
rect 41936 42308 41984 42364
rect 42040 42308 42088 42364
rect 42144 42308 42192 42364
rect 42248 42308 42296 42364
rect 41776 42298 42352 42308
rect 40236 41972 40292 41982
rect 2056 41580 2632 41590
rect 2112 41524 2160 41580
rect 2216 41524 2264 41580
rect 2320 41524 2368 41580
rect 2424 41524 2472 41580
rect 2528 41524 2576 41580
rect 2056 41514 2632 41524
rect 38056 41580 38632 41590
rect 38112 41524 38160 41580
rect 38216 41524 38264 41580
rect 38320 41524 38368 41580
rect 38424 41524 38472 41580
rect 38528 41524 38576 41580
rect 38056 41514 38632 41524
rect 3052 41186 3108 41198
rect 3052 41134 3054 41186
rect 3106 41134 3108 41186
rect 2156 41074 2212 41086
rect 2156 41022 2158 41074
rect 2210 41022 2212 41074
rect 2156 40516 2212 41022
rect 3052 40964 3108 41134
rect 3052 40898 3108 40908
rect 3500 40964 3556 40974
rect 3500 40870 3556 40908
rect 17948 40964 18004 40974
rect 5776 40796 6352 40806
rect 5832 40740 5880 40796
rect 5936 40740 5984 40796
rect 6040 40740 6088 40796
rect 6144 40740 6192 40796
rect 6248 40740 6296 40796
rect 5776 40730 6352 40740
rect 2156 40450 2212 40460
rect 2056 40012 2632 40022
rect 2112 39956 2160 40012
rect 2216 39956 2264 40012
rect 2320 39956 2368 40012
rect 2424 39956 2472 40012
rect 2528 39956 2576 40012
rect 2056 39946 2632 39956
rect 5776 39228 6352 39238
rect 5832 39172 5880 39228
rect 5936 39172 5984 39228
rect 6040 39172 6088 39228
rect 6144 39172 6192 39228
rect 6248 39172 6296 39228
rect 5776 39162 6352 39172
rect 2056 38444 2632 38454
rect 2112 38388 2160 38444
rect 2216 38388 2264 38444
rect 2320 38388 2368 38444
rect 2424 38388 2472 38444
rect 2528 38388 2576 38444
rect 2056 38378 2632 38388
rect 5776 37660 6352 37670
rect 5832 37604 5880 37660
rect 5936 37604 5984 37660
rect 6040 37604 6088 37660
rect 6144 37604 6192 37660
rect 6248 37604 6296 37660
rect 5776 37594 6352 37604
rect 2056 36876 2632 36886
rect 2112 36820 2160 36876
rect 2216 36820 2264 36876
rect 2320 36820 2368 36876
rect 2424 36820 2472 36876
rect 2528 36820 2576 36876
rect 2056 36810 2632 36820
rect 17388 36372 17444 36382
rect 17388 36258 17444 36316
rect 17948 36370 18004 40908
rect 38056 40012 38632 40022
rect 38112 39956 38160 40012
rect 38216 39956 38264 40012
rect 38320 39956 38368 40012
rect 38424 39956 38472 40012
rect 38528 39956 38576 40012
rect 38056 39946 38632 39956
rect 38056 38444 38632 38454
rect 38112 38388 38160 38444
rect 38216 38388 38264 38444
rect 38320 38388 38368 38444
rect 38424 38388 38472 38444
rect 38528 38388 38576 38444
rect 38056 38378 38632 38388
rect 38056 36876 38632 36886
rect 38112 36820 38160 36876
rect 38216 36820 38264 36876
rect 38320 36820 38368 36876
rect 38424 36820 38472 36876
rect 38528 36820 38576 36876
rect 38056 36810 38632 36820
rect 17948 36318 17950 36370
rect 18002 36318 18004 36370
rect 17948 36306 18004 36318
rect 18284 36372 18340 36382
rect 18284 36278 18340 36316
rect 17388 36206 17390 36258
rect 17442 36206 17444 36258
rect 5776 36092 6352 36102
rect 5832 36036 5880 36092
rect 5936 36036 5984 36092
rect 6040 36036 6088 36092
rect 6144 36036 6192 36092
rect 6248 36036 6296 36092
rect 5776 36026 6352 36036
rect 2056 35308 2632 35318
rect 2112 35252 2160 35308
rect 2216 35252 2264 35308
rect 2320 35252 2368 35308
rect 2424 35252 2472 35308
rect 2528 35252 2576 35308
rect 2056 35242 2632 35252
rect 1820 34690 1876 34702
rect 1820 34638 1822 34690
rect 1874 34638 1876 34690
rect 1820 34356 1876 34638
rect 5776 34524 6352 34534
rect 5832 34468 5880 34524
rect 5936 34468 5984 34524
rect 6040 34468 6088 34524
rect 6144 34468 6192 34524
rect 6248 34468 6296 34524
rect 5776 34458 6352 34468
rect 1820 34290 1876 34300
rect 2056 33740 2632 33750
rect 2112 33684 2160 33740
rect 2216 33684 2264 33740
rect 2320 33684 2368 33740
rect 2424 33684 2472 33740
rect 2528 33684 2576 33740
rect 2056 33674 2632 33684
rect 5776 32956 6352 32966
rect 5832 32900 5880 32956
rect 5936 32900 5984 32956
rect 6040 32900 6088 32956
rect 6144 32900 6192 32956
rect 6248 32900 6296 32956
rect 5776 32890 6352 32900
rect 2056 32172 2632 32182
rect 2112 32116 2160 32172
rect 2216 32116 2264 32172
rect 2320 32116 2368 32172
rect 2424 32116 2472 32172
rect 2528 32116 2576 32172
rect 2056 32106 2632 32116
rect 5776 31388 6352 31398
rect 5832 31332 5880 31388
rect 5936 31332 5984 31388
rect 6040 31332 6088 31388
rect 6144 31332 6192 31388
rect 6248 31332 6296 31388
rect 5776 31322 6352 31332
rect 2056 30604 2632 30614
rect 2112 30548 2160 30604
rect 2216 30548 2264 30604
rect 2320 30548 2368 30604
rect 2424 30548 2472 30604
rect 2528 30548 2576 30604
rect 2056 30538 2632 30548
rect 5776 29820 6352 29830
rect 5832 29764 5880 29820
rect 5936 29764 5984 29820
rect 6040 29764 6088 29820
rect 6144 29764 6192 29820
rect 6248 29764 6296 29820
rect 5776 29754 6352 29764
rect 2056 29036 2632 29046
rect 2112 28980 2160 29036
rect 2216 28980 2264 29036
rect 2320 28980 2368 29036
rect 2424 28980 2472 29036
rect 2528 28980 2576 29036
rect 2056 28970 2632 28980
rect 1820 28530 1876 28542
rect 1820 28478 1822 28530
rect 1874 28478 1876 28530
rect 1820 28084 1876 28478
rect 2156 28420 2212 28430
rect 2156 28418 2884 28420
rect 2156 28366 2158 28418
rect 2210 28366 2884 28418
rect 2156 28364 2884 28366
rect 2156 28354 2212 28364
rect 1820 27990 1876 28028
rect 2056 27468 2632 27478
rect 2112 27412 2160 27468
rect 2216 27412 2264 27468
rect 2320 27412 2368 27468
rect 2424 27412 2472 27468
rect 2528 27412 2576 27468
rect 2056 27402 2632 27412
rect 2056 25900 2632 25910
rect 2112 25844 2160 25900
rect 2216 25844 2264 25900
rect 2320 25844 2368 25900
rect 2424 25844 2472 25900
rect 2528 25844 2576 25900
rect 2056 25834 2632 25844
rect 2056 24332 2632 24342
rect 2112 24276 2160 24332
rect 2216 24276 2264 24332
rect 2320 24276 2368 24332
rect 2424 24276 2472 24332
rect 2528 24276 2576 24332
rect 2056 24266 2632 24276
rect 2056 22764 2632 22774
rect 2112 22708 2160 22764
rect 2216 22708 2264 22764
rect 2320 22708 2368 22764
rect 2424 22708 2472 22764
rect 2528 22708 2576 22764
rect 2056 22698 2632 22708
rect 1820 22146 1876 22158
rect 1820 22094 1822 22146
rect 1874 22094 1876 22146
rect 1820 22036 1876 22094
rect 1820 21970 1876 21980
rect 2056 21196 2632 21206
rect 2112 21140 2160 21196
rect 2216 21140 2264 21196
rect 2320 21140 2368 21196
rect 2424 21140 2472 21196
rect 2528 21140 2576 21196
rect 2056 21130 2632 21140
rect 2056 19628 2632 19638
rect 2112 19572 2160 19628
rect 2216 19572 2264 19628
rect 2320 19572 2368 19628
rect 2424 19572 2472 19628
rect 2528 19572 2576 19628
rect 2056 19562 2632 19572
rect 2056 18060 2632 18070
rect 2112 18004 2160 18060
rect 2216 18004 2264 18060
rect 2320 18004 2368 18060
rect 2424 18004 2472 18060
rect 2528 18004 2576 18060
rect 2056 17994 2632 18004
rect 2056 16492 2632 16502
rect 2112 16436 2160 16492
rect 2216 16436 2264 16492
rect 2320 16436 2368 16492
rect 2424 16436 2472 16492
rect 2528 16436 2576 16492
rect 2056 16426 2632 16436
rect 1820 15986 1876 15998
rect 1820 15934 1822 15986
rect 1874 15934 1876 15986
rect 1820 15652 1876 15934
rect 2156 15876 2212 15886
rect 2156 15874 2772 15876
rect 2156 15822 2158 15874
rect 2210 15822 2772 15874
rect 2156 15820 2772 15822
rect 2156 15810 2212 15820
rect 1820 15538 1876 15596
rect 1820 15486 1822 15538
rect 1874 15486 1876 15538
rect 1820 15474 1876 15486
rect 2056 14924 2632 14934
rect 2112 14868 2160 14924
rect 2216 14868 2264 14924
rect 2320 14868 2368 14924
rect 2424 14868 2472 14924
rect 2528 14868 2576 14924
rect 2056 14858 2632 14868
rect 2056 13356 2632 13366
rect 2112 13300 2160 13356
rect 2216 13300 2264 13356
rect 2320 13300 2368 13356
rect 2424 13300 2472 13356
rect 2528 13300 2576 13356
rect 2056 13290 2632 13300
rect 2056 11788 2632 11798
rect 2112 11732 2160 11788
rect 2216 11732 2264 11788
rect 2320 11732 2368 11788
rect 2424 11732 2472 11788
rect 2528 11732 2576 11788
rect 2056 11722 2632 11732
rect 2716 10500 2772 15820
rect 2828 10834 2884 28364
rect 5776 28252 6352 28262
rect 5832 28196 5880 28252
rect 5936 28196 5984 28252
rect 6040 28196 6088 28252
rect 6144 28196 6192 28252
rect 6248 28196 6296 28252
rect 5776 28186 6352 28196
rect 5776 26684 6352 26694
rect 5832 26628 5880 26684
rect 5936 26628 5984 26684
rect 6040 26628 6088 26684
rect 6144 26628 6192 26684
rect 6248 26628 6296 26684
rect 5776 26618 6352 26628
rect 5776 25116 6352 25126
rect 5832 25060 5880 25116
rect 5936 25060 5984 25116
rect 6040 25060 6088 25116
rect 6144 25060 6192 25116
rect 6248 25060 6296 25116
rect 5776 25050 6352 25060
rect 5776 23548 6352 23558
rect 5832 23492 5880 23548
rect 5936 23492 5984 23548
rect 6040 23492 6088 23548
rect 6144 23492 6192 23548
rect 6248 23492 6296 23548
rect 5776 23482 6352 23492
rect 12908 22260 12964 22270
rect 5776 21980 6352 21990
rect 5832 21924 5880 21980
rect 5936 21924 5984 21980
rect 6040 21924 6088 21980
rect 6144 21924 6192 21980
rect 6248 21924 6296 21980
rect 5776 21914 6352 21924
rect 5776 20412 6352 20422
rect 5832 20356 5880 20412
rect 5936 20356 5984 20412
rect 6040 20356 6088 20412
rect 6144 20356 6192 20412
rect 6248 20356 6296 20412
rect 5776 20346 6352 20356
rect 5776 18844 6352 18854
rect 5832 18788 5880 18844
rect 5936 18788 5984 18844
rect 6040 18788 6088 18844
rect 6144 18788 6192 18844
rect 6248 18788 6296 18844
rect 5776 18778 6352 18788
rect 5776 17276 6352 17286
rect 5832 17220 5880 17276
rect 5936 17220 5984 17276
rect 6040 17220 6088 17276
rect 6144 17220 6192 17276
rect 6248 17220 6296 17276
rect 5776 17210 6352 17220
rect 5776 15708 6352 15718
rect 5832 15652 5880 15708
rect 5936 15652 5984 15708
rect 6040 15652 6088 15708
rect 6144 15652 6192 15708
rect 6248 15652 6296 15708
rect 5776 15642 6352 15652
rect 5776 14140 6352 14150
rect 5832 14084 5880 14140
rect 5936 14084 5984 14140
rect 6040 14084 6088 14140
rect 6144 14084 6192 14140
rect 6248 14084 6296 14140
rect 5776 14074 6352 14084
rect 5776 12572 6352 12582
rect 5832 12516 5880 12572
rect 5936 12516 5984 12572
rect 6040 12516 6088 12572
rect 6144 12516 6192 12572
rect 6248 12516 6296 12572
rect 5776 12506 6352 12516
rect 5776 11004 6352 11014
rect 5832 10948 5880 11004
rect 5936 10948 5984 11004
rect 6040 10948 6088 11004
rect 6144 10948 6192 11004
rect 6248 10948 6296 11004
rect 5776 10938 6352 10948
rect 2828 10782 2830 10834
rect 2882 10782 2884 10834
rect 2828 10724 2884 10782
rect 2828 10658 2884 10668
rect 4172 10724 4228 10734
rect 4172 10630 4228 10668
rect 3500 10612 3556 10622
rect 3500 10610 3668 10612
rect 3500 10558 3502 10610
rect 3554 10558 3668 10610
rect 3500 10556 3668 10558
rect 3500 10546 3556 10556
rect 2716 10444 2996 10500
rect 2056 10220 2632 10230
rect 2112 10164 2160 10220
rect 2216 10164 2264 10220
rect 2320 10164 2368 10220
rect 2424 10164 2472 10220
rect 2528 10164 2576 10220
rect 2056 10154 2632 10164
rect 2156 9826 2212 9838
rect 2156 9774 2158 9826
rect 2210 9774 2212 9826
rect 2156 9604 2212 9774
rect 2156 9538 2212 9548
rect 2828 9714 2884 9726
rect 2828 9662 2830 9714
rect 2882 9662 2884 9714
rect 1820 9492 1876 9502
rect 1820 9266 1876 9436
rect 1820 9214 1822 9266
rect 1874 9214 1876 9266
rect 1820 9202 1876 9214
rect 2056 8652 2632 8662
rect 2112 8596 2160 8652
rect 2216 8596 2264 8652
rect 2320 8596 2368 8652
rect 2424 8596 2472 8652
rect 2528 8596 2576 8652
rect 2056 8586 2632 8596
rect 2044 8370 2100 8382
rect 2044 8318 2046 8370
rect 2098 8318 2100 8370
rect 2044 8148 2100 8318
rect 2044 8082 2100 8092
rect 2056 7084 2632 7094
rect 2112 7028 2160 7084
rect 2216 7028 2264 7084
rect 2320 7028 2368 7084
rect 2424 7028 2472 7084
rect 2528 7028 2576 7084
rect 2056 7018 2632 7028
rect 2056 5516 2632 5526
rect 2112 5460 2160 5516
rect 2216 5460 2264 5516
rect 2320 5460 2368 5516
rect 2424 5460 2472 5516
rect 2528 5460 2576 5516
rect 2056 5450 2632 5460
rect 1820 4226 1876 4238
rect 1820 4174 1822 4226
rect 1874 4174 1876 4226
rect 1820 3556 1876 4174
rect 2056 3948 2632 3958
rect 2112 3892 2160 3948
rect 2216 3892 2264 3948
rect 2320 3892 2368 3948
rect 2424 3892 2472 3948
rect 2528 3892 2576 3948
rect 2056 3882 2632 3892
rect 1820 3462 1876 3500
rect 2156 3332 2212 3342
rect 2828 3332 2884 9662
rect 2940 9266 2996 10444
rect 2940 9214 2942 9266
rect 2994 9214 2996 9266
rect 2940 9156 2996 9214
rect 2940 9090 2996 9100
rect 3612 9604 3668 10556
rect 6300 10498 6356 10510
rect 6300 10446 6302 10498
rect 6354 10446 6356 10498
rect 2156 3330 2884 3332
rect 2156 3278 2158 3330
rect 2210 3278 2884 3330
rect 2156 3276 2884 3278
rect 3052 9044 3108 9054
rect 2156 3266 2212 3276
rect 3052 480 3108 8988
rect 3612 9042 3668 9548
rect 4956 9938 5012 9950
rect 4956 9886 4958 9938
rect 5010 9886 5012 9938
rect 4284 9156 4340 9166
rect 4284 9062 4340 9100
rect 3612 8990 3614 9042
rect 3666 8990 3668 9042
rect 3612 8978 3668 8990
rect 4956 8428 5012 9886
rect 6300 9716 6356 10446
rect 6748 10500 6804 10510
rect 6748 10498 6916 10500
rect 6748 10446 6750 10498
rect 6802 10446 6916 10498
rect 6748 10444 6916 10446
rect 6748 10434 6804 10444
rect 6300 9660 6580 9716
rect 5628 9604 5684 9614
rect 5628 9510 5684 9548
rect 5776 9436 6352 9446
rect 5832 9380 5880 9436
rect 5936 9380 5984 9436
rect 6040 9380 6088 9436
rect 6144 9380 6192 9436
rect 6248 9380 6296 9436
rect 5776 9370 6352 9380
rect 4172 8372 5012 8428
rect 6412 8930 6468 8942
rect 6412 8878 6414 8930
rect 6466 8878 6468 8930
rect 4172 8370 4228 8372
rect 4172 8318 4174 8370
rect 4226 8318 4228 8370
rect 4172 8306 4228 8318
rect 4956 8260 5012 8270
rect 4956 8166 5012 8204
rect 5628 8260 5684 8270
rect 5740 8260 5796 8270
rect 5684 8258 5796 8260
rect 5684 8206 5742 8258
rect 5794 8206 5796 8258
rect 5684 8204 5796 8206
rect 5180 7364 5236 7374
rect 5180 7270 5236 7308
rect 5628 7364 5684 8204
rect 5740 8194 5796 8204
rect 5776 7868 6352 7878
rect 5832 7812 5880 7868
rect 5936 7812 5984 7868
rect 6040 7812 6088 7868
rect 6144 7812 6192 7868
rect 6248 7812 6296 7868
rect 5776 7802 6352 7812
rect 6412 7588 6468 8878
rect 6524 8370 6580 9660
rect 6860 9604 6916 10444
rect 6860 8932 6916 9548
rect 6860 8838 6916 8876
rect 8988 8930 9044 8942
rect 8988 8878 8990 8930
rect 9042 8878 9044 8930
rect 6524 8318 6526 8370
rect 6578 8318 6580 8370
rect 6524 8306 6580 8318
rect 8652 8372 8708 8382
rect 8652 8278 8708 8316
rect 8988 8260 9044 8878
rect 11788 8932 11844 8942
rect 11788 8838 11844 8876
rect 12572 8932 12628 8942
rect 8988 8194 9044 8204
rect 9660 8260 9716 8270
rect 9548 8148 9604 8158
rect 9548 8054 9604 8092
rect 9660 7698 9716 8204
rect 9996 8260 10052 8270
rect 9996 8166 10052 8204
rect 10780 8148 10836 8158
rect 10780 8054 10836 8092
rect 9660 7646 9662 7698
rect 9714 7646 9716 7698
rect 6412 7522 6468 7532
rect 6860 7588 6916 7598
rect 6860 7494 6916 7532
rect 5628 7298 5684 7308
rect 6188 7474 6244 7486
rect 6188 7422 6190 7474
rect 6242 7422 6244 7474
rect 6188 7364 6244 7422
rect 6188 7298 6244 7308
rect 8988 7362 9044 7374
rect 8988 7310 8990 7362
rect 9042 7310 9044 7362
rect 5776 6300 6352 6310
rect 5832 6244 5880 6300
rect 5936 6244 5984 6300
rect 6040 6244 6088 6300
rect 6144 6244 6192 6300
rect 6248 6244 6296 6300
rect 5776 6234 6352 6244
rect 8988 5236 9044 7310
rect 9660 7364 9716 7646
rect 9660 7298 9716 7308
rect 11788 7364 11844 7374
rect 11788 7270 11844 7308
rect 12460 6466 12516 6478
rect 12460 6414 12462 6466
rect 12514 6414 12516 6466
rect 12460 6132 12516 6414
rect 12572 6132 12628 8876
rect 12908 8370 12964 22204
rect 16380 22148 16436 22158
rect 14476 19012 14532 19022
rect 14028 10610 14084 10622
rect 14028 10558 14030 10610
rect 14082 10558 14084 10610
rect 13468 10500 13524 10510
rect 14028 10500 14084 10558
rect 13468 10498 14084 10500
rect 13468 10446 13470 10498
rect 13522 10446 14084 10498
rect 13468 10444 14084 10446
rect 13468 9940 13524 10444
rect 13468 8932 13524 9884
rect 13468 8866 13524 8876
rect 12908 8318 12910 8370
rect 12962 8318 12964 8370
rect 12908 8306 12964 8318
rect 13020 8372 13076 8382
rect 13020 6692 13076 8316
rect 13580 8036 13636 8046
rect 13580 7364 13636 7980
rect 13580 7298 13636 7308
rect 13020 6560 13076 6636
rect 13804 6690 13860 6702
rect 13804 6638 13806 6690
rect 13858 6638 13860 6690
rect 12684 6132 12740 6142
rect 12460 6076 12684 6132
rect 12684 5906 12740 6076
rect 13804 6132 13860 6638
rect 14476 6692 14532 18956
rect 15484 16884 15540 16894
rect 14812 10724 14868 10734
rect 14812 10630 14868 10668
rect 14476 6598 14532 6636
rect 13804 6066 13860 6076
rect 13356 6020 13412 6030
rect 13356 5926 13412 5964
rect 12684 5854 12686 5906
rect 12738 5854 12740 5906
rect 12684 5842 12740 5854
rect 15484 5794 15540 16828
rect 16156 12962 16212 12974
rect 16156 12910 16158 12962
rect 16210 12910 16212 12962
rect 15596 12740 15652 12750
rect 16156 12740 16212 12910
rect 15596 12738 16212 12740
rect 15596 12686 15598 12738
rect 15650 12686 16212 12738
rect 15596 12684 16212 12686
rect 15596 9940 15652 12684
rect 15596 9874 15652 9884
rect 16044 9940 16100 9950
rect 16044 9846 16100 9884
rect 15932 6132 15988 6142
rect 15932 6038 15988 6076
rect 16380 6130 16436 22092
rect 17388 20580 17444 36206
rect 38056 35308 38632 35318
rect 38112 35252 38160 35308
rect 38216 35252 38264 35308
rect 38320 35252 38368 35308
rect 38424 35252 38472 35308
rect 38528 35252 38576 35308
rect 38056 35242 38632 35252
rect 38056 33740 38632 33750
rect 38112 33684 38160 33740
rect 38216 33684 38264 33740
rect 38320 33684 38368 33740
rect 38424 33684 38472 33740
rect 38528 33684 38576 33740
rect 38056 33674 38632 33684
rect 38056 32172 38632 32182
rect 38112 32116 38160 32172
rect 38216 32116 38264 32172
rect 38320 32116 38368 32172
rect 38424 32116 38472 32172
rect 38528 32116 38576 32172
rect 38056 32106 38632 32116
rect 38056 30604 38632 30614
rect 38112 30548 38160 30604
rect 38216 30548 38264 30604
rect 38320 30548 38368 30604
rect 38424 30548 38472 30604
rect 38528 30548 38576 30604
rect 38056 30538 38632 30548
rect 39004 29540 39060 29550
rect 38332 29428 38388 29438
rect 37436 29426 38388 29428
rect 37436 29374 38334 29426
rect 38386 29374 38388 29426
rect 37436 29372 38388 29374
rect 36876 29314 36932 29326
rect 36876 29262 36878 29314
rect 36930 29262 36932 29314
rect 32956 28756 33012 28766
rect 30380 28644 30436 28654
rect 29484 27972 29540 27982
rect 27916 25396 27972 25406
rect 17388 16884 17444 20524
rect 20524 21476 20580 21486
rect 17388 16818 17444 16828
rect 19740 19348 19796 19358
rect 19068 13076 19124 13086
rect 19068 12982 19124 13020
rect 16940 12852 16996 12862
rect 16940 12758 16996 12796
rect 19628 12852 19684 12862
rect 19628 12758 19684 12796
rect 18396 12404 18452 12414
rect 18396 11506 18452 12348
rect 18396 11454 18398 11506
rect 18450 11454 18452 11506
rect 18396 11442 18452 11454
rect 17612 11394 17668 11406
rect 17612 11342 17614 11394
rect 17666 11342 17668 11394
rect 17052 11172 17108 11182
rect 17612 11172 17668 11342
rect 17052 11170 17668 11172
rect 17052 11118 17054 11170
rect 17106 11118 17668 11170
rect 17052 11116 17668 11118
rect 16940 11060 16996 11070
rect 16940 10498 16996 11004
rect 16940 10446 16942 10498
rect 16994 10446 16996 10498
rect 16940 10434 16996 10446
rect 16604 9940 16660 9950
rect 16604 9826 16660 9884
rect 17052 9940 17108 11116
rect 17612 10724 17668 10734
rect 17612 10630 17668 10668
rect 19516 10610 19572 10622
rect 19516 10558 19518 10610
rect 19570 10558 19572 10610
rect 17052 9874 17108 9884
rect 18956 10500 19012 10510
rect 19516 10500 19572 10558
rect 18956 10498 19572 10500
rect 18956 10446 18958 10498
rect 19010 10446 19572 10498
rect 18956 10444 19572 10446
rect 18956 9940 19012 10444
rect 19740 10388 19796 19292
rect 20524 11506 20580 21420
rect 22428 21364 22484 21374
rect 20860 18340 20916 18350
rect 20748 12404 20804 12414
rect 20748 12310 20804 12348
rect 20524 11454 20526 11506
rect 20578 11454 20580 11506
rect 20524 11442 20580 11454
rect 20300 10836 20356 10846
rect 20300 10722 20356 10780
rect 20300 10670 20302 10722
rect 20354 10670 20356 10722
rect 20300 10658 20356 10670
rect 18956 9874 19012 9884
rect 19516 10332 19796 10388
rect 19516 9938 19572 10332
rect 19516 9886 19518 9938
rect 19570 9886 19572 9938
rect 19516 9874 19572 9886
rect 16604 9774 16606 9826
rect 16658 9774 16660 9826
rect 16604 9762 16660 9774
rect 17388 9716 17444 9726
rect 17388 9622 17444 9660
rect 20076 9716 20132 9726
rect 20076 9622 20132 9660
rect 19964 9268 20020 9278
rect 16716 9042 16772 9054
rect 16716 8990 16718 9042
rect 16770 8990 16772 9042
rect 16716 8932 16772 8990
rect 19180 9044 19236 9054
rect 19180 8950 19236 8988
rect 19628 9044 19684 9054
rect 19628 8950 19684 8988
rect 16492 8036 16548 8046
rect 16492 7942 16548 7980
rect 16716 7474 16772 8876
rect 17724 8932 17780 8942
rect 17052 8258 17108 8270
rect 17052 8206 17054 8258
rect 17106 8206 17108 8258
rect 17052 8036 17108 8206
rect 17052 7970 17108 7980
rect 17388 8036 17444 8046
rect 16716 7422 16718 7474
rect 16770 7422 16772 7474
rect 16716 7410 16772 7422
rect 16604 6802 16660 6814
rect 16604 6750 16606 6802
rect 16658 6750 16660 6802
rect 16604 6692 16660 6750
rect 16604 6626 16660 6636
rect 17388 6804 17444 7980
rect 17612 7700 17668 7710
rect 17724 7700 17780 8876
rect 19964 8370 20020 9212
rect 19964 8318 19966 8370
rect 20018 8318 20020 8370
rect 19964 8306 20020 8318
rect 17836 8146 17892 8158
rect 17836 8094 17838 8146
rect 17890 8094 17892 8146
rect 17836 8036 17892 8094
rect 17836 7970 17892 7980
rect 20524 8036 20580 8046
rect 20524 7942 20580 7980
rect 17612 7698 17780 7700
rect 17612 7646 17614 7698
rect 17666 7646 17780 7698
rect 17612 7644 17780 7646
rect 17612 7634 17668 7644
rect 20300 6916 20356 6926
rect 16380 6078 16382 6130
rect 16434 6078 16436 6130
rect 16380 6020 16436 6078
rect 16380 5954 16436 5964
rect 15484 5742 15486 5794
rect 15538 5742 15540 5794
rect 15484 5730 15540 5742
rect 8988 5170 9044 5180
rect 16492 5346 16548 5358
rect 16492 5294 16494 5346
rect 16546 5294 16548 5346
rect 16492 5234 16548 5294
rect 17164 5348 17220 5358
rect 17388 5348 17444 6748
rect 17948 6804 18004 6814
rect 17948 6690 18004 6748
rect 17948 6638 17950 6690
rect 18002 6638 18004 6690
rect 17948 6626 18004 6638
rect 18732 6580 18788 6590
rect 18732 6486 18788 6524
rect 17164 5346 17444 5348
rect 17164 5294 17166 5346
rect 17218 5294 17444 5346
rect 17164 5292 17444 5294
rect 17164 5282 17220 5292
rect 16492 5182 16494 5234
rect 16546 5182 16548 5234
rect 16492 5170 16548 5182
rect 16940 5236 16996 5246
rect 16940 5142 16996 5180
rect 17388 5122 17444 5292
rect 18172 5236 18228 5246
rect 18172 5142 18228 5180
rect 20300 5234 20356 6860
rect 20860 6802 20916 18284
rect 21644 11508 21700 11518
rect 21644 11414 21700 11452
rect 22428 10498 22484 21308
rect 22428 10446 22430 10498
rect 22482 10446 22484 10498
rect 22428 10434 22484 10446
rect 22652 20244 22708 20254
rect 20860 6750 20862 6802
rect 20914 6750 20916 6802
rect 20860 6738 20916 6750
rect 21644 10052 21700 10062
rect 21644 6580 21700 9996
rect 22652 10052 22708 20188
rect 25676 19908 25732 19918
rect 23660 19796 23716 19806
rect 23660 13076 23716 19740
rect 23660 13010 23716 13020
rect 23772 15876 23828 15886
rect 23772 11506 23828 15820
rect 23772 11454 23774 11506
rect 23826 11454 23828 11506
rect 23772 11442 23828 11454
rect 25004 15652 25060 15662
rect 24556 11396 24612 11406
rect 24556 11302 24612 11340
rect 24780 11396 24836 11406
rect 22876 10836 22932 10846
rect 22876 10742 22932 10780
rect 24780 10834 24836 11340
rect 24780 10782 24782 10834
rect 24834 10782 24836 10834
rect 24780 10770 24836 10782
rect 22652 9986 22708 9996
rect 25004 9268 25060 15596
rect 25676 11508 25732 19852
rect 27916 16212 27972 25340
rect 28364 22258 28420 22270
rect 28364 22206 28366 22258
rect 28418 22206 28420 22258
rect 28028 22148 28084 22158
rect 28028 22054 28084 22092
rect 27468 16210 27972 16212
rect 27468 16158 27918 16210
rect 27970 16158 27972 16210
rect 27468 16156 27972 16158
rect 27468 16098 27524 16156
rect 27916 16146 27972 16156
rect 28028 21924 28084 21934
rect 27468 16046 27470 16098
rect 27522 16046 27524 16098
rect 27468 16034 27524 16046
rect 27132 15876 27188 15886
rect 27132 15782 27188 15820
rect 27916 12066 27972 12078
rect 27916 12014 27918 12066
rect 27970 12014 27972 12066
rect 25676 11442 25732 11452
rect 25900 11508 25956 11518
rect 25900 11414 25956 11452
rect 25116 11396 25172 11406
rect 25116 11302 25172 11340
rect 27468 11396 27524 11406
rect 27468 10610 27524 11340
rect 27916 11396 27972 12014
rect 28028 11506 28084 21868
rect 28364 21028 28420 22206
rect 28364 20962 28420 20972
rect 28812 20580 28868 20590
rect 28812 20486 28868 20524
rect 29372 20132 29428 20142
rect 29372 20038 29428 20076
rect 29484 18676 29540 27916
rect 30044 26068 30100 26078
rect 29820 21028 29876 21038
rect 29820 20934 29876 20972
rect 30044 18900 30100 26012
rect 30156 20802 30212 20814
rect 30156 20750 30158 20802
rect 30210 20750 30212 20802
rect 30156 20580 30212 20750
rect 30156 20514 30212 20524
rect 30044 18844 30212 18900
rect 30044 18676 30100 18686
rect 29484 18674 30100 18676
rect 29484 18622 30046 18674
rect 30098 18622 30100 18674
rect 29484 18620 30100 18622
rect 29148 18564 29204 18574
rect 29148 18562 29316 18564
rect 29148 18510 29150 18562
rect 29202 18510 29316 18562
rect 29148 18508 29316 18510
rect 29148 18498 29204 18508
rect 28476 16100 28532 16110
rect 28028 11454 28030 11506
rect 28082 11454 28084 11506
rect 28028 11442 28084 11454
rect 28252 15876 28308 15886
rect 27916 11330 27972 11340
rect 28252 10722 28308 15820
rect 28476 12404 28532 16044
rect 28924 15764 28980 15774
rect 28812 13748 28868 13758
rect 28476 12348 28644 12404
rect 28476 12180 28532 12190
rect 28364 12178 28532 12180
rect 28364 12126 28478 12178
rect 28530 12126 28532 12178
rect 28364 12124 28532 12126
rect 28364 11396 28420 12124
rect 28476 12114 28532 12124
rect 28588 11956 28644 12348
rect 28364 11330 28420 11340
rect 28476 11900 28644 11956
rect 28252 10670 28254 10722
rect 28306 10670 28308 10722
rect 28252 10658 28308 10670
rect 27468 10558 27470 10610
rect 27522 10558 27524 10610
rect 27468 10546 27524 10558
rect 25004 9202 25060 9212
rect 23436 8932 23492 8942
rect 23436 7476 23492 8876
rect 23436 7410 23492 7420
rect 24444 7476 24500 7486
rect 21644 6486 21700 6524
rect 22876 7252 22932 7262
rect 20300 5182 20302 5234
rect 20354 5182 20356 5234
rect 20300 5170 20356 5182
rect 22876 5236 22932 7196
rect 22876 5170 22932 5180
rect 17388 5070 17390 5122
rect 17442 5070 17444 5122
rect 17388 5058 17444 5070
rect 24444 5122 24500 7420
rect 26236 7476 26292 7486
rect 26236 7382 26292 7420
rect 28252 7476 28308 7486
rect 28252 7382 28308 7420
rect 26012 6690 26068 6702
rect 26012 6638 26014 6690
rect 26066 6638 26068 6690
rect 25788 5908 25844 5918
rect 26012 5908 26068 6638
rect 26684 6580 26740 6590
rect 26684 6486 26740 6524
rect 25788 5906 26068 5908
rect 25788 5854 25790 5906
rect 25842 5854 26068 5906
rect 25788 5852 26068 5854
rect 25788 5842 25844 5852
rect 24444 5070 24446 5122
rect 24498 5070 24500 5122
rect 24444 5058 24500 5070
rect 26012 5012 26068 5852
rect 26460 5908 26516 5918
rect 26460 5814 26516 5852
rect 25788 4956 26012 5012
rect 5776 4732 6352 4742
rect 5832 4676 5880 4732
rect 5936 4676 5984 4732
rect 6040 4676 6088 4732
rect 6144 4676 6192 4732
rect 6248 4676 6296 4732
rect 5776 4666 6352 4676
rect 22540 4676 22596 4686
rect 20412 4452 20468 4462
rect 20412 4226 20468 4396
rect 22540 4450 22596 4620
rect 24220 4676 24276 4686
rect 24220 4562 24276 4620
rect 24220 4510 24222 4562
rect 24274 4510 24276 4562
rect 24220 4498 24276 4510
rect 22540 4398 22542 4450
rect 22594 4398 22596 4450
rect 22540 4386 22596 4398
rect 23324 4340 23380 4350
rect 23324 4246 23380 4284
rect 23772 4340 23828 4350
rect 23772 4246 23828 4284
rect 25676 4340 25732 4350
rect 25788 4340 25844 4956
rect 26012 4946 26068 4956
rect 28028 5012 28084 5022
rect 28028 4918 28084 4956
rect 26460 4564 26516 4574
rect 26460 4450 26516 4508
rect 26460 4398 26462 4450
rect 26514 4398 26516 4450
rect 26460 4386 26516 4398
rect 25732 4338 25844 4340
rect 25732 4286 25790 4338
rect 25842 4286 25844 4338
rect 25732 4284 25844 4286
rect 20412 4174 20414 4226
rect 20466 4174 20468 4226
rect 20412 4162 20468 4174
rect 25676 3554 25732 4284
rect 25788 4274 25844 4284
rect 28476 3666 28532 11900
rect 28588 11508 28644 11518
rect 28588 11414 28644 11452
rect 28812 6802 28868 13692
rect 28812 6750 28814 6802
rect 28866 6750 28868 6802
rect 28812 6738 28868 6750
rect 28588 5796 28644 5806
rect 28924 5796 28980 15708
rect 29148 15428 29204 15438
rect 29148 15334 29204 15372
rect 29260 12290 29316 18508
rect 29484 18562 29540 18620
rect 30044 18610 30100 18620
rect 29484 18510 29486 18562
rect 29538 18510 29540 18562
rect 29484 18498 29540 18510
rect 29708 17668 29764 17678
rect 29708 17574 29764 17612
rect 30156 17556 30212 18844
rect 30380 17778 30436 28588
rect 31500 27860 31556 27870
rect 30828 25284 30884 25294
rect 30380 17726 30382 17778
rect 30434 17726 30436 17778
rect 30380 17668 30436 17726
rect 30380 17602 30436 17612
rect 30492 23380 30548 23390
rect 30044 17500 30212 17556
rect 29932 17442 29988 17454
rect 29932 17390 29934 17442
rect 29986 17390 29988 17442
rect 29932 16324 29988 17390
rect 29932 16258 29988 16268
rect 30044 15538 30100 17500
rect 30380 16324 30436 16334
rect 30044 15486 30046 15538
rect 30098 15486 30100 15538
rect 29484 15426 29540 15438
rect 29484 15374 29486 15426
rect 29538 15374 29540 15426
rect 29484 13524 29540 15374
rect 30044 15428 30100 15486
rect 30044 15362 30100 15372
rect 30156 15874 30212 15886
rect 30156 15822 30158 15874
rect 30210 15822 30212 15874
rect 29484 13458 29540 13468
rect 30044 14644 30100 14654
rect 29260 12238 29262 12290
rect 29314 12238 29316 12290
rect 29260 12226 29316 12238
rect 29596 12962 29652 12974
rect 29596 12910 29598 12962
rect 29650 12910 29652 12962
rect 29596 11396 29652 12910
rect 29596 9828 29652 11340
rect 29932 9828 29988 9838
rect 29596 9826 29932 9828
rect 29596 9774 29598 9826
rect 29650 9774 29932 9826
rect 29596 9772 29932 9774
rect 29596 9762 29652 9772
rect 29932 9042 29988 9772
rect 29932 8990 29934 9042
rect 29986 8990 29988 9042
rect 29932 8978 29988 8990
rect 29148 7476 29204 7486
rect 29036 5908 29092 5918
rect 29036 5814 29092 5852
rect 28588 5794 28980 5796
rect 28588 5742 28590 5794
rect 28642 5742 28980 5794
rect 28588 5740 28980 5742
rect 28588 5730 28644 5740
rect 28700 5236 28756 5246
rect 29148 5236 29204 7420
rect 29596 6580 29652 6590
rect 29596 6486 29652 6524
rect 29932 6466 29988 6478
rect 29932 6414 29934 6466
rect 29986 6414 29988 6466
rect 28700 5234 29204 5236
rect 28700 5182 28702 5234
rect 28754 5182 29204 5234
rect 28700 5180 29204 5182
rect 29484 5794 29540 5806
rect 29484 5742 29486 5794
rect 29538 5742 29540 5794
rect 28700 5170 28756 5180
rect 29260 5012 29316 5022
rect 29260 4562 29316 4956
rect 29484 5012 29540 5742
rect 29484 4946 29540 4956
rect 29708 5122 29764 5134
rect 29708 5070 29710 5122
rect 29762 5070 29764 5122
rect 29708 5012 29764 5070
rect 29708 4946 29764 4956
rect 29932 5012 29988 6414
rect 29932 4946 29988 4956
rect 29260 4510 29262 4562
rect 29314 4510 29316 4562
rect 28588 4226 28644 4238
rect 28588 4174 28590 4226
rect 28642 4174 28644 4226
rect 28588 3892 28644 4174
rect 28588 3836 29092 3892
rect 29036 3778 29092 3836
rect 29036 3726 29038 3778
rect 29090 3726 29092 3778
rect 29036 3714 29092 3726
rect 28476 3614 28478 3666
rect 28530 3614 28532 3666
rect 28476 3602 28532 3614
rect 29260 3668 29316 4510
rect 29708 4564 29764 4574
rect 29708 4470 29764 4508
rect 30044 3778 30100 14588
rect 30156 13524 30212 15822
rect 30156 13468 30324 13524
rect 30268 11508 30324 13468
rect 30380 13074 30436 16268
rect 30492 16098 30548 23324
rect 30828 20690 30884 25228
rect 31500 20916 31556 27804
rect 30940 20914 31556 20916
rect 30940 20862 31502 20914
rect 31554 20862 31556 20914
rect 30940 20860 31556 20862
rect 30940 20802 30996 20860
rect 31500 20850 31556 20860
rect 31612 27748 31668 27758
rect 30940 20750 30942 20802
rect 30994 20750 30996 20802
rect 30940 20738 30996 20750
rect 31612 20692 31668 27692
rect 32396 26180 32452 26190
rect 30828 20638 30830 20690
rect 30882 20638 30884 20690
rect 30828 20132 30884 20638
rect 30828 20066 30884 20076
rect 31388 20636 31668 20692
rect 31836 23156 31892 23166
rect 31276 19124 31332 19134
rect 31276 19030 31332 19068
rect 30940 19012 30996 19022
rect 30940 19010 31108 19012
rect 30940 18958 30942 19010
rect 30994 18958 31108 19010
rect 30940 18956 31108 18958
rect 30940 18946 30996 18956
rect 30940 18562 30996 18574
rect 30940 18510 30942 18562
rect 30994 18510 30996 18562
rect 30940 16436 30996 18510
rect 30940 16370 30996 16380
rect 31052 16212 31108 18956
rect 31276 18564 31332 18574
rect 31276 18470 31332 18508
rect 31276 17442 31332 17454
rect 31276 17390 31278 17442
rect 31330 17390 31332 17442
rect 30492 16046 30494 16098
rect 30546 16046 30548 16098
rect 30492 15540 30548 16046
rect 30940 16156 31108 16212
rect 31164 16994 31220 17006
rect 31164 16942 31166 16994
rect 31218 16942 31220 16994
rect 30828 15540 30884 15550
rect 30492 15538 30884 15540
rect 30492 15486 30830 15538
rect 30882 15486 30884 15538
rect 30492 15484 30884 15486
rect 30828 15474 30884 15484
rect 30380 13022 30382 13074
rect 30434 13022 30436 13074
rect 30380 13010 30436 13022
rect 30492 13524 30548 13534
rect 30380 11508 30436 11518
rect 30268 11506 30436 11508
rect 30268 11454 30382 11506
rect 30434 11454 30436 11506
rect 30268 11452 30436 11454
rect 30380 11442 30436 11452
rect 30380 10612 30436 10622
rect 30380 10498 30436 10556
rect 30380 10446 30382 10498
rect 30434 10446 30436 10498
rect 30380 10434 30436 10446
rect 30380 9940 30436 9950
rect 30492 9940 30548 13468
rect 30940 12740 30996 16156
rect 31052 15876 31108 15886
rect 31052 15782 31108 15820
rect 30940 12674 30996 12684
rect 31052 15540 31108 15550
rect 30380 9938 30548 9940
rect 30380 9886 30382 9938
rect 30434 9886 30548 9938
rect 30380 9884 30548 9886
rect 30828 10498 30884 10510
rect 30828 10446 30830 10498
rect 30882 10446 30884 10498
rect 30380 9874 30436 9884
rect 30828 9828 30884 10446
rect 30716 8932 30772 8942
rect 30716 8838 30772 8876
rect 30828 7586 30884 9772
rect 31052 9716 31108 15484
rect 31164 11508 31220 16942
rect 31164 11442 31220 11452
rect 31276 10836 31332 17390
rect 31388 16212 31444 20636
rect 31836 18788 31892 23100
rect 32172 20580 32228 20590
rect 31836 18732 32004 18788
rect 31836 18564 31892 18574
rect 31724 18562 31892 18564
rect 31724 18510 31838 18562
rect 31890 18510 31892 18562
rect 31724 18508 31892 18510
rect 31612 17780 31668 17790
rect 31612 17666 31668 17724
rect 31612 17614 31614 17666
rect 31666 17614 31668 17666
rect 31612 17602 31668 17614
rect 31500 17108 31556 17118
rect 31500 16994 31556 17052
rect 31500 16942 31502 16994
rect 31554 16942 31556 16994
rect 31500 16930 31556 16942
rect 31388 16156 31556 16212
rect 31388 15988 31444 15998
rect 31388 15894 31444 15932
rect 31500 15148 31556 16156
rect 31388 15092 31556 15148
rect 31724 15148 31780 18508
rect 31836 18498 31892 18508
rect 31948 18340 32004 18732
rect 32172 18562 32228 20524
rect 32172 18510 32174 18562
rect 32226 18510 32228 18562
rect 32172 18498 32228 18510
rect 32284 20130 32340 20142
rect 32284 20078 32286 20130
rect 32338 20078 32340 20130
rect 31836 18284 32004 18340
rect 31836 16210 31892 18284
rect 32060 17780 32116 17790
rect 32060 17686 32116 17724
rect 32060 17108 32116 17118
rect 32060 17014 32116 17052
rect 31836 16158 31838 16210
rect 31890 16158 31892 16210
rect 31836 15988 31892 16158
rect 31836 15922 31892 15932
rect 31724 15092 31892 15148
rect 31388 12066 31444 15092
rect 31836 12404 31892 15092
rect 31836 12338 31892 12348
rect 31388 12014 31390 12066
rect 31442 12014 31444 12066
rect 31388 12002 31444 12014
rect 31836 12180 31892 12190
rect 31836 12066 31892 12124
rect 31836 12014 31838 12066
rect 31890 12014 31892 12066
rect 31276 10770 31332 10780
rect 31836 9828 31892 12014
rect 32284 10724 32340 20078
rect 32284 10658 32340 10668
rect 32396 9940 32452 26124
rect 32620 20018 32676 20030
rect 32620 19966 32622 20018
rect 32674 19966 32676 20018
rect 32620 18340 32676 19966
rect 32620 18274 32676 18284
rect 32844 16100 32900 16110
rect 32844 16006 32900 16044
rect 32956 15148 33012 28700
rect 36764 28756 36820 28766
rect 36876 28756 36932 29262
rect 37324 29316 37380 29326
rect 37436 29316 37492 29372
rect 38332 29362 38388 29372
rect 38780 29426 38836 29438
rect 38780 29374 38782 29426
rect 38834 29374 38836 29426
rect 37324 29314 37492 29316
rect 37324 29262 37326 29314
rect 37378 29262 37492 29314
rect 37324 29260 37492 29262
rect 37324 29250 37380 29260
rect 36820 28700 36932 28756
rect 36764 28662 36820 28700
rect 35196 28084 35252 28094
rect 34636 27636 34692 27646
rect 34636 25396 34692 27580
rect 34636 25330 34692 25340
rect 35196 25284 35252 28028
rect 36652 28084 36708 28094
rect 36652 27990 36708 28028
rect 36204 27748 36260 27758
rect 36204 27654 36260 27692
rect 37436 27748 37492 29260
rect 37996 29204 38052 29214
rect 37884 29202 38052 29204
rect 37884 29150 37998 29202
rect 38050 29150 38052 29202
rect 37884 29148 38052 29150
rect 37660 28084 37716 28094
rect 37660 27858 37716 28028
rect 37884 27972 37940 29148
rect 37996 29138 38052 29148
rect 38056 29036 38632 29046
rect 38112 28980 38160 29036
rect 38216 28980 38264 29036
rect 38320 28980 38368 29036
rect 38424 28980 38472 29036
rect 38528 28980 38576 29036
rect 38056 28970 38632 28980
rect 38332 28756 38388 28766
rect 38332 28662 38388 28700
rect 37996 28644 38052 28654
rect 37996 28550 38052 28588
rect 38556 28530 38612 28542
rect 38556 28478 38558 28530
rect 38610 28478 38612 28530
rect 37884 27906 37940 27916
rect 38220 27972 38276 27982
rect 37660 27806 37662 27858
rect 37714 27806 37716 27858
rect 37660 27794 37716 27806
rect 38108 27860 38164 27870
rect 38108 27766 38164 27804
rect 37436 27682 37492 27692
rect 38220 27748 38276 27916
rect 38556 27860 38612 28478
rect 38556 27794 38612 27804
rect 38780 28532 38836 29374
rect 39004 28644 39060 29484
rect 39676 29316 39732 29326
rect 39676 29314 39844 29316
rect 39676 29262 39678 29314
rect 39730 29262 39844 29314
rect 39676 29260 39844 29262
rect 39676 29250 39732 29260
rect 39004 28578 39060 28588
rect 39676 28866 39732 28878
rect 39676 28814 39678 28866
rect 39730 28814 39732 28866
rect 38780 27860 38836 28476
rect 38220 27682 38276 27692
rect 37324 27636 37380 27646
rect 37324 27542 37380 27580
rect 38056 27468 38632 27478
rect 38112 27412 38160 27468
rect 38216 27412 38264 27468
rect 38320 27412 38368 27468
rect 38424 27412 38472 27468
rect 38528 27412 38576 27468
rect 38056 27402 38632 27412
rect 38780 27186 38836 27804
rect 38780 27134 38782 27186
rect 38834 27134 38836 27186
rect 38780 27122 38836 27134
rect 38892 28530 38948 28542
rect 38892 28478 38894 28530
rect 38946 28478 38948 28530
rect 38892 28420 38948 28478
rect 39676 28420 39732 28814
rect 39788 28532 39844 29260
rect 40236 28866 40292 41916
rect 41776 40796 42352 40806
rect 41832 40740 41880 40796
rect 41936 40740 41984 40796
rect 42040 40740 42088 40796
rect 42144 40740 42192 40796
rect 42248 40740 42296 40796
rect 41776 40730 42352 40740
rect 41776 39228 42352 39238
rect 41832 39172 41880 39228
rect 41936 39172 41984 39228
rect 42040 39172 42088 39228
rect 42144 39172 42192 39228
rect 42248 39172 42296 39228
rect 41776 39162 42352 39172
rect 40236 28814 40238 28866
rect 40290 28814 40292 28866
rect 40236 28802 40292 28814
rect 41132 38724 41188 38734
rect 39788 28466 39844 28476
rect 40124 28532 40180 28542
rect 40124 28438 40180 28476
rect 38892 28418 39732 28420
rect 38892 28366 39678 28418
rect 39730 28366 39732 28418
rect 38892 28364 39732 28366
rect 35196 25218 35252 25228
rect 37100 26404 37156 26414
rect 37100 26178 37156 26348
rect 37100 26126 37102 26178
rect 37154 26126 37156 26178
rect 37100 24724 37156 26126
rect 37548 26180 37604 26190
rect 37548 26086 37604 26124
rect 38556 26180 38612 26190
rect 38220 26068 38276 26106
rect 38556 26086 38612 26124
rect 38892 26180 38948 28364
rect 39676 28354 39732 28364
rect 39116 27860 39172 27870
rect 39116 27766 39172 27804
rect 39676 27860 39732 27870
rect 39676 27858 39844 27860
rect 39676 27806 39678 27858
rect 39730 27806 39844 27858
rect 39676 27804 39844 27806
rect 39676 27794 39732 27804
rect 39676 26964 39732 26974
rect 39340 26962 39732 26964
rect 39340 26910 39678 26962
rect 39730 26910 39732 26962
rect 39340 26908 39732 26910
rect 39116 26404 39172 26414
rect 39116 26310 39172 26348
rect 39340 26292 39396 26908
rect 39676 26898 39732 26908
rect 39788 26852 39844 27804
rect 39788 26786 39844 26796
rect 40236 26852 40292 26862
rect 40236 26758 40292 26796
rect 40796 26852 40852 26862
rect 38892 26114 38948 26124
rect 39228 26290 39396 26292
rect 39228 26238 39342 26290
rect 39394 26238 39396 26290
rect 39228 26236 39396 26238
rect 38220 26002 38276 26012
rect 38056 25900 38632 25910
rect 38112 25844 38160 25900
rect 38216 25844 38264 25900
rect 38320 25844 38368 25900
rect 38424 25844 38472 25900
rect 38528 25844 38576 25900
rect 38056 25834 38632 25844
rect 39116 24836 39172 24846
rect 38444 24724 38500 24734
rect 37100 24722 38500 24724
rect 37100 24670 38446 24722
rect 38498 24670 38500 24722
rect 37100 24668 38500 24670
rect 36988 24610 37044 24622
rect 36988 24558 36990 24610
rect 37042 24558 37044 24610
rect 36988 23940 37044 24558
rect 36764 23716 36820 23726
rect 36988 23716 37044 23884
rect 36652 23714 37044 23716
rect 36652 23662 36766 23714
rect 36818 23662 37044 23714
rect 36652 23660 37044 23662
rect 37436 24610 37492 24668
rect 38444 24658 38500 24668
rect 37436 24558 37438 24610
rect 37490 24558 37492 24610
rect 34972 22148 35028 22158
rect 33404 21812 33460 21822
rect 32508 15092 33012 15148
rect 33180 20578 33236 20590
rect 33180 20526 33182 20578
rect 33234 20526 33236 20578
rect 32508 13074 32564 15092
rect 32508 13022 32510 13074
rect 32562 13022 32564 13074
rect 32508 13010 32564 13022
rect 32620 13524 32676 13534
rect 32508 11732 32564 11742
rect 32508 11506 32564 11676
rect 32508 11454 32510 11506
rect 32562 11454 32564 11506
rect 32508 11442 32564 11454
rect 32508 9940 32564 9950
rect 32396 9938 32564 9940
rect 32396 9886 32510 9938
rect 32562 9886 32564 9938
rect 32396 9884 32564 9886
rect 32508 9874 32564 9884
rect 31836 9762 31892 9772
rect 31052 9650 31108 9660
rect 32620 8932 32676 13468
rect 32956 12740 33012 12750
rect 32732 12738 33012 12740
rect 32732 12686 32958 12738
rect 33010 12686 33012 12738
rect 32732 12684 33012 12686
rect 32732 12402 32788 12684
rect 32956 12674 33012 12684
rect 32732 12350 32734 12402
rect 32786 12350 32788 12402
rect 32732 12180 32788 12350
rect 32732 12114 32788 12124
rect 33180 11620 33236 20526
rect 33292 15874 33348 15886
rect 33292 15822 33294 15874
rect 33346 15822 33348 15874
rect 33292 15764 33348 15822
rect 33292 15698 33348 15708
rect 33292 14756 33348 14766
rect 33292 14642 33348 14700
rect 33292 14590 33294 14642
rect 33346 14590 33348 14642
rect 33292 14578 33348 14590
rect 33404 11732 33460 21756
rect 33516 20690 33572 20702
rect 33516 20638 33518 20690
rect 33570 20638 33572 20690
rect 33516 18676 33572 20638
rect 34300 20692 34356 20702
rect 33628 20244 33684 20254
rect 33628 20150 33684 20188
rect 33964 20018 34020 20030
rect 33964 19966 33966 20018
rect 34018 19966 34020 20018
rect 33740 19012 33796 19022
rect 33516 18610 33572 18620
rect 33628 19010 33796 19012
rect 33628 18958 33742 19010
rect 33794 18958 33796 19010
rect 33628 18956 33796 18958
rect 33516 16100 33572 16110
rect 33516 15538 33572 16044
rect 33516 15486 33518 15538
rect 33570 15486 33572 15538
rect 33516 15474 33572 15486
rect 33628 14420 33684 18956
rect 33740 18900 33796 18956
rect 33740 18834 33796 18844
rect 33964 18004 34020 19966
rect 34300 19458 34356 20636
rect 34524 20132 34580 20142
rect 34524 20130 34692 20132
rect 34524 20078 34526 20130
rect 34578 20078 34692 20130
rect 34524 20076 34692 20078
rect 34524 20066 34580 20076
rect 34300 19406 34302 19458
rect 34354 19406 34356 19458
rect 34300 19394 34356 19406
rect 34188 19122 34244 19134
rect 34188 19070 34190 19122
rect 34242 19070 34244 19122
rect 34188 19012 34244 19070
rect 34188 18946 34244 18956
rect 34300 19010 34356 19022
rect 34300 18958 34302 19010
rect 34354 18958 34356 19010
rect 34300 18900 34356 18958
rect 34300 18834 34356 18844
rect 33964 17938 34020 17948
rect 33964 17442 34020 17454
rect 34524 17444 34580 17454
rect 33964 17390 33966 17442
rect 34018 17390 34020 17442
rect 33964 16884 34020 17390
rect 33964 16818 34020 16828
rect 34076 17442 34580 17444
rect 34076 17390 34526 17442
rect 34578 17390 34580 17442
rect 34076 17388 34580 17390
rect 34076 15148 34132 17388
rect 34524 17378 34580 17388
rect 34636 17220 34692 20076
rect 34748 20018 34804 20030
rect 34748 19966 34750 20018
rect 34802 19966 34804 20018
rect 34748 17892 34804 19966
rect 34860 19012 34916 19022
rect 34860 18918 34916 18956
rect 34748 17826 34804 17836
rect 34860 18452 34916 18462
rect 34524 17164 34692 17220
rect 34748 17666 34804 17678
rect 34748 17614 34750 17666
rect 34802 17614 34804 17666
rect 34300 16996 34356 17006
rect 34300 16770 34356 16940
rect 34300 16718 34302 16770
rect 34354 16718 34356 16770
rect 34188 16100 34244 16110
rect 34188 15986 34244 16044
rect 34188 15934 34190 15986
rect 34242 15934 34244 15986
rect 34188 15922 34244 15934
rect 34300 15764 34356 16718
rect 34300 15698 34356 15708
rect 34412 15986 34468 15998
rect 34412 15934 34414 15986
rect 34466 15934 34468 15986
rect 33964 15092 34132 15148
rect 34300 15540 34356 15550
rect 34300 15426 34356 15484
rect 34300 15374 34302 15426
rect 34354 15374 34356 15426
rect 33740 14756 33796 14766
rect 33740 14642 33796 14700
rect 33740 14590 33742 14642
rect 33794 14590 33796 14642
rect 33740 14578 33796 14590
rect 33628 14364 33796 14420
rect 33404 11666 33460 11676
rect 33180 11564 33348 11620
rect 33180 11394 33236 11406
rect 33180 11342 33182 11394
rect 33234 11342 33236 11394
rect 33180 11284 33236 11342
rect 32732 11228 33180 11284
rect 32732 10834 32788 11228
rect 32732 10782 32734 10834
rect 32786 10782 32788 10834
rect 32732 10770 32788 10782
rect 32956 9940 33012 11228
rect 33180 11218 33236 11228
rect 32956 9808 33012 9884
rect 32844 8932 32900 8942
rect 32620 8930 32900 8932
rect 32620 8878 32846 8930
rect 32898 8878 32900 8930
rect 32620 8876 32900 8878
rect 32844 8866 32900 8876
rect 33292 8428 33348 11564
rect 33516 9940 33572 9950
rect 33516 9846 33572 9884
rect 33516 9380 33572 9390
rect 33516 9266 33572 9324
rect 33516 9214 33518 9266
rect 33570 9214 33572 9266
rect 33516 8932 33572 9214
rect 33516 8866 33572 8876
rect 33740 8428 33796 14364
rect 33964 11956 34020 15092
rect 34300 14756 34356 15374
rect 34412 15316 34468 15934
rect 34412 15250 34468 15260
rect 34524 14980 34580 17164
rect 34748 16996 34804 17614
rect 34860 17668 34916 18396
rect 34860 17602 34916 17612
rect 34300 14690 34356 14700
rect 34412 14924 34580 14980
rect 34636 16940 34804 16996
rect 34076 13636 34132 13646
rect 34076 13542 34132 13580
rect 34412 12180 34468 14924
rect 34524 14756 34580 14766
rect 34636 14756 34692 16940
rect 34860 16884 34916 16894
rect 34748 16828 34860 16884
rect 34748 16770 34804 16828
rect 34860 16818 34916 16828
rect 34748 16718 34750 16770
rect 34802 16718 34804 16770
rect 34748 16706 34804 16718
rect 34972 16324 35028 22092
rect 36428 21476 36484 21486
rect 36428 21382 36484 21420
rect 36652 20692 36708 23660
rect 36764 23650 36820 23660
rect 36876 23268 36932 23278
rect 36876 23042 36932 23212
rect 36876 22990 36878 23042
rect 36930 22990 36932 23042
rect 36764 21476 36820 21486
rect 36764 21028 36820 21420
rect 36876 21474 36932 22990
rect 37324 23042 37380 23054
rect 37324 22990 37326 23042
rect 37378 22990 37380 23042
rect 37324 22932 37380 22990
rect 37324 21924 37380 22876
rect 37324 21858 37380 21868
rect 37436 21812 37492 24558
rect 38108 24500 38164 24510
rect 37884 24498 38164 24500
rect 37884 24446 38110 24498
rect 38162 24446 38164 24498
rect 37884 24444 38164 24446
rect 37884 23380 37940 24444
rect 38108 24434 38164 24444
rect 38056 24332 38632 24342
rect 38112 24276 38160 24332
rect 38216 24276 38264 24332
rect 38320 24276 38368 24332
rect 38424 24276 38472 24332
rect 38528 24276 38576 24332
rect 38056 24266 38632 24276
rect 39116 24164 39172 24780
rect 39116 24098 39172 24108
rect 39228 24722 39284 26236
rect 39340 26226 39396 26236
rect 40348 25618 40404 25630
rect 40348 25566 40350 25618
rect 40402 25566 40404 25618
rect 39228 24670 39230 24722
rect 39282 24670 39284 24722
rect 38332 23940 38388 23950
rect 38332 23846 38388 23884
rect 39116 23940 39172 23950
rect 39228 23940 39284 24670
rect 39116 23938 39284 23940
rect 39116 23886 39118 23938
rect 39170 23886 39284 23938
rect 39116 23884 39284 23886
rect 39676 25284 39732 25294
rect 39676 24050 39732 25228
rect 40348 24052 40404 25566
rect 39676 23998 39678 24050
rect 39730 23998 39732 24050
rect 39004 23826 39060 23838
rect 39004 23774 39006 23826
rect 39058 23774 39060 23826
rect 37884 23314 37940 23324
rect 37996 23714 38052 23726
rect 37996 23662 37998 23714
rect 38050 23662 38052 23714
rect 37996 23156 38052 23662
rect 37996 23090 38052 23100
rect 38332 23492 38388 23502
rect 37996 22932 38052 22942
rect 37436 21746 37492 21756
rect 37772 22930 38052 22932
rect 37772 22878 37998 22930
rect 38050 22878 38052 22930
rect 37772 22876 38052 22878
rect 36876 21422 36878 21474
rect 36930 21422 36932 21474
rect 36876 21364 36932 21422
rect 36876 21298 36932 21308
rect 37548 21362 37604 21374
rect 37548 21310 37550 21362
rect 37602 21310 37604 21362
rect 36764 20914 36820 20972
rect 36764 20862 36766 20914
rect 36818 20862 36820 20914
rect 36764 20850 36820 20862
rect 36652 20636 36932 20692
rect 36316 20580 36372 20590
rect 36316 20578 36484 20580
rect 36316 20526 36318 20578
rect 36370 20526 36484 20578
rect 36316 20524 36484 20526
rect 36316 20514 36372 20524
rect 36428 20244 36484 20524
rect 35980 19906 36036 19918
rect 35980 19854 35982 19906
rect 36034 19854 36036 19906
rect 35980 19796 36036 19854
rect 35980 19730 36036 19740
rect 36428 19906 36484 20188
rect 36428 19854 36430 19906
rect 36482 19854 36484 19906
rect 36428 19348 36484 19854
rect 36428 19282 36484 19292
rect 36764 19796 36820 19806
rect 36764 19460 36820 19740
rect 36764 19346 36820 19404
rect 36764 19294 36766 19346
rect 36818 19294 36820 19346
rect 36764 19282 36820 19294
rect 35756 19010 35812 19022
rect 35756 18958 35758 19010
rect 35810 18958 35812 19010
rect 35756 18788 35812 18958
rect 36204 19012 36260 19022
rect 36204 18918 36260 18956
rect 35420 18562 35476 18574
rect 35420 18510 35422 18562
rect 35474 18510 35476 18562
rect 34860 16268 35028 16324
rect 35084 18452 35140 18462
rect 35084 16322 35140 18396
rect 35420 18116 35476 18510
rect 35644 18452 35700 18462
rect 35644 18358 35700 18396
rect 35420 18050 35476 18060
rect 35532 18004 35588 18014
rect 35420 17892 35476 17902
rect 35084 16270 35086 16322
rect 35138 16270 35140 16322
rect 34748 16098 34804 16110
rect 34748 16046 34750 16098
rect 34802 16046 34804 16098
rect 34748 15764 34804 16046
rect 34748 15698 34804 15708
rect 34860 15540 34916 16268
rect 35084 16258 35140 16270
rect 35308 17556 35364 17566
rect 34860 15474 34916 15484
rect 34972 16100 35028 16110
rect 34748 15426 34804 15438
rect 34748 15374 34750 15426
rect 34802 15374 34804 15426
rect 34748 15316 34804 15374
rect 34748 15250 34804 15260
rect 34972 15314 35028 16044
rect 35308 15538 35364 17500
rect 35420 17106 35476 17836
rect 35532 17890 35588 17948
rect 35532 17838 35534 17890
rect 35586 17838 35588 17890
rect 35532 17826 35588 17838
rect 35756 17668 35812 18732
rect 36764 18788 36820 18798
rect 36652 18452 36708 18462
rect 36428 18340 36484 18350
rect 36428 18246 36484 18284
rect 36204 18116 36260 18126
rect 35420 17054 35422 17106
rect 35474 17054 35476 17106
rect 35420 17042 35476 17054
rect 35532 17612 35812 17668
rect 35868 17668 35924 17678
rect 35532 16884 35588 17612
rect 35308 15486 35310 15538
rect 35362 15486 35364 15538
rect 35308 15474 35364 15486
rect 35420 16828 35588 16884
rect 35644 17444 35700 17454
rect 34972 15262 34974 15314
rect 35026 15262 35028 15314
rect 34972 15250 35028 15262
rect 34524 14754 34692 14756
rect 34524 14702 34526 14754
rect 34578 14702 34692 14754
rect 34524 14700 34692 14702
rect 34860 14756 34916 14766
rect 34524 14690 34580 14700
rect 34860 14662 34916 14700
rect 34412 12124 34580 12180
rect 33964 11900 34244 11956
rect 33852 11508 33908 11518
rect 33852 11414 33908 11452
rect 34076 11396 34132 11406
rect 33964 11340 34076 11396
rect 33964 10610 34020 11340
rect 34076 11330 34132 11340
rect 33964 10558 33966 10610
rect 34018 10558 34020 10610
rect 33964 9268 34020 10558
rect 33964 9136 34020 9212
rect 33180 8372 33348 8428
rect 33628 8372 33796 8428
rect 33180 8036 33236 8372
rect 33180 7970 33236 7980
rect 30828 7534 30830 7586
rect 30882 7534 30884 7586
rect 30828 7522 30884 7534
rect 33628 6692 33684 8372
rect 33628 6626 33684 6636
rect 33068 6020 33124 6030
rect 32508 5234 32564 5246
rect 32508 5182 32510 5234
rect 32562 5182 32564 5234
rect 30380 5124 30436 5134
rect 30380 5030 30436 5068
rect 32508 4788 32564 5182
rect 33068 5234 33124 5964
rect 33068 5182 33070 5234
rect 33122 5182 33124 5234
rect 33068 5124 33124 5182
rect 33068 5058 33124 5068
rect 33852 5122 33908 5134
rect 33852 5070 33854 5122
rect 33906 5070 33908 5122
rect 32508 4722 32564 4732
rect 33516 5012 33572 5022
rect 33516 4562 33572 4956
rect 33852 5012 33908 5070
rect 33908 4956 34132 5012
rect 33852 4946 33908 4956
rect 33516 4510 33518 4562
rect 33570 4510 33572 4562
rect 33516 4498 33572 4510
rect 34076 4562 34132 4956
rect 34076 4510 34078 4562
rect 34130 4510 34132 4562
rect 34076 4340 34132 4510
rect 34188 4564 34244 11900
rect 34524 8428 34580 12124
rect 35308 12178 35364 12190
rect 35308 12126 35310 12178
rect 35362 12126 35364 12178
rect 34636 12068 34692 12078
rect 35308 12068 35364 12126
rect 34636 12066 35364 12068
rect 34636 12014 34638 12066
rect 34690 12014 35364 12066
rect 34636 12012 35364 12014
rect 34636 12002 34692 12012
rect 35308 11396 35364 12012
rect 35308 11330 35364 11340
rect 35420 11060 35476 16828
rect 35644 16212 35700 17388
rect 35868 17220 35924 17612
rect 35868 17154 35924 17164
rect 35756 16884 35812 16894
rect 35812 16828 35924 16884
rect 35756 16790 35812 16828
rect 35644 16210 35812 16212
rect 35644 16158 35646 16210
rect 35698 16158 35812 16210
rect 35644 16156 35812 16158
rect 35644 16146 35700 16156
rect 35644 15316 35700 15326
rect 35532 15092 35588 15102
rect 35532 14418 35588 15036
rect 35644 14530 35700 15260
rect 35756 15092 35812 16156
rect 35756 15026 35812 15036
rect 35868 14980 35924 16828
rect 36204 16660 36260 18060
rect 36428 17668 36484 17678
rect 36652 17668 36708 18396
rect 36764 18450 36820 18732
rect 36764 18398 36766 18450
rect 36818 18398 36820 18450
rect 36764 18386 36820 18398
rect 36876 18228 36932 20636
rect 37436 20244 37492 20254
rect 37436 20018 37492 20188
rect 37436 19966 37438 20018
rect 37490 19966 37492 20018
rect 37436 19954 37492 19966
rect 37100 19794 37156 19806
rect 37100 19742 37102 19794
rect 37154 19742 37156 19794
rect 37100 18564 37156 19742
rect 37324 19012 37380 19022
rect 37100 18498 37156 18508
rect 37212 18676 37268 18686
rect 36428 17554 36484 17612
rect 36428 17502 36430 17554
rect 36482 17502 36484 17554
rect 36316 16996 36372 17006
rect 36316 16902 36372 16940
rect 36428 16884 36484 17502
rect 36428 16818 36484 16828
rect 36540 17666 36708 17668
rect 36540 17614 36654 17666
rect 36706 17614 36708 17666
rect 36540 17612 36708 17614
rect 36540 16882 36596 17612
rect 36652 17602 36708 17612
rect 36764 18172 36932 18228
rect 36540 16830 36542 16882
rect 36594 16830 36596 16882
rect 36540 16818 36596 16830
rect 36204 16604 36596 16660
rect 36428 16100 36484 16110
rect 36092 16098 36484 16100
rect 36092 16046 36430 16098
rect 36482 16046 36484 16098
rect 36092 16044 36484 16046
rect 36092 15538 36148 16044
rect 36428 16034 36484 16044
rect 36092 15486 36094 15538
rect 36146 15486 36148 15538
rect 36092 15474 36148 15486
rect 36204 15874 36260 15886
rect 36204 15822 36206 15874
rect 36258 15822 36260 15874
rect 36204 15148 36260 15822
rect 36204 15092 36372 15148
rect 36204 14980 36260 14990
rect 35868 14924 36036 14980
rect 35980 14532 36036 14924
rect 35644 14478 35646 14530
rect 35698 14478 35700 14530
rect 35644 14466 35700 14478
rect 35868 14476 36036 14532
rect 36092 14756 36148 14766
rect 35532 14366 35534 14418
rect 35586 14366 35588 14418
rect 35532 13636 35588 14366
rect 35532 13570 35588 13580
rect 35420 10994 35476 11004
rect 34636 10724 34692 10734
rect 34636 10630 34692 10668
rect 35196 9268 35252 9278
rect 35196 9174 35252 9212
rect 35756 9268 35812 9278
rect 35756 9042 35812 9212
rect 35756 8990 35758 9042
rect 35810 8990 35812 9042
rect 35756 8978 35812 8990
rect 35868 8428 35924 14476
rect 35980 14308 36036 14318
rect 35980 12290 36036 14252
rect 36092 13970 36148 14700
rect 36092 13918 36094 13970
rect 36146 13918 36148 13970
rect 36092 13906 36148 13918
rect 36204 14306 36260 14924
rect 36204 14254 36206 14306
rect 36258 14254 36260 14306
rect 36204 13524 36260 14254
rect 36204 13458 36260 13468
rect 35980 12238 35982 12290
rect 36034 12238 36036 12290
rect 35980 12226 36036 12238
rect 36092 12740 36148 12750
rect 35980 11508 36036 11518
rect 36092 11508 36148 12684
rect 35980 11506 36148 11508
rect 35980 11454 35982 11506
rect 36034 11454 36148 11506
rect 35980 11452 36148 11454
rect 35980 11442 36036 11452
rect 36316 8428 36372 15092
rect 36428 15092 36484 15102
rect 36428 14998 36484 15036
rect 36428 13634 36484 13646
rect 36428 13582 36430 13634
rect 36482 13582 36484 13634
rect 36428 13524 36484 13582
rect 36428 13458 36484 13468
rect 36540 12516 36596 16604
rect 36764 14980 36820 18172
rect 37212 17108 37268 18620
rect 37324 18564 37380 18956
rect 37548 18788 37604 21310
rect 37660 20580 37716 20590
rect 37660 20486 37716 20524
rect 37660 19124 37716 19134
rect 37660 19030 37716 19068
rect 37324 18470 37380 18508
rect 37436 18732 37604 18788
rect 37436 17780 37492 18732
rect 37660 18564 37716 18574
rect 37548 18452 37604 18462
rect 37548 18358 37604 18396
rect 37436 17714 37492 17724
rect 37548 17442 37604 17454
rect 37548 17390 37550 17442
rect 37602 17390 37604 17442
rect 37436 17220 37492 17230
rect 37324 17108 37380 17118
rect 37212 17106 37380 17108
rect 37212 17054 37326 17106
rect 37378 17054 37380 17106
rect 37212 17052 37380 17054
rect 37324 17042 37380 17052
rect 37436 16322 37492 17164
rect 37436 16270 37438 16322
rect 37490 16270 37492 16322
rect 37436 16258 37492 16270
rect 37436 15874 37492 15886
rect 37436 15822 37438 15874
rect 37490 15822 37492 15874
rect 37436 15652 37492 15822
rect 37436 15586 37492 15596
rect 36988 15426 37044 15438
rect 36988 15374 36990 15426
rect 37042 15374 37044 15426
rect 36876 15316 36932 15326
rect 36876 15222 36932 15260
rect 36988 14980 37044 15374
rect 36764 14924 36932 14980
rect 36764 14756 36820 14766
rect 36764 14642 36820 14700
rect 36764 14590 36766 14642
rect 36818 14590 36820 14642
rect 36652 12740 36708 12750
rect 36652 12646 36708 12684
rect 36540 12460 36708 12516
rect 36540 11508 36596 11518
rect 36540 11414 36596 11452
rect 36540 11284 36596 11294
rect 36540 9154 36596 11228
rect 36540 9102 36542 9154
rect 36594 9102 36596 9154
rect 36540 9090 36596 9102
rect 34412 8372 34580 8428
rect 35756 8372 35924 8428
rect 36204 8372 36372 8428
rect 34412 4676 34468 8372
rect 35644 7474 35700 7486
rect 35644 7422 35646 7474
rect 35698 7422 35700 7474
rect 35196 7364 35252 7374
rect 35644 7364 35700 7422
rect 35196 7362 35700 7364
rect 35196 7310 35198 7362
rect 35250 7310 35700 7362
rect 35196 7308 35700 7310
rect 34860 5796 34916 5806
rect 35196 5796 35252 7308
rect 35420 5906 35476 5918
rect 35420 5854 35422 5906
rect 35474 5854 35476 5906
rect 35420 5796 35476 5854
rect 34860 5794 35476 5796
rect 34860 5742 34862 5794
rect 34914 5742 35476 5794
rect 34860 5740 35476 5742
rect 34636 5010 34692 5022
rect 34636 4958 34638 5010
rect 34690 4958 34692 5010
rect 34636 4900 34692 4958
rect 34636 4834 34692 4844
rect 34860 5012 34916 5740
rect 34412 4610 34468 4620
rect 34188 4498 34244 4508
rect 34076 4274 34132 4284
rect 34636 4340 34692 4350
rect 34860 4340 34916 4956
rect 35756 4452 35812 8372
rect 36204 6580 36260 8372
rect 36428 7700 36484 7710
rect 36428 7586 36484 7644
rect 36428 7534 36430 7586
rect 36482 7534 36484 7586
rect 36428 7522 36484 7534
rect 36204 6514 36260 6524
rect 36204 6132 36260 6142
rect 36204 6018 36260 6076
rect 36204 5966 36206 6018
rect 36258 5966 36260 6018
rect 36204 5954 36260 5966
rect 36652 5908 36708 12460
rect 36764 10498 36820 14590
rect 36876 10612 36932 14924
rect 36988 14644 37044 14924
rect 36988 14578 37044 14588
rect 37324 14756 37380 14766
rect 37324 13858 37380 14700
rect 37324 13806 37326 13858
rect 37378 13806 37380 13858
rect 37324 13794 37380 13806
rect 37548 12964 37604 17390
rect 37660 16658 37716 18508
rect 37772 17108 37828 22876
rect 37996 22866 38052 22876
rect 38332 22932 38388 23436
rect 39004 23492 39060 23774
rect 39004 23426 39060 23436
rect 39004 23268 39060 23278
rect 39004 23174 39060 23212
rect 39116 23154 39172 23884
rect 39676 23492 39732 23998
rect 40236 23996 40404 24052
rect 40796 25282 40852 26796
rect 40796 25230 40798 25282
rect 40850 25230 40852 25282
rect 40236 23604 40292 23996
rect 40796 23940 40852 25230
rect 41132 25284 41188 38668
rect 41776 37660 42352 37670
rect 41832 37604 41880 37660
rect 41936 37604 41984 37660
rect 42040 37604 42088 37660
rect 42144 37604 42192 37660
rect 42248 37604 42296 37660
rect 41776 37594 42352 37604
rect 44156 36260 44212 45612
rect 46172 45444 46228 45836
rect 46844 45826 46900 45836
rect 45836 45388 46228 45444
rect 47740 45778 47796 45790
rect 47740 45726 47742 45778
rect 47794 45726 47796 45778
rect 45836 45330 45892 45388
rect 45836 45278 45838 45330
rect 45890 45278 45892 45330
rect 44156 36194 44212 36204
rect 45612 37156 45668 37166
rect 41776 36092 42352 36102
rect 41832 36036 41880 36092
rect 41936 36036 41984 36092
rect 42040 36036 42088 36092
rect 42144 36036 42192 36092
rect 42248 36036 42296 36092
rect 41776 36026 42352 36036
rect 41776 34524 42352 34534
rect 41832 34468 41880 34524
rect 41936 34468 41984 34524
rect 42040 34468 42088 34524
rect 42144 34468 42192 34524
rect 42248 34468 42296 34524
rect 41776 34458 42352 34468
rect 41776 32956 42352 32966
rect 41832 32900 41880 32956
rect 41936 32900 41984 32956
rect 42040 32900 42088 32956
rect 42144 32900 42192 32956
rect 42248 32900 42296 32956
rect 41776 32890 42352 32900
rect 44492 32452 44548 32462
rect 41776 31388 42352 31398
rect 41832 31332 41880 31388
rect 41936 31332 41984 31388
rect 42040 31332 42088 31388
rect 42144 31332 42192 31388
rect 42248 31332 42296 31388
rect 41776 31322 42352 31332
rect 41776 29820 42352 29830
rect 41832 29764 41880 29820
rect 41936 29764 41984 29820
rect 42040 29764 42088 29820
rect 42144 29764 42192 29820
rect 42248 29764 42296 29820
rect 41776 29754 42352 29764
rect 41132 25218 41188 25228
rect 41244 29316 41300 29326
rect 40684 23938 40852 23940
rect 40684 23886 40798 23938
rect 40850 23886 40852 23938
rect 40684 23884 40852 23886
rect 40348 23826 40404 23838
rect 40348 23774 40350 23826
rect 40402 23774 40404 23826
rect 40348 23716 40404 23774
rect 40348 23660 40516 23716
rect 40236 23548 40404 23604
rect 39676 23426 39732 23436
rect 39116 23102 39118 23154
rect 39170 23102 39172 23154
rect 39116 23090 39172 23102
rect 38332 22866 38388 22876
rect 38056 22764 38632 22774
rect 38112 22708 38160 22764
rect 38216 22708 38264 22764
rect 38320 22708 38368 22764
rect 38424 22708 38472 22764
rect 38528 22708 38576 22764
rect 38056 22698 38632 22708
rect 38108 22260 38164 22270
rect 38108 22166 38164 22204
rect 38668 22260 38724 22270
rect 38668 22166 38724 22204
rect 38220 22146 38276 22158
rect 38220 22094 38222 22146
rect 38274 22094 38276 22146
rect 37884 21364 37940 21374
rect 37884 21270 37940 21308
rect 38220 21364 38276 22094
rect 38444 21698 38500 21710
rect 38444 21646 38446 21698
rect 38498 21646 38500 21698
rect 38444 21476 38500 21646
rect 38668 21588 38724 21598
rect 40348 21588 40404 23548
rect 38724 21532 38836 21588
rect 38668 21494 38724 21532
rect 38444 21410 38500 21420
rect 38220 21298 38276 21308
rect 38056 21196 38632 21206
rect 38112 21140 38160 21196
rect 38216 21140 38264 21196
rect 38320 21140 38368 21196
rect 38424 21140 38472 21196
rect 38528 21140 38576 21196
rect 38056 21130 38632 21140
rect 37996 21028 38052 21038
rect 37996 20934 38052 20972
rect 38332 21028 38388 21038
rect 38332 20244 38388 20972
rect 38668 21028 38724 21038
rect 38668 20690 38724 20972
rect 38668 20638 38670 20690
rect 38722 20638 38724 20690
rect 38668 20626 38724 20638
rect 38780 20802 38836 21532
rect 40348 21522 40404 21532
rect 38780 20750 38782 20802
rect 38834 20750 38836 20802
rect 38332 20178 38388 20188
rect 37996 20132 38052 20142
rect 37884 20076 37996 20132
rect 37884 19460 37940 20076
rect 37996 20000 38052 20076
rect 38220 20020 38276 20030
rect 38220 19926 38276 19964
rect 38780 20020 38836 20750
rect 39900 21364 39956 21374
rect 39452 20692 39508 20702
rect 39452 20598 39508 20636
rect 39900 20690 39956 21308
rect 40460 20916 40516 23660
rect 40348 20860 40516 20916
rect 39900 20638 39902 20690
rect 39954 20638 39956 20690
rect 39900 20626 39956 20638
rect 40012 20692 40068 20702
rect 40012 20598 40068 20636
rect 38056 19628 38632 19638
rect 38112 19572 38160 19628
rect 38216 19572 38264 19628
rect 38320 19572 38368 19628
rect 38424 19572 38472 19628
rect 38528 19572 38576 19628
rect 38056 19562 38632 19572
rect 37996 19460 38052 19470
rect 38780 19460 38836 19964
rect 39116 20580 39172 20590
rect 39116 19908 39172 20524
rect 39676 20580 39732 20590
rect 39676 20486 39732 20524
rect 37884 19404 37996 19460
rect 37996 19366 38052 19404
rect 38668 19404 38836 19460
rect 39004 19906 39172 19908
rect 39004 19854 39118 19906
rect 39170 19854 39172 19906
rect 39004 19852 39172 19854
rect 38668 19234 38724 19404
rect 38668 19182 38670 19234
rect 38722 19182 38724 19234
rect 38668 19170 38724 19182
rect 38780 19124 38836 19134
rect 38108 18788 38164 18798
rect 38108 18450 38164 18732
rect 38780 18788 38836 19068
rect 38780 18722 38836 18732
rect 38108 18398 38110 18450
rect 38162 18398 38164 18450
rect 38108 18386 38164 18398
rect 38556 18452 38612 18462
rect 38556 18358 38612 18396
rect 38780 18452 38836 18462
rect 38056 18060 38632 18070
rect 38112 18004 38160 18060
rect 38216 18004 38264 18060
rect 38320 18004 38368 18060
rect 38424 18004 38472 18060
rect 38528 18004 38576 18060
rect 38056 17994 38632 18004
rect 38780 17892 38836 18396
rect 38332 17836 38836 17892
rect 38332 17778 38388 17836
rect 38332 17726 38334 17778
rect 38386 17726 38388 17778
rect 37884 17556 37940 17566
rect 37884 17462 37940 17500
rect 37772 17042 37828 17052
rect 38220 17220 38276 17230
rect 38220 16994 38276 17164
rect 38220 16942 38222 16994
rect 38274 16942 38276 16994
rect 38220 16930 38276 16942
rect 38332 16882 38388 17726
rect 38332 16830 38334 16882
rect 38386 16830 38388 16882
rect 38332 16660 38388 16830
rect 37660 16606 37662 16658
rect 37714 16606 37716 16658
rect 37660 15652 37716 16606
rect 37884 16604 38388 16660
rect 37884 16212 37940 16604
rect 38056 16492 38632 16502
rect 38112 16436 38160 16492
rect 38216 16436 38264 16492
rect 38320 16436 38368 16492
rect 38424 16436 38472 16492
rect 38528 16436 38576 16492
rect 38056 16426 38632 16436
rect 38332 16322 38388 16334
rect 38332 16270 38334 16322
rect 38386 16270 38388 16322
rect 37996 16212 38052 16222
rect 37884 16210 38052 16212
rect 37884 16158 37998 16210
rect 38050 16158 38052 16210
rect 37884 16156 38052 16158
rect 37996 16146 38052 16156
rect 38332 16210 38388 16270
rect 38332 16158 38334 16210
rect 38386 16158 38388 16210
rect 38332 16146 38388 16158
rect 38780 16212 38836 17836
rect 39004 16884 39060 19852
rect 39116 19842 39172 19852
rect 40348 18452 40404 20860
rect 40684 20804 40740 23884
rect 40796 23874 40852 23884
rect 40460 20748 40740 20804
rect 40460 20690 40516 20748
rect 40460 20638 40462 20690
rect 40514 20638 40516 20690
rect 40460 20626 40516 20638
rect 40796 20692 40852 20702
rect 40796 20598 40852 20636
rect 41244 19012 41300 29260
rect 41776 28252 42352 28262
rect 41832 28196 41880 28252
rect 41936 28196 41984 28252
rect 42040 28196 42088 28252
rect 42144 28196 42192 28252
rect 42248 28196 42296 28252
rect 41776 28186 42352 28196
rect 42812 26964 42868 26974
rect 41776 26684 42352 26694
rect 41832 26628 41880 26684
rect 41936 26628 41984 26684
rect 42040 26628 42088 26684
rect 42144 26628 42192 26684
rect 42248 26628 42296 26684
rect 41776 26618 42352 26628
rect 41776 25116 42352 25126
rect 41832 25060 41880 25116
rect 41936 25060 41984 25116
rect 42040 25060 42088 25116
rect 42144 25060 42192 25116
rect 42248 25060 42296 25116
rect 41776 25050 42352 25060
rect 41776 23548 42352 23558
rect 41832 23492 41880 23548
rect 41936 23492 41984 23548
rect 42040 23492 42088 23548
rect 42144 23492 42192 23548
rect 42248 23492 42296 23548
rect 41776 23482 42352 23492
rect 41776 21980 42352 21990
rect 41832 21924 41880 21980
rect 41936 21924 41984 21980
rect 42040 21924 42088 21980
rect 42144 21924 42192 21980
rect 42248 21924 42296 21980
rect 41776 21914 42352 21924
rect 41244 18946 41300 18956
rect 41580 20692 41636 20702
rect 40348 18386 40404 18396
rect 39116 17108 39172 17118
rect 39116 17106 39844 17108
rect 39116 17054 39118 17106
rect 39170 17054 39844 17106
rect 39116 17052 39844 17054
rect 39116 17042 39172 17052
rect 39004 16828 39284 16884
rect 38892 16212 38948 16222
rect 38780 16210 38948 16212
rect 38780 16158 38894 16210
rect 38946 16158 38948 16210
rect 38780 16156 38948 16158
rect 38892 16146 38948 16156
rect 37660 15586 37716 15596
rect 37884 15988 37940 15998
rect 37660 15092 37716 15102
rect 37660 14420 37716 15036
rect 37884 14756 37940 15932
rect 39116 15540 39172 15550
rect 39116 15446 39172 15484
rect 38220 15426 38276 15438
rect 38220 15374 38222 15426
rect 38274 15374 38276 15426
rect 37996 15314 38052 15326
rect 37996 15262 37998 15314
rect 38050 15262 38052 15314
rect 37996 15092 38052 15262
rect 38220 15204 38276 15374
rect 38892 15428 38948 15438
rect 38220 15138 38276 15148
rect 38780 15314 38836 15326
rect 38780 15262 38782 15314
rect 38834 15262 38836 15314
rect 37996 15026 38052 15036
rect 38780 15092 38836 15262
rect 38780 15026 38836 15036
rect 38056 14924 38632 14934
rect 38112 14868 38160 14924
rect 38216 14868 38264 14924
rect 38320 14868 38368 14924
rect 38424 14868 38472 14924
rect 38528 14868 38576 14924
rect 38056 14858 38632 14868
rect 38780 14756 38836 14766
rect 38892 14756 38948 15372
rect 37884 14700 38276 14756
rect 37660 13858 37716 14364
rect 37660 13806 37662 13858
rect 37714 13806 37716 13858
rect 37660 13794 37716 13806
rect 37884 14418 37940 14430
rect 37884 14366 37886 14418
rect 37938 14366 37940 14418
rect 37884 14196 37940 14366
rect 38108 14420 38164 14430
rect 38108 14326 38164 14364
rect 36876 10546 36932 10556
rect 37100 12908 37604 12964
rect 37884 13746 37940 14140
rect 38220 13970 38276 14700
rect 38780 14754 38948 14756
rect 38780 14702 38782 14754
rect 38834 14702 38948 14754
rect 38780 14700 38948 14702
rect 38780 14690 38836 14700
rect 38444 14644 38500 14654
rect 38444 14550 38500 14588
rect 38220 13918 38222 13970
rect 38274 13918 38276 13970
rect 38220 13906 38276 13918
rect 39004 13972 39060 13982
rect 39004 13878 39060 13916
rect 37884 13694 37886 13746
rect 37938 13694 37940 13746
rect 36764 10446 36766 10498
rect 36818 10446 36820 10498
rect 36764 10434 36820 10446
rect 36652 5842 36708 5852
rect 36764 6580 36820 6590
rect 36764 5234 36820 6524
rect 36764 5182 36766 5234
rect 36818 5182 36820 5234
rect 36764 5170 36820 5182
rect 35756 4386 35812 4396
rect 34692 4284 34916 4340
rect 34636 4246 34692 4284
rect 30044 3726 30046 3778
rect 30098 3726 30100 3778
rect 30044 3714 30100 3726
rect 35420 4226 35476 4238
rect 35420 4174 35422 4226
rect 35474 4174 35476 4226
rect 25676 3502 25678 3554
rect 25730 3502 25732 3554
rect 29260 3536 29316 3612
rect 30156 3668 30212 3678
rect 30156 3574 30212 3612
rect 35420 3668 35476 4174
rect 35420 3602 35476 3612
rect 25676 3490 25732 3502
rect 26348 3444 26404 3454
rect 26348 3350 26404 3388
rect 29708 3444 29764 3454
rect 29708 3350 29764 3388
rect 37100 3444 37156 12908
rect 37436 12740 37492 12750
rect 37884 12740 37940 13694
rect 38056 13356 38632 13366
rect 38112 13300 38160 13356
rect 38216 13300 38264 13356
rect 38320 13300 38368 13356
rect 38424 13300 38472 13356
rect 38528 13300 38576 13356
rect 38056 13290 38632 13300
rect 38556 13188 38612 13198
rect 38556 13076 38612 13132
rect 37492 12684 37940 12740
rect 38108 13074 38612 13076
rect 38108 13022 38558 13074
rect 38610 13022 38612 13074
rect 38108 13020 38612 13022
rect 37436 12608 37492 12684
rect 38108 12066 38164 13020
rect 38556 13010 38612 13020
rect 38108 12014 38110 12066
rect 38162 12014 38164 12066
rect 38108 12002 38164 12014
rect 38056 11788 38632 11798
rect 39228 11788 39284 16828
rect 39340 16882 39396 16894
rect 39340 16830 39342 16882
rect 39394 16830 39396 16882
rect 39340 15428 39396 16830
rect 39340 15362 39396 15372
rect 39452 16884 39508 16894
rect 39340 15204 39396 15214
rect 39340 13522 39396 15148
rect 39452 15092 39508 16828
rect 39452 15026 39508 15036
rect 39676 15874 39732 15886
rect 39676 15822 39678 15874
rect 39730 15822 39732 15874
rect 39676 14644 39732 15822
rect 39340 13470 39342 13522
rect 39394 13470 39396 13522
rect 39340 13188 39396 13470
rect 39340 13122 39396 13132
rect 39564 14588 39732 14644
rect 38112 11732 38160 11788
rect 38216 11732 38264 11788
rect 38320 11732 38368 11788
rect 38424 11732 38472 11788
rect 38528 11732 38576 11788
rect 38056 11722 38632 11732
rect 38892 11732 39284 11788
rect 38332 11620 38388 11630
rect 38332 11506 38388 11564
rect 38332 11454 38334 11506
rect 38386 11454 38388 11506
rect 38332 11442 38388 11454
rect 37212 11396 37268 11406
rect 37548 11396 37604 11406
rect 37268 11394 37604 11396
rect 37268 11342 37550 11394
rect 37602 11342 37604 11394
rect 37268 11340 37604 11342
rect 37212 10834 37268 11340
rect 37548 11330 37604 11340
rect 37660 11396 37716 11406
rect 37212 10782 37214 10834
rect 37266 10782 37268 10834
rect 37212 10770 37268 10782
rect 37660 10834 37716 11340
rect 37660 10782 37662 10834
rect 37714 10782 37716 10834
rect 37660 10724 37716 10782
rect 37660 10658 37716 10668
rect 38780 10500 38836 10510
rect 38056 10220 38632 10230
rect 38112 10164 38160 10220
rect 38216 10164 38264 10220
rect 38320 10164 38368 10220
rect 38424 10164 38472 10220
rect 38528 10164 38576 10220
rect 38056 10154 38632 10164
rect 37548 9604 37604 9614
rect 37548 6802 37604 9548
rect 38668 8932 38724 8942
rect 38780 8932 38836 10444
rect 38668 8930 38836 8932
rect 38668 8878 38670 8930
rect 38722 8878 38836 8930
rect 38668 8876 38836 8878
rect 38668 8866 38724 8876
rect 38056 8652 38632 8662
rect 38112 8596 38160 8652
rect 38216 8596 38264 8652
rect 38320 8596 38368 8652
rect 38424 8596 38472 8652
rect 38528 8596 38576 8652
rect 38056 8586 38632 8596
rect 38556 8484 38612 8494
rect 38556 7362 38612 8428
rect 38892 8148 38948 11732
rect 39564 11508 39620 14588
rect 39676 14308 39732 14318
rect 39676 14214 39732 14252
rect 39564 11442 39620 11452
rect 39788 9380 39844 17052
rect 41580 16994 41636 20636
rect 41776 20412 42352 20422
rect 41832 20356 41880 20412
rect 41936 20356 41984 20412
rect 42040 20356 42088 20412
rect 42144 20356 42192 20412
rect 42248 20356 42296 20412
rect 41776 20346 42352 20356
rect 41776 18844 42352 18854
rect 41832 18788 41880 18844
rect 41936 18788 41984 18844
rect 42040 18788 42088 18844
rect 42144 18788 42192 18844
rect 42248 18788 42296 18844
rect 41776 18778 42352 18788
rect 42812 17668 42868 26908
rect 44492 20132 44548 32396
rect 45500 31108 45556 31118
rect 45500 24836 45556 31052
rect 45500 24770 45556 24780
rect 45612 23268 45668 37100
rect 45612 23202 45668 23212
rect 45724 28644 45780 28654
rect 44492 20066 44548 20076
rect 42812 17602 42868 17612
rect 41776 17276 42352 17286
rect 41832 17220 41880 17276
rect 41936 17220 41984 17276
rect 42040 17220 42088 17276
rect 42144 17220 42192 17276
rect 42248 17220 42296 17276
rect 41776 17210 42352 17220
rect 45724 17108 45780 28588
rect 45836 27972 45892 45278
rect 47740 45332 47796 45726
rect 47740 45266 47796 45276
rect 46844 45108 46900 45118
rect 46396 45106 46900 45108
rect 46396 45054 46846 45106
rect 46898 45054 46900 45106
rect 46396 45052 46900 45054
rect 46396 44994 46452 45052
rect 46844 45042 46900 45052
rect 46396 44942 46398 44994
rect 46450 44942 46452 44994
rect 46396 44548 46452 44942
rect 47852 44994 47908 46732
rect 47852 44942 47854 44994
rect 47906 44942 47908 44994
rect 47852 44930 47908 44942
rect 45948 44492 46452 44548
rect 45948 28084 46004 44492
rect 46284 44324 46340 44334
rect 46844 44324 46900 44334
rect 46284 44322 46900 44324
rect 46284 44270 46286 44322
rect 46338 44270 46846 44322
rect 46898 44270 46900 44322
rect 46284 44268 46900 44270
rect 46284 43708 46340 44268
rect 46844 44258 46900 44268
rect 47740 44210 47796 44222
rect 47740 44158 47742 44210
rect 47794 44158 47796 44210
rect 47740 43876 47796 44158
rect 47740 43810 47796 43820
rect 46060 43652 46340 43708
rect 46060 29540 46116 43652
rect 46844 42754 46900 42766
rect 46844 42702 46846 42754
rect 46898 42702 46900 42754
rect 46284 42530 46340 42542
rect 46284 42478 46286 42530
rect 46338 42478 46340 42530
rect 46284 41972 46340 42478
rect 46284 41906 46340 41916
rect 46844 41972 46900 42702
rect 47740 42642 47796 42654
rect 47740 42590 47742 42642
rect 47794 42590 47796 42642
rect 47740 42420 47796 42590
rect 47740 42354 47796 42364
rect 46844 41906 46900 41916
rect 46844 41188 46900 41198
rect 46284 41186 46900 41188
rect 46284 41134 46846 41186
rect 46898 41134 46900 41186
rect 46284 41132 46900 41134
rect 46284 40964 46340 41132
rect 46844 41122 46900 41132
rect 46172 40962 46340 40964
rect 46172 40910 46286 40962
rect 46338 40910 46340 40962
rect 46172 40908 46340 40910
rect 46172 37940 46228 40908
rect 46284 40898 46340 40908
rect 47740 41074 47796 41086
rect 47740 41022 47742 41074
rect 47794 41022 47796 41074
rect 47740 40964 47796 41022
rect 47740 40898 47796 40908
rect 46844 39620 46900 39630
rect 46732 39618 46900 39620
rect 46732 39566 46846 39618
rect 46898 39566 46900 39618
rect 46732 39564 46900 39566
rect 46284 39396 46340 39406
rect 46732 39396 46788 39564
rect 46844 39554 46900 39564
rect 47740 39508 47796 39518
rect 47740 39414 47796 39452
rect 46284 39394 46788 39396
rect 46284 39342 46286 39394
rect 46338 39342 46788 39394
rect 46284 39340 46788 39342
rect 46284 39330 46340 39340
rect 46396 38724 46452 38734
rect 46396 38630 46452 38668
rect 46172 37884 46564 37940
rect 46396 37156 46452 37166
rect 46396 37062 46452 37100
rect 46396 35700 46452 35710
rect 46396 35606 46452 35644
rect 46396 34020 46452 34030
rect 46284 34018 46452 34020
rect 46284 33966 46398 34018
rect 46450 33966 46452 34018
rect 46284 33964 46452 33966
rect 46284 33906 46340 33964
rect 46396 33954 46452 33964
rect 46284 33854 46286 33906
rect 46338 33854 46340 33906
rect 46284 31948 46340 33854
rect 46396 32452 46452 32462
rect 46396 32358 46452 32396
rect 46060 29474 46116 29484
rect 46172 31892 46340 31948
rect 46508 31948 46564 37884
rect 46508 31892 46676 31948
rect 45948 28018 46004 28028
rect 45836 27906 45892 27916
rect 46172 26908 46228 31892
rect 46396 30994 46452 31006
rect 46396 30942 46398 30994
rect 46450 30942 46452 30994
rect 46396 30884 46452 30942
rect 46508 30884 46564 30894
rect 46396 30882 46564 30884
rect 46396 30830 46510 30882
rect 46562 30830 46564 30882
rect 46396 30828 46564 30830
rect 46508 30818 46564 30828
rect 46396 29316 46452 29326
rect 46396 29222 46452 29260
rect 46284 28644 46340 28654
rect 46284 28550 46340 28588
rect 46060 26852 46228 26908
rect 46284 26964 46340 26974
rect 46284 26870 46340 26908
rect 45836 25732 45892 25742
rect 45836 19124 45892 25676
rect 46060 21028 46116 26852
rect 46620 26404 46676 31892
rect 46732 31108 46788 39340
rect 46844 38834 46900 38846
rect 46844 38782 46846 38834
rect 46898 38782 46900 38834
rect 46844 38724 46900 38782
rect 46844 38658 46900 38668
rect 47852 38724 47908 38734
rect 47852 38630 47908 38668
rect 46844 37266 46900 37278
rect 46844 37214 46846 37266
rect 46898 37214 46900 37266
rect 46844 37156 46900 37214
rect 46844 37090 46900 37100
rect 47852 37154 47908 37166
rect 47852 37102 47854 37154
rect 47906 37102 47908 37154
rect 47852 36596 47908 37102
rect 47852 36530 47908 36540
rect 46956 35700 47012 35710
rect 47012 35644 47124 35700
rect 46956 35568 47012 35644
rect 46956 34130 47012 34142
rect 46956 34078 46958 34130
rect 47010 34078 47012 34130
rect 46844 34020 46900 34030
rect 46956 34020 47012 34078
rect 46844 34018 47012 34020
rect 46844 33966 46846 34018
rect 46898 33966 47012 34018
rect 46844 33964 47012 33966
rect 46844 33954 46900 33964
rect 46844 32562 46900 32574
rect 46844 32510 46846 32562
rect 46898 32510 46900 32562
rect 46844 32452 46900 32510
rect 46844 32386 46900 32396
rect 46732 31042 46788 31052
rect 46956 30994 47012 31006
rect 46956 30942 46958 30994
rect 47010 30942 47012 30994
rect 46844 30884 46900 30894
rect 46956 30884 47012 30942
rect 46844 30882 47012 30884
rect 46844 30830 46846 30882
rect 46898 30830 47012 30882
rect 46844 30828 47012 30830
rect 46844 30818 46900 30828
rect 46844 29426 46900 29438
rect 46844 29374 46846 29426
rect 46898 29374 46900 29426
rect 46844 29316 46900 29374
rect 46844 29250 46900 29260
rect 46844 28644 46900 28654
rect 46844 28550 46900 28588
rect 46844 27074 46900 27086
rect 46844 27022 46846 27074
rect 46898 27022 46900 27074
rect 46844 26964 46900 27022
rect 46844 26898 46900 26908
rect 46620 26338 46676 26348
rect 46956 25732 47012 30828
rect 46956 25666 47012 25676
rect 46956 25506 47012 25518
rect 46956 25454 46958 25506
rect 47010 25454 47012 25506
rect 46284 25284 46340 25294
rect 46956 25284 47012 25454
rect 46284 25282 47012 25284
rect 46284 25230 46286 25282
rect 46338 25230 47012 25282
rect 46284 25228 47012 25230
rect 46284 25218 46340 25228
rect 46844 23938 46900 23950
rect 46844 23886 46846 23938
rect 46898 23886 46900 23938
rect 46284 23716 46340 23726
rect 46844 23716 46900 23886
rect 46284 23714 46900 23716
rect 46284 23662 46286 23714
rect 46338 23662 46900 23714
rect 46284 23660 46900 23662
rect 46284 22372 46340 23660
rect 46060 20962 46116 20972
rect 46172 22316 46340 22372
rect 46844 22370 46900 22382
rect 46844 22318 46846 22370
rect 46898 22318 46900 22370
rect 46172 20804 46228 22316
rect 46284 22148 46340 22158
rect 46284 22054 46340 22092
rect 46844 22148 46900 22318
rect 46844 22082 46900 22092
rect 46844 20804 46900 20814
rect 45836 19058 45892 19068
rect 45948 20748 46228 20804
rect 46284 20802 46900 20804
rect 46284 20750 46846 20802
rect 46898 20750 46900 20802
rect 46284 20748 46900 20750
rect 45724 17042 45780 17052
rect 41580 16942 41582 16994
rect 41634 16942 41636 16994
rect 41580 16930 41636 16942
rect 41916 16994 41972 17006
rect 41916 16942 41918 16994
rect 41970 16942 41972 16994
rect 40796 16098 40852 16110
rect 40796 16046 40798 16098
rect 40850 16046 40852 16098
rect 40012 15988 40068 15998
rect 40012 15894 40068 15932
rect 40572 15876 40628 15886
rect 40348 15874 40628 15876
rect 40348 15822 40574 15874
rect 40626 15822 40628 15874
rect 40348 15820 40628 15822
rect 40012 15316 40068 15326
rect 40012 15222 40068 15260
rect 39900 14530 39956 14542
rect 39900 14478 39902 14530
rect 39954 14478 39956 14530
rect 39900 13972 39956 14478
rect 39900 13906 39956 13916
rect 40012 14420 40068 14430
rect 40012 13746 40068 14364
rect 40012 13694 40014 13746
rect 40066 13694 40068 13746
rect 40012 13682 40068 13694
rect 40124 13858 40180 13870
rect 40124 13806 40126 13858
rect 40178 13806 40180 13858
rect 40124 13748 40180 13806
rect 40124 13682 40180 13692
rect 40348 12964 40404 15820
rect 40572 15810 40628 15820
rect 40796 15540 40852 16046
rect 41916 15876 41972 16942
rect 45948 16100 46004 20748
rect 46284 20580 46340 20748
rect 46844 20738 46900 20748
rect 46060 20578 46340 20580
rect 46060 20526 46286 20578
rect 46338 20526 46340 20578
rect 46060 20524 46340 20526
rect 46060 17444 46116 20524
rect 46284 20514 46340 20524
rect 46844 19236 46900 19246
rect 46284 19234 46900 19236
rect 46284 19182 46846 19234
rect 46898 19182 46900 19234
rect 46284 19180 46900 19182
rect 46284 19012 46340 19180
rect 46844 19170 46900 19180
rect 46060 17378 46116 17388
rect 46172 19010 46340 19012
rect 46172 18958 46286 19010
rect 46338 18958 46340 19010
rect 46172 18956 46340 18958
rect 45948 16034 46004 16044
rect 40796 15474 40852 15484
rect 41356 15820 41972 15876
rect 40572 15314 40628 15326
rect 40572 15262 40574 15314
rect 40626 15262 40628 15314
rect 40572 15148 40628 15262
rect 41356 15148 41412 15820
rect 41776 15708 42352 15718
rect 41832 15652 41880 15708
rect 41936 15652 41984 15708
rect 42040 15652 42088 15708
rect 42144 15652 42192 15708
rect 42248 15652 42296 15708
rect 41776 15642 42352 15652
rect 41468 15316 41524 15326
rect 41468 15222 41524 15260
rect 40572 15092 41412 15148
rect 40572 14420 40628 14430
rect 40572 14326 40628 14364
rect 41132 14306 41188 15092
rect 46172 14644 46228 18956
rect 46284 18946 46340 18956
rect 46844 18452 46900 18462
rect 46508 18450 46900 18452
rect 46508 18398 46846 18450
rect 46898 18398 46900 18450
rect 46508 18396 46900 18398
rect 46396 18340 46452 18350
rect 46508 18340 46564 18396
rect 46844 18386 46900 18396
rect 46396 18338 46564 18340
rect 46396 18286 46398 18338
rect 46450 18286 46564 18338
rect 46396 18284 46564 18286
rect 46396 18274 46452 18284
rect 46396 16884 46452 16894
rect 46396 16790 46452 16828
rect 46284 15316 46340 15326
rect 46284 15222 46340 15260
rect 46172 14578 46228 14588
rect 41132 14254 41134 14306
rect 41186 14254 41188 14306
rect 40684 13748 40740 13758
rect 40684 13654 40740 13692
rect 41132 12964 41188 14254
rect 46508 14308 46564 18284
rect 46956 16996 47012 25228
rect 47068 20916 47124 35644
rect 47852 35586 47908 35598
rect 47852 35534 47854 35586
rect 47906 35534 47908 35586
rect 47852 35364 47908 35534
rect 47852 35298 47908 35308
rect 47852 34018 47908 34030
rect 47852 33966 47854 34018
rect 47906 33966 47908 34018
rect 47852 33684 47908 33966
rect 47852 33618 47908 33628
rect 47852 32450 47908 32462
rect 47852 32398 47854 32450
rect 47906 32398 47908 32450
rect 47852 32228 47908 32398
rect 47852 32162 47908 32172
rect 47852 30882 47908 30894
rect 47852 30830 47854 30882
rect 47906 30830 47908 30882
rect 47852 30772 47908 30830
rect 47852 30706 47908 30716
rect 47852 29316 47908 29326
rect 47852 29222 47908 29260
rect 47852 28754 47908 28766
rect 47852 28702 47854 28754
rect 47906 28702 47908 28754
rect 47852 27860 47908 28702
rect 47852 27794 47908 27804
rect 47740 26962 47796 26974
rect 47740 26910 47742 26962
rect 47794 26910 47796 26962
rect 47740 26404 47796 26910
rect 47740 26338 47796 26348
rect 47740 25394 47796 25406
rect 47740 25342 47742 25394
rect 47794 25342 47796 25394
rect 47740 24948 47796 25342
rect 47740 24882 47796 24892
rect 47740 23826 47796 23838
rect 47740 23774 47742 23826
rect 47794 23774 47796 23826
rect 47740 23492 47796 23774
rect 47740 23426 47796 23436
rect 47740 22258 47796 22270
rect 47740 22206 47742 22258
rect 47794 22206 47796 22258
rect 47740 22036 47796 22206
rect 47740 21970 47796 21980
rect 47068 20850 47124 20860
rect 47740 20690 47796 20702
rect 47740 20638 47742 20690
rect 47794 20638 47796 20690
rect 47740 20580 47796 20638
rect 47740 20514 47796 20524
rect 47740 19124 47796 19134
rect 47740 19030 47796 19068
rect 47852 18338 47908 18350
rect 47852 18286 47854 18338
rect 47906 18286 47908 18338
rect 47852 17668 47908 18286
rect 47852 17602 47908 17612
rect 46956 16930 47012 16940
rect 46844 16884 46900 16894
rect 46844 16790 46900 16828
rect 47740 16884 47796 16894
rect 47740 16790 47796 16828
rect 46844 15316 46900 15326
rect 46844 15222 46900 15260
rect 47852 15202 47908 15214
rect 47852 15150 47854 15202
rect 47906 15150 47908 15202
rect 47852 14756 47908 15150
rect 47852 14690 47908 14700
rect 46508 14242 46564 14252
rect 41776 14140 42352 14150
rect 41832 14084 41880 14140
rect 41936 14084 41984 14140
rect 42040 14084 42088 14140
rect 42144 14084 42192 14140
rect 42248 14084 42296 14140
rect 41776 14074 42352 14084
rect 42476 13748 42532 13758
rect 41468 12964 41524 12974
rect 40348 12908 40740 12964
rect 41132 12962 41524 12964
rect 41132 12910 41470 12962
rect 41522 12910 41524 12962
rect 41132 12908 41524 12910
rect 40460 12740 40516 12750
rect 40348 12738 40516 12740
rect 40348 12686 40462 12738
rect 40514 12686 40516 12738
rect 40348 12684 40516 12686
rect 40348 11844 40404 12684
rect 40460 12674 40516 12684
rect 40460 12292 40516 12302
rect 40460 12290 40628 12292
rect 40460 12238 40462 12290
rect 40514 12238 40628 12290
rect 40460 12236 40628 12238
rect 40460 12226 40516 12236
rect 40348 11778 40404 11788
rect 40460 11732 40516 11742
rect 40460 11506 40516 11676
rect 40460 11454 40462 11506
rect 40514 11454 40516 11506
rect 40460 11442 40516 11454
rect 40572 11284 40628 12236
rect 40684 11396 40740 12908
rect 40796 12850 40852 12862
rect 40796 12798 40798 12850
rect 40850 12798 40852 12850
rect 40796 12404 40852 12798
rect 40796 12338 40852 12348
rect 41468 12292 41524 12908
rect 41916 12852 41972 12862
rect 41916 12758 41972 12796
rect 41776 12572 42352 12582
rect 41832 12516 41880 12572
rect 41936 12516 41984 12572
rect 42040 12516 42088 12572
rect 42144 12516 42192 12572
rect 42248 12516 42296 12572
rect 41776 12506 42352 12516
rect 42476 12404 42532 13692
rect 46284 13748 46340 13758
rect 46284 13654 46340 13692
rect 46844 13748 46900 13758
rect 46844 13654 46900 13692
rect 47852 13634 47908 13646
rect 47852 13582 47854 13634
rect 47906 13582 47908 13634
rect 47852 13524 47908 13582
rect 47852 13458 47908 13468
rect 42028 12348 42532 12404
rect 42700 12852 42756 12862
rect 41468 12236 41860 12292
rect 40796 12180 40852 12190
rect 40796 12178 41636 12180
rect 40796 12126 40798 12178
rect 40850 12126 41636 12178
rect 40796 12124 41636 12126
rect 40796 12114 40852 12124
rect 41132 11844 41188 11854
rect 41132 11506 41188 11788
rect 41132 11454 41134 11506
rect 41186 11454 41188 11506
rect 41132 11442 41188 11454
rect 40684 11330 40740 11340
rect 40572 11218 40628 11228
rect 41468 11284 41524 11294
rect 40796 10500 40852 10510
rect 40796 10406 40852 10444
rect 41244 9604 41300 9614
rect 39788 9314 39844 9324
rect 41132 9602 41300 9604
rect 41132 9550 41246 9602
rect 41298 9550 41300 9602
rect 41132 9548 41300 9550
rect 41132 8484 41188 9548
rect 41244 9538 41300 9548
rect 41132 8370 41188 8428
rect 41132 8318 41134 8370
rect 41186 8318 41188 8370
rect 41132 8306 41188 8318
rect 38892 8082 38948 8092
rect 40684 8148 40740 8158
rect 39004 7700 39060 7710
rect 40684 7700 40740 8092
rect 40796 7700 40852 7710
rect 41468 7700 41524 11228
rect 41580 10836 41636 12124
rect 41692 12068 41748 12078
rect 41692 11974 41748 12012
rect 41804 11394 41860 12236
rect 42028 12178 42084 12348
rect 42588 12292 42644 12302
rect 42028 12126 42030 12178
rect 42082 12126 42084 12178
rect 42028 11844 42084 12126
rect 42028 11778 42084 11788
rect 42476 12236 42588 12292
rect 41804 11342 41806 11394
rect 41858 11342 41860 11394
rect 41804 11330 41860 11342
rect 42364 11284 42420 11294
rect 42364 11190 42420 11228
rect 41776 11004 42352 11014
rect 41832 10948 41880 11004
rect 41936 10948 41984 11004
rect 42040 10948 42088 11004
rect 42144 10948 42192 11004
rect 42248 10948 42296 11004
rect 41776 10938 42352 10948
rect 41692 10836 41748 10846
rect 41580 10834 41748 10836
rect 41580 10782 41694 10834
rect 41746 10782 41748 10834
rect 41580 10780 41748 10782
rect 41692 10770 41748 10780
rect 42028 10500 42084 10510
rect 42028 10406 42084 10444
rect 42476 10500 42532 12236
rect 42588 12160 42644 12236
rect 42700 12178 42756 12796
rect 43372 12292 43428 12302
rect 43372 12198 43428 12236
rect 46284 12292 46340 12302
rect 46284 12198 46340 12236
rect 46844 12292 46900 12302
rect 42700 12126 42702 12178
rect 42754 12126 42756 12178
rect 42476 10434 42532 10444
rect 42588 10722 42644 10734
rect 42588 10670 42590 10722
rect 42642 10670 42644 10722
rect 42588 10052 42644 10670
rect 42476 9714 42532 9726
rect 42476 9662 42478 9714
rect 42530 9662 42532 9714
rect 42140 9604 42196 9642
rect 42140 9538 42196 9548
rect 41776 9436 42352 9446
rect 41832 9380 41880 9436
rect 41936 9380 41984 9436
rect 42040 9380 42088 9436
rect 42144 9380 42192 9436
rect 42248 9380 42296 9436
rect 41776 9370 42352 9380
rect 40684 7698 40852 7700
rect 40684 7646 40798 7698
rect 40850 7646 40852 7698
rect 40684 7644 40852 7646
rect 39004 7606 39060 7644
rect 38556 7310 38558 7362
rect 38610 7310 38612 7362
rect 38556 7298 38612 7310
rect 38056 7084 38632 7094
rect 38112 7028 38160 7084
rect 38216 7028 38264 7084
rect 38320 7028 38368 7084
rect 38424 7028 38472 7084
rect 38528 7028 38576 7084
rect 38056 7018 38632 7028
rect 37548 6750 37550 6802
rect 37602 6750 37604 6802
rect 37548 6132 37604 6750
rect 38332 6804 38388 6814
rect 38108 6580 38164 6590
rect 38108 6486 38164 6524
rect 37548 6066 37604 6076
rect 37660 6356 37716 6366
rect 37548 5122 37604 5134
rect 37548 5070 37550 5122
rect 37602 5070 37604 5122
rect 37324 5012 37380 5022
rect 37324 3666 37380 4956
rect 37548 5012 37604 5070
rect 37548 4946 37604 4956
rect 37548 4228 37604 4238
rect 37660 4228 37716 6300
rect 38332 5794 38388 6748
rect 40796 6804 40852 7644
rect 40796 6738 40852 6748
rect 41356 7698 41524 7700
rect 41356 7646 41470 7698
rect 41522 7646 41524 7698
rect 41356 7644 41524 7646
rect 40348 6690 40404 6702
rect 40348 6638 40350 6690
rect 40402 6638 40404 6690
rect 38556 6580 38612 6590
rect 38556 6486 38612 6524
rect 39788 6580 39844 6590
rect 40124 6580 40180 6590
rect 39844 6524 39956 6580
rect 38892 6466 38948 6478
rect 38892 6414 38894 6466
rect 38946 6414 38948 6466
rect 38892 6356 38948 6414
rect 38892 6132 38948 6300
rect 38892 6066 38948 6076
rect 39676 6468 39732 6478
rect 39788 6448 39844 6524
rect 38332 5742 38334 5794
rect 38386 5742 38388 5794
rect 38332 5730 38388 5742
rect 39340 6018 39396 6030
rect 39340 5966 39342 6018
rect 39394 5966 39396 6018
rect 38056 5516 38632 5526
rect 38112 5460 38160 5516
rect 38216 5460 38264 5516
rect 38320 5460 38368 5516
rect 38424 5460 38472 5516
rect 38528 5460 38576 5516
rect 38056 5450 38632 5460
rect 38332 5236 38388 5246
rect 38332 5142 38388 5180
rect 38108 5012 38164 5022
rect 38108 4562 38164 4956
rect 38892 5012 38948 5022
rect 38108 4510 38110 4562
rect 38162 4510 38164 4562
rect 38108 4498 38164 4510
rect 38444 4564 38500 4574
rect 38444 4470 38500 4508
rect 38892 4562 38948 4956
rect 38892 4510 38894 4562
rect 38946 4510 38948 4562
rect 38892 4498 38948 4510
rect 39340 4788 39396 5966
rect 39676 6018 39732 6412
rect 39676 5966 39678 6018
rect 39730 5966 39732 6018
rect 39676 5954 39732 5966
rect 39900 5684 39956 6524
rect 40124 6486 40180 6524
rect 40348 6132 40404 6638
rect 40684 6692 40740 6702
rect 40684 6598 40740 6636
rect 41356 6580 41412 7644
rect 41468 7634 41524 7644
rect 41580 8260 41636 8270
rect 41580 6690 41636 8204
rect 42028 8260 42084 8270
rect 42028 8166 42084 8204
rect 41916 8148 41972 8158
rect 41916 8054 41972 8092
rect 41776 7868 42352 7878
rect 41832 7812 41880 7868
rect 41936 7812 41984 7868
rect 42040 7812 42088 7868
rect 42144 7812 42192 7868
rect 42248 7812 42296 7868
rect 41776 7802 42352 7812
rect 41580 6638 41582 6690
rect 41634 6638 41636 6690
rect 41580 6626 41636 6638
rect 41916 7362 41972 7374
rect 41916 7310 41918 7362
rect 41970 7310 41972 7362
rect 40348 6066 40404 6076
rect 41244 6132 41300 6142
rect 40796 5794 40852 5806
rect 40796 5742 40798 5794
rect 40850 5742 40852 5794
rect 39900 5590 39956 5628
rect 40236 5682 40292 5694
rect 40236 5630 40238 5682
rect 40290 5630 40292 5682
rect 40236 5012 40292 5630
rect 40684 5460 40740 5470
rect 40460 5348 40516 5358
rect 40460 5234 40516 5292
rect 40460 5182 40462 5234
rect 40514 5182 40516 5234
rect 40460 5170 40516 5182
rect 40236 4946 40292 4956
rect 39340 4452 39396 4732
rect 40684 4562 40740 5404
rect 40684 4510 40686 4562
rect 40738 4510 40740 4562
rect 40684 4498 40740 4510
rect 39340 4386 39396 4396
rect 40124 4452 40180 4462
rect 40124 4358 40180 4396
rect 40796 4452 40852 5742
rect 41244 4452 41300 6076
rect 41356 5908 41412 6524
rect 41692 6580 41748 6590
rect 41692 6468 41748 6524
rect 41916 6580 41972 7310
rect 42252 7028 42308 7038
rect 42252 6914 42308 6972
rect 42252 6862 42254 6914
rect 42306 6862 42308 6914
rect 42252 6850 42308 6862
rect 42476 6692 42532 9662
rect 42588 8484 42644 9996
rect 42588 8370 42644 8428
rect 42588 8318 42590 8370
rect 42642 8318 42644 8370
rect 42588 8306 42644 8318
rect 42700 10610 42756 12126
rect 46844 12178 46900 12236
rect 46844 12126 46846 12178
rect 46898 12126 46900 12178
rect 46844 12114 46900 12126
rect 47852 12066 47908 12078
rect 47852 12014 47854 12066
rect 47906 12014 47908 12066
rect 47852 11844 47908 12014
rect 47852 11778 47908 11788
rect 43148 11396 43204 11406
rect 43036 11394 43204 11396
rect 43036 11342 43150 11394
rect 43202 11342 43204 11394
rect 43036 11340 43204 11342
rect 42924 11172 42980 11182
rect 42700 10558 42702 10610
rect 42754 10558 42756 10610
rect 42700 8260 42756 10558
rect 42700 8194 42756 8204
rect 42812 11170 42980 11172
rect 42812 11118 42926 11170
rect 42978 11118 42980 11170
rect 42812 11116 42980 11118
rect 42588 8148 42644 8158
rect 42588 7028 42644 8092
rect 42812 7700 42868 11116
rect 42924 11106 42980 11116
rect 42924 8372 42980 8382
rect 43036 8372 43092 11340
rect 43148 11330 43204 11340
rect 46844 10610 46900 10622
rect 46844 10558 46846 10610
rect 46898 10558 46900 10610
rect 46284 10498 46340 10510
rect 46284 10446 46286 10498
rect 46338 10446 46340 10498
rect 46284 10052 46340 10446
rect 46284 9986 46340 9996
rect 46844 10052 46900 10558
rect 47852 10498 47908 10510
rect 47852 10446 47854 10498
rect 47906 10446 47908 10498
rect 47852 10388 47908 10446
rect 47852 10322 47908 10332
rect 46844 9986 46900 9996
rect 42924 8370 43092 8372
rect 42924 8318 42926 8370
rect 42978 8318 43092 8370
rect 42924 8316 43092 8318
rect 46396 9044 46452 9054
rect 46844 9044 46900 9054
rect 46396 9042 46900 9044
rect 46396 8990 46398 9042
rect 46450 8990 46846 9042
rect 46898 8990 46900 9042
rect 46396 8988 46900 8990
rect 42924 8306 42980 8316
rect 46396 8148 46452 8988
rect 46844 8978 46900 8988
rect 47852 8932 47908 8942
rect 47852 8838 47908 8876
rect 46396 8082 46452 8092
rect 46844 8258 46900 8270
rect 46844 8206 46846 8258
rect 46898 8206 46900 8258
rect 46284 8034 46340 8046
rect 46284 7982 46286 8034
rect 46338 7982 46340 8034
rect 46284 7924 46340 7982
rect 46844 7924 46900 8206
rect 46284 7868 46900 7924
rect 47740 8146 47796 8158
rect 47740 8094 47742 8146
rect 47794 8094 47796 8146
rect 42812 7634 42868 7644
rect 42812 7362 42868 7374
rect 42812 7310 42814 7362
rect 42866 7310 42868 7362
rect 42812 7252 42868 7310
rect 42812 7186 42868 7196
rect 43260 7364 43316 7374
rect 43708 7364 43764 7374
rect 43260 7362 43764 7364
rect 43260 7310 43262 7362
rect 43314 7310 43710 7362
rect 43762 7310 43764 7362
rect 43260 7308 43764 7310
rect 42588 6962 42644 6972
rect 43260 6916 43316 7308
rect 43708 7298 43764 7308
rect 43932 7252 43988 7262
rect 43932 7158 43988 7196
rect 44268 7250 44324 7262
rect 44268 7198 44270 7250
rect 44322 7198 44324 7250
rect 43260 6850 43316 6860
rect 42588 6692 42644 6702
rect 42476 6690 42644 6692
rect 42476 6638 42590 6690
rect 42642 6638 42644 6690
rect 42476 6636 42644 6638
rect 42588 6626 42644 6636
rect 43484 6692 43540 6702
rect 43484 6598 43540 6636
rect 41916 6514 41972 6524
rect 41356 5842 41412 5852
rect 41468 6412 41748 6468
rect 42476 6468 42532 6478
rect 43260 6468 43316 6478
rect 41468 5348 41524 6412
rect 41776 6300 42352 6310
rect 41832 6244 41880 6300
rect 41936 6244 41984 6300
rect 42040 6244 42088 6300
rect 42144 6244 42192 6300
rect 42248 6244 42296 6300
rect 41776 6234 42352 6244
rect 41916 6132 41972 6142
rect 41916 6018 41972 6076
rect 41916 5966 41918 6018
rect 41970 5966 41972 6018
rect 41916 5954 41972 5966
rect 41356 5124 41412 5134
rect 41356 5010 41412 5068
rect 41356 4958 41358 5010
rect 41410 4958 41412 5010
rect 41356 4946 41412 4958
rect 41468 4564 41524 5292
rect 41692 5908 41748 5918
rect 41692 5460 41748 5852
rect 42476 5906 42532 6412
rect 43148 6466 43316 6468
rect 43148 6414 43262 6466
rect 43314 6414 43316 6466
rect 43148 6412 43316 6414
rect 42476 5854 42478 5906
rect 42530 5854 42532 5906
rect 42476 5842 42532 5854
rect 42812 5908 42868 5918
rect 42812 5814 42868 5852
rect 41692 5010 41748 5404
rect 42700 5460 42756 5470
rect 42252 5348 42308 5358
rect 42252 5254 42308 5292
rect 41692 4958 41694 5010
rect 41746 4958 41748 5010
rect 41692 4946 41748 4958
rect 41916 5122 41972 5134
rect 41916 5070 41918 5122
rect 41970 5070 41972 5122
rect 41916 4900 41972 5070
rect 41916 4844 42532 4900
rect 42476 4788 42532 4844
rect 41776 4732 42352 4742
rect 41832 4676 41880 4732
rect 41936 4676 41984 4732
rect 42040 4676 42088 4732
rect 42144 4676 42192 4732
rect 42248 4676 42296 4732
rect 41776 4666 42352 4676
rect 41580 4564 41636 4574
rect 41468 4562 41636 4564
rect 41468 4510 41582 4562
rect 41634 4510 41636 4562
rect 41468 4508 41636 4510
rect 41580 4498 41636 4508
rect 42476 4452 42532 4732
rect 42700 4562 42756 5404
rect 42924 4900 42980 4910
rect 42924 4806 42980 4844
rect 42700 4510 42702 4562
rect 42754 4510 42756 4562
rect 42700 4498 42756 4510
rect 41244 4396 41524 4452
rect 40796 4386 40852 4396
rect 41468 4340 41524 4396
rect 42476 4386 42532 4396
rect 41916 4340 41972 4350
rect 41468 4338 41972 4340
rect 41468 4286 41918 4338
rect 41970 4286 41972 4338
rect 41468 4284 41972 4286
rect 41916 4274 41972 4284
rect 37548 4226 37716 4228
rect 37548 4174 37550 4226
rect 37602 4174 37716 4226
rect 37548 4172 37716 4174
rect 37548 4162 37604 4172
rect 38056 3948 38632 3958
rect 38112 3892 38160 3948
rect 38216 3892 38264 3948
rect 38320 3892 38368 3948
rect 38424 3892 38472 3948
rect 38528 3892 38576 3948
rect 38056 3882 38632 3892
rect 37324 3614 37326 3666
rect 37378 3614 37380 3666
rect 37324 3602 37380 3614
rect 37884 3668 37940 3678
rect 37884 3574 37940 3612
rect 43148 3668 43204 6412
rect 43260 6402 43316 6412
rect 43484 6020 43540 6030
rect 43484 5926 43540 5964
rect 43708 5906 43764 5918
rect 43708 5854 43710 5906
rect 43762 5854 43764 5906
rect 43596 5460 43652 5470
rect 43596 5124 43652 5404
rect 43708 5348 43764 5854
rect 43708 5282 43764 5292
rect 43708 5124 43764 5134
rect 43596 5122 43764 5124
rect 43596 5070 43710 5122
rect 43762 5070 43764 5122
rect 43596 5068 43764 5070
rect 43708 5058 43764 5068
rect 44268 5124 44324 7198
rect 46284 6692 46340 6702
rect 46284 6132 46340 6636
rect 46396 6580 46452 7868
rect 47740 7476 47796 8094
rect 47740 7410 47796 7420
rect 46844 6692 46900 6702
rect 46844 6598 46900 6636
rect 46396 6514 46452 6524
rect 47740 6578 47796 6590
rect 47740 6526 47742 6578
rect 47794 6526 47796 6578
rect 46284 6066 46340 6076
rect 44380 6018 44436 6030
rect 44380 5966 44382 6018
rect 44434 5966 44436 6018
rect 44380 5236 44436 5966
rect 47740 6020 47796 6526
rect 47740 5954 47796 5964
rect 44604 5908 44660 5918
rect 44604 5814 44660 5852
rect 44380 5170 44436 5180
rect 46396 5684 46452 5694
rect 44268 5058 44324 5068
rect 46396 5124 46452 5628
rect 47852 5234 47908 5246
rect 47852 5182 47854 5234
rect 47906 5182 47908 5234
rect 46844 5124 46900 5134
rect 46396 5122 46900 5124
rect 46396 5070 46398 5122
rect 46450 5070 46846 5122
rect 46898 5070 46900 5122
rect 46396 5068 46900 5070
rect 46396 5058 46452 5068
rect 46844 5058 46900 5068
rect 43260 5012 43316 5022
rect 43260 4918 43316 4956
rect 43148 3602 43204 3612
rect 46396 4788 46452 4798
rect 46396 3556 46452 4732
rect 47852 4676 47908 5182
rect 47852 4610 47908 4620
rect 47180 4564 47236 4574
rect 47180 4470 47236 4508
rect 47740 4564 47796 4574
rect 47740 4470 47796 4508
rect 48076 4450 48132 4462
rect 48076 4398 48078 4450
rect 48130 4398 48132 4450
rect 46844 3556 46900 3566
rect 46396 3554 46900 3556
rect 46396 3502 46398 3554
rect 46450 3502 46846 3554
rect 46898 3502 46900 3554
rect 46396 3500 46900 3502
rect 46396 3490 46452 3500
rect 46844 3490 46900 3500
rect 37100 3378 37156 3388
rect 47740 3442 47796 3454
rect 47740 3390 47742 3442
rect 47794 3390 47796 3442
rect 8652 3332 8708 3342
rect 14140 3332 14196 3342
rect 19628 3332 19684 3342
rect 8540 3330 8708 3332
rect 8540 3278 8654 3330
rect 8706 3278 8708 3330
rect 8540 3276 8708 3278
rect 5776 3164 6352 3174
rect 5832 3108 5880 3164
rect 5936 3108 5984 3164
rect 6040 3108 6088 3164
rect 6144 3108 6192 3164
rect 6248 3108 6296 3164
rect 5776 3098 6352 3108
rect 8540 480 8596 3276
rect 8652 3266 8708 3276
rect 14028 3330 14196 3332
rect 14028 3278 14142 3330
rect 14194 3278 14196 3330
rect 14028 3276 14196 3278
rect 14028 480 14084 3276
rect 14140 3266 14196 3276
rect 19516 3330 19684 3332
rect 19516 3278 19630 3330
rect 19682 3278 19684 3330
rect 19516 3276 19684 3278
rect 19516 480 19572 3276
rect 19628 3266 19684 3276
rect 24556 3332 24612 3342
rect 24556 3330 24836 3332
rect 24556 3278 24558 3330
rect 24610 3278 24836 3330
rect 24556 3276 24836 3278
rect 24556 3266 24612 3276
rect 2856 392 3108 480
rect 8344 392 8596 480
rect 13832 392 14084 480
rect 19320 392 19572 480
rect 24780 480 24836 3276
rect 41776 3164 42352 3174
rect 41832 3108 41880 3164
rect 41936 3108 41984 3164
rect 42040 3108 42088 3164
rect 42144 3108 42192 3164
rect 42248 3108 42296 3164
rect 41776 3098 42352 3108
rect 47740 3108 47796 3390
rect 47740 3042 47796 3052
rect 48076 1652 48132 4398
rect 48076 1586 48132 1596
rect 24780 392 25032 480
rect 2856 -960 3080 392
rect 8344 -960 8568 392
rect 13832 -960 14056 392
rect 19320 -960 19544 392
rect 24808 -960 25032 392
rect 30296 -960 30520 480
rect 35784 -960 36008 480
rect 41272 -960 41496 480
rect 46760 -960 46984 480
<< via2 >>
rect 46060 48188 46116 48244
rect 1820 46396 1876 46452
rect 2056 46282 2112 46284
rect 2056 46230 2058 46282
rect 2058 46230 2110 46282
rect 2110 46230 2112 46282
rect 2056 46228 2112 46230
rect 2160 46282 2216 46284
rect 2160 46230 2162 46282
rect 2162 46230 2214 46282
rect 2214 46230 2216 46282
rect 2160 46228 2216 46230
rect 2264 46282 2320 46284
rect 2264 46230 2266 46282
rect 2266 46230 2318 46282
rect 2318 46230 2320 46282
rect 2264 46228 2320 46230
rect 2368 46282 2424 46284
rect 2368 46230 2370 46282
rect 2370 46230 2422 46282
rect 2422 46230 2424 46282
rect 2368 46228 2424 46230
rect 2472 46282 2528 46284
rect 2472 46230 2474 46282
rect 2474 46230 2526 46282
rect 2526 46230 2528 46282
rect 2472 46228 2528 46230
rect 2576 46282 2632 46284
rect 2576 46230 2578 46282
rect 2578 46230 2630 46282
rect 2630 46230 2632 46282
rect 2576 46228 2632 46230
rect 38056 46282 38112 46284
rect 38056 46230 38058 46282
rect 38058 46230 38110 46282
rect 38110 46230 38112 46282
rect 38056 46228 38112 46230
rect 38160 46282 38216 46284
rect 38160 46230 38162 46282
rect 38162 46230 38214 46282
rect 38214 46230 38216 46282
rect 38160 46228 38216 46230
rect 38264 46282 38320 46284
rect 38264 46230 38266 46282
rect 38266 46230 38318 46282
rect 38318 46230 38320 46282
rect 38264 46228 38320 46230
rect 38368 46282 38424 46284
rect 38368 46230 38370 46282
rect 38370 46230 38422 46282
rect 38422 46230 38424 46282
rect 38368 46228 38424 46230
rect 38472 46282 38528 46284
rect 38472 46230 38474 46282
rect 38474 46230 38526 46282
rect 38526 46230 38528 46282
rect 38472 46228 38528 46230
rect 38576 46282 38632 46284
rect 38576 46230 38578 46282
rect 38578 46230 38630 46282
rect 38630 46230 38632 46282
rect 38576 46228 38632 46230
rect 47852 46732 47908 46788
rect 5776 45498 5832 45500
rect 5776 45446 5778 45498
rect 5778 45446 5830 45498
rect 5830 45446 5832 45498
rect 5776 45444 5832 45446
rect 5880 45498 5936 45500
rect 5880 45446 5882 45498
rect 5882 45446 5934 45498
rect 5934 45446 5936 45498
rect 5880 45444 5936 45446
rect 5984 45498 6040 45500
rect 5984 45446 5986 45498
rect 5986 45446 6038 45498
rect 6038 45446 6040 45498
rect 5984 45444 6040 45446
rect 6088 45498 6144 45500
rect 6088 45446 6090 45498
rect 6090 45446 6142 45498
rect 6142 45446 6144 45498
rect 6088 45444 6144 45446
rect 6192 45498 6248 45500
rect 6192 45446 6194 45498
rect 6194 45446 6246 45498
rect 6246 45446 6248 45498
rect 6192 45444 6248 45446
rect 6296 45498 6352 45500
rect 6296 45446 6298 45498
rect 6298 45446 6350 45498
rect 6350 45446 6352 45498
rect 6296 45444 6352 45446
rect 41776 45498 41832 45500
rect 41776 45446 41778 45498
rect 41778 45446 41830 45498
rect 41830 45446 41832 45498
rect 41776 45444 41832 45446
rect 41880 45498 41936 45500
rect 41880 45446 41882 45498
rect 41882 45446 41934 45498
rect 41934 45446 41936 45498
rect 41880 45444 41936 45446
rect 41984 45498 42040 45500
rect 41984 45446 41986 45498
rect 41986 45446 42038 45498
rect 42038 45446 42040 45498
rect 41984 45444 42040 45446
rect 42088 45498 42144 45500
rect 42088 45446 42090 45498
rect 42090 45446 42142 45498
rect 42142 45446 42144 45498
rect 42088 45444 42144 45446
rect 42192 45498 42248 45500
rect 42192 45446 42194 45498
rect 42194 45446 42246 45498
rect 42246 45446 42248 45498
rect 42192 45444 42248 45446
rect 42296 45498 42352 45500
rect 42296 45446 42298 45498
rect 42298 45446 42350 45498
rect 42350 45446 42352 45498
rect 42296 45444 42352 45446
rect 2056 44714 2112 44716
rect 2056 44662 2058 44714
rect 2058 44662 2110 44714
rect 2110 44662 2112 44714
rect 2056 44660 2112 44662
rect 2160 44714 2216 44716
rect 2160 44662 2162 44714
rect 2162 44662 2214 44714
rect 2214 44662 2216 44714
rect 2160 44660 2216 44662
rect 2264 44714 2320 44716
rect 2264 44662 2266 44714
rect 2266 44662 2318 44714
rect 2318 44662 2320 44714
rect 2264 44660 2320 44662
rect 2368 44714 2424 44716
rect 2368 44662 2370 44714
rect 2370 44662 2422 44714
rect 2422 44662 2424 44714
rect 2368 44660 2424 44662
rect 2472 44714 2528 44716
rect 2472 44662 2474 44714
rect 2474 44662 2526 44714
rect 2526 44662 2528 44714
rect 2472 44660 2528 44662
rect 2576 44714 2632 44716
rect 2576 44662 2578 44714
rect 2578 44662 2630 44714
rect 2630 44662 2632 44714
rect 2576 44660 2632 44662
rect 38056 44714 38112 44716
rect 38056 44662 38058 44714
rect 38058 44662 38110 44714
rect 38110 44662 38112 44714
rect 38056 44660 38112 44662
rect 38160 44714 38216 44716
rect 38160 44662 38162 44714
rect 38162 44662 38214 44714
rect 38214 44662 38216 44714
rect 38160 44660 38216 44662
rect 38264 44714 38320 44716
rect 38264 44662 38266 44714
rect 38266 44662 38318 44714
rect 38318 44662 38320 44714
rect 38264 44660 38320 44662
rect 38368 44714 38424 44716
rect 38368 44662 38370 44714
rect 38370 44662 38422 44714
rect 38422 44662 38424 44714
rect 38368 44660 38424 44662
rect 38472 44714 38528 44716
rect 38472 44662 38474 44714
rect 38474 44662 38526 44714
rect 38526 44662 38528 44714
rect 38472 44660 38528 44662
rect 38576 44714 38632 44716
rect 38576 44662 38578 44714
rect 38578 44662 38630 44714
rect 38630 44662 38632 44714
rect 38576 44660 38632 44662
rect 5776 43930 5832 43932
rect 5776 43878 5778 43930
rect 5778 43878 5830 43930
rect 5830 43878 5832 43930
rect 5776 43876 5832 43878
rect 5880 43930 5936 43932
rect 5880 43878 5882 43930
rect 5882 43878 5934 43930
rect 5934 43878 5936 43930
rect 5880 43876 5936 43878
rect 5984 43930 6040 43932
rect 5984 43878 5986 43930
rect 5986 43878 6038 43930
rect 6038 43878 6040 43930
rect 5984 43876 6040 43878
rect 6088 43930 6144 43932
rect 6088 43878 6090 43930
rect 6090 43878 6142 43930
rect 6142 43878 6144 43930
rect 6088 43876 6144 43878
rect 6192 43930 6248 43932
rect 6192 43878 6194 43930
rect 6194 43878 6246 43930
rect 6246 43878 6248 43930
rect 6192 43876 6248 43878
rect 6296 43930 6352 43932
rect 6296 43878 6298 43930
rect 6298 43878 6350 43930
rect 6350 43878 6352 43930
rect 6296 43876 6352 43878
rect 41776 43930 41832 43932
rect 41776 43878 41778 43930
rect 41778 43878 41830 43930
rect 41830 43878 41832 43930
rect 41776 43876 41832 43878
rect 41880 43930 41936 43932
rect 41880 43878 41882 43930
rect 41882 43878 41934 43930
rect 41934 43878 41936 43930
rect 41880 43876 41936 43878
rect 41984 43930 42040 43932
rect 41984 43878 41986 43930
rect 41986 43878 42038 43930
rect 42038 43878 42040 43930
rect 41984 43876 42040 43878
rect 42088 43930 42144 43932
rect 42088 43878 42090 43930
rect 42090 43878 42142 43930
rect 42142 43878 42144 43930
rect 42088 43876 42144 43878
rect 42192 43930 42248 43932
rect 42192 43878 42194 43930
rect 42194 43878 42246 43930
rect 42246 43878 42248 43930
rect 42192 43876 42248 43878
rect 42296 43930 42352 43932
rect 42296 43878 42298 43930
rect 42298 43878 42350 43930
rect 42350 43878 42352 43930
rect 42296 43876 42352 43878
rect 2056 43146 2112 43148
rect 2056 43094 2058 43146
rect 2058 43094 2110 43146
rect 2110 43094 2112 43146
rect 2056 43092 2112 43094
rect 2160 43146 2216 43148
rect 2160 43094 2162 43146
rect 2162 43094 2214 43146
rect 2214 43094 2216 43146
rect 2160 43092 2216 43094
rect 2264 43146 2320 43148
rect 2264 43094 2266 43146
rect 2266 43094 2318 43146
rect 2318 43094 2320 43146
rect 2264 43092 2320 43094
rect 2368 43146 2424 43148
rect 2368 43094 2370 43146
rect 2370 43094 2422 43146
rect 2422 43094 2424 43146
rect 2368 43092 2424 43094
rect 2472 43146 2528 43148
rect 2472 43094 2474 43146
rect 2474 43094 2526 43146
rect 2526 43094 2528 43146
rect 2472 43092 2528 43094
rect 2576 43146 2632 43148
rect 2576 43094 2578 43146
rect 2578 43094 2630 43146
rect 2630 43094 2632 43146
rect 2576 43092 2632 43094
rect 38056 43146 38112 43148
rect 38056 43094 38058 43146
rect 38058 43094 38110 43146
rect 38110 43094 38112 43146
rect 38056 43092 38112 43094
rect 38160 43146 38216 43148
rect 38160 43094 38162 43146
rect 38162 43094 38214 43146
rect 38214 43094 38216 43146
rect 38160 43092 38216 43094
rect 38264 43146 38320 43148
rect 38264 43094 38266 43146
rect 38266 43094 38318 43146
rect 38318 43094 38320 43146
rect 38264 43092 38320 43094
rect 38368 43146 38424 43148
rect 38368 43094 38370 43146
rect 38370 43094 38422 43146
rect 38422 43094 38424 43146
rect 38368 43092 38424 43094
rect 38472 43146 38528 43148
rect 38472 43094 38474 43146
rect 38474 43094 38526 43146
rect 38526 43094 38528 43146
rect 38472 43092 38528 43094
rect 38576 43146 38632 43148
rect 38576 43094 38578 43146
rect 38578 43094 38630 43146
rect 38630 43094 38632 43146
rect 38576 43092 38632 43094
rect 5776 42362 5832 42364
rect 5776 42310 5778 42362
rect 5778 42310 5830 42362
rect 5830 42310 5832 42362
rect 5776 42308 5832 42310
rect 5880 42362 5936 42364
rect 5880 42310 5882 42362
rect 5882 42310 5934 42362
rect 5934 42310 5936 42362
rect 5880 42308 5936 42310
rect 5984 42362 6040 42364
rect 5984 42310 5986 42362
rect 5986 42310 6038 42362
rect 6038 42310 6040 42362
rect 5984 42308 6040 42310
rect 6088 42362 6144 42364
rect 6088 42310 6090 42362
rect 6090 42310 6142 42362
rect 6142 42310 6144 42362
rect 6088 42308 6144 42310
rect 6192 42362 6248 42364
rect 6192 42310 6194 42362
rect 6194 42310 6246 42362
rect 6246 42310 6248 42362
rect 6192 42308 6248 42310
rect 6296 42362 6352 42364
rect 6296 42310 6298 42362
rect 6298 42310 6350 42362
rect 6350 42310 6352 42362
rect 6296 42308 6352 42310
rect 41776 42362 41832 42364
rect 41776 42310 41778 42362
rect 41778 42310 41830 42362
rect 41830 42310 41832 42362
rect 41776 42308 41832 42310
rect 41880 42362 41936 42364
rect 41880 42310 41882 42362
rect 41882 42310 41934 42362
rect 41934 42310 41936 42362
rect 41880 42308 41936 42310
rect 41984 42362 42040 42364
rect 41984 42310 41986 42362
rect 41986 42310 42038 42362
rect 42038 42310 42040 42362
rect 41984 42308 42040 42310
rect 42088 42362 42144 42364
rect 42088 42310 42090 42362
rect 42090 42310 42142 42362
rect 42142 42310 42144 42362
rect 42088 42308 42144 42310
rect 42192 42362 42248 42364
rect 42192 42310 42194 42362
rect 42194 42310 42246 42362
rect 42246 42310 42248 42362
rect 42192 42308 42248 42310
rect 42296 42362 42352 42364
rect 42296 42310 42298 42362
rect 42298 42310 42350 42362
rect 42350 42310 42352 42362
rect 42296 42308 42352 42310
rect 40236 41916 40292 41972
rect 2056 41578 2112 41580
rect 2056 41526 2058 41578
rect 2058 41526 2110 41578
rect 2110 41526 2112 41578
rect 2056 41524 2112 41526
rect 2160 41578 2216 41580
rect 2160 41526 2162 41578
rect 2162 41526 2214 41578
rect 2214 41526 2216 41578
rect 2160 41524 2216 41526
rect 2264 41578 2320 41580
rect 2264 41526 2266 41578
rect 2266 41526 2318 41578
rect 2318 41526 2320 41578
rect 2264 41524 2320 41526
rect 2368 41578 2424 41580
rect 2368 41526 2370 41578
rect 2370 41526 2422 41578
rect 2422 41526 2424 41578
rect 2368 41524 2424 41526
rect 2472 41578 2528 41580
rect 2472 41526 2474 41578
rect 2474 41526 2526 41578
rect 2526 41526 2528 41578
rect 2472 41524 2528 41526
rect 2576 41578 2632 41580
rect 2576 41526 2578 41578
rect 2578 41526 2630 41578
rect 2630 41526 2632 41578
rect 2576 41524 2632 41526
rect 38056 41578 38112 41580
rect 38056 41526 38058 41578
rect 38058 41526 38110 41578
rect 38110 41526 38112 41578
rect 38056 41524 38112 41526
rect 38160 41578 38216 41580
rect 38160 41526 38162 41578
rect 38162 41526 38214 41578
rect 38214 41526 38216 41578
rect 38160 41524 38216 41526
rect 38264 41578 38320 41580
rect 38264 41526 38266 41578
rect 38266 41526 38318 41578
rect 38318 41526 38320 41578
rect 38264 41524 38320 41526
rect 38368 41578 38424 41580
rect 38368 41526 38370 41578
rect 38370 41526 38422 41578
rect 38422 41526 38424 41578
rect 38368 41524 38424 41526
rect 38472 41578 38528 41580
rect 38472 41526 38474 41578
rect 38474 41526 38526 41578
rect 38526 41526 38528 41578
rect 38472 41524 38528 41526
rect 38576 41578 38632 41580
rect 38576 41526 38578 41578
rect 38578 41526 38630 41578
rect 38630 41526 38632 41578
rect 38576 41524 38632 41526
rect 3052 40908 3108 40964
rect 3500 40962 3556 40964
rect 3500 40910 3502 40962
rect 3502 40910 3554 40962
rect 3554 40910 3556 40962
rect 3500 40908 3556 40910
rect 17948 40908 18004 40964
rect 5776 40794 5832 40796
rect 5776 40742 5778 40794
rect 5778 40742 5830 40794
rect 5830 40742 5832 40794
rect 5776 40740 5832 40742
rect 5880 40794 5936 40796
rect 5880 40742 5882 40794
rect 5882 40742 5934 40794
rect 5934 40742 5936 40794
rect 5880 40740 5936 40742
rect 5984 40794 6040 40796
rect 5984 40742 5986 40794
rect 5986 40742 6038 40794
rect 6038 40742 6040 40794
rect 5984 40740 6040 40742
rect 6088 40794 6144 40796
rect 6088 40742 6090 40794
rect 6090 40742 6142 40794
rect 6142 40742 6144 40794
rect 6088 40740 6144 40742
rect 6192 40794 6248 40796
rect 6192 40742 6194 40794
rect 6194 40742 6246 40794
rect 6246 40742 6248 40794
rect 6192 40740 6248 40742
rect 6296 40794 6352 40796
rect 6296 40742 6298 40794
rect 6298 40742 6350 40794
rect 6350 40742 6352 40794
rect 6296 40740 6352 40742
rect 2156 40460 2212 40516
rect 2056 40010 2112 40012
rect 2056 39958 2058 40010
rect 2058 39958 2110 40010
rect 2110 39958 2112 40010
rect 2056 39956 2112 39958
rect 2160 40010 2216 40012
rect 2160 39958 2162 40010
rect 2162 39958 2214 40010
rect 2214 39958 2216 40010
rect 2160 39956 2216 39958
rect 2264 40010 2320 40012
rect 2264 39958 2266 40010
rect 2266 39958 2318 40010
rect 2318 39958 2320 40010
rect 2264 39956 2320 39958
rect 2368 40010 2424 40012
rect 2368 39958 2370 40010
rect 2370 39958 2422 40010
rect 2422 39958 2424 40010
rect 2368 39956 2424 39958
rect 2472 40010 2528 40012
rect 2472 39958 2474 40010
rect 2474 39958 2526 40010
rect 2526 39958 2528 40010
rect 2472 39956 2528 39958
rect 2576 40010 2632 40012
rect 2576 39958 2578 40010
rect 2578 39958 2630 40010
rect 2630 39958 2632 40010
rect 2576 39956 2632 39958
rect 5776 39226 5832 39228
rect 5776 39174 5778 39226
rect 5778 39174 5830 39226
rect 5830 39174 5832 39226
rect 5776 39172 5832 39174
rect 5880 39226 5936 39228
rect 5880 39174 5882 39226
rect 5882 39174 5934 39226
rect 5934 39174 5936 39226
rect 5880 39172 5936 39174
rect 5984 39226 6040 39228
rect 5984 39174 5986 39226
rect 5986 39174 6038 39226
rect 6038 39174 6040 39226
rect 5984 39172 6040 39174
rect 6088 39226 6144 39228
rect 6088 39174 6090 39226
rect 6090 39174 6142 39226
rect 6142 39174 6144 39226
rect 6088 39172 6144 39174
rect 6192 39226 6248 39228
rect 6192 39174 6194 39226
rect 6194 39174 6246 39226
rect 6246 39174 6248 39226
rect 6192 39172 6248 39174
rect 6296 39226 6352 39228
rect 6296 39174 6298 39226
rect 6298 39174 6350 39226
rect 6350 39174 6352 39226
rect 6296 39172 6352 39174
rect 2056 38442 2112 38444
rect 2056 38390 2058 38442
rect 2058 38390 2110 38442
rect 2110 38390 2112 38442
rect 2056 38388 2112 38390
rect 2160 38442 2216 38444
rect 2160 38390 2162 38442
rect 2162 38390 2214 38442
rect 2214 38390 2216 38442
rect 2160 38388 2216 38390
rect 2264 38442 2320 38444
rect 2264 38390 2266 38442
rect 2266 38390 2318 38442
rect 2318 38390 2320 38442
rect 2264 38388 2320 38390
rect 2368 38442 2424 38444
rect 2368 38390 2370 38442
rect 2370 38390 2422 38442
rect 2422 38390 2424 38442
rect 2368 38388 2424 38390
rect 2472 38442 2528 38444
rect 2472 38390 2474 38442
rect 2474 38390 2526 38442
rect 2526 38390 2528 38442
rect 2472 38388 2528 38390
rect 2576 38442 2632 38444
rect 2576 38390 2578 38442
rect 2578 38390 2630 38442
rect 2630 38390 2632 38442
rect 2576 38388 2632 38390
rect 5776 37658 5832 37660
rect 5776 37606 5778 37658
rect 5778 37606 5830 37658
rect 5830 37606 5832 37658
rect 5776 37604 5832 37606
rect 5880 37658 5936 37660
rect 5880 37606 5882 37658
rect 5882 37606 5934 37658
rect 5934 37606 5936 37658
rect 5880 37604 5936 37606
rect 5984 37658 6040 37660
rect 5984 37606 5986 37658
rect 5986 37606 6038 37658
rect 6038 37606 6040 37658
rect 5984 37604 6040 37606
rect 6088 37658 6144 37660
rect 6088 37606 6090 37658
rect 6090 37606 6142 37658
rect 6142 37606 6144 37658
rect 6088 37604 6144 37606
rect 6192 37658 6248 37660
rect 6192 37606 6194 37658
rect 6194 37606 6246 37658
rect 6246 37606 6248 37658
rect 6192 37604 6248 37606
rect 6296 37658 6352 37660
rect 6296 37606 6298 37658
rect 6298 37606 6350 37658
rect 6350 37606 6352 37658
rect 6296 37604 6352 37606
rect 2056 36874 2112 36876
rect 2056 36822 2058 36874
rect 2058 36822 2110 36874
rect 2110 36822 2112 36874
rect 2056 36820 2112 36822
rect 2160 36874 2216 36876
rect 2160 36822 2162 36874
rect 2162 36822 2214 36874
rect 2214 36822 2216 36874
rect 2160 36820 2216 36822
rect 2264 36874 2320 36876
rect 2264 36822 2266 36874
rect 2266 36822 2318 36874
rect 2318 36822 2320 36874
rect 2264 36820 2320 36822
rect 2368 36874 2424 36876
rect 2368 36822 2370 36874
rect 2370 36822 2422 36874
rect 2422 36822 2424 36874
rect 2368 36820 2424 36822
rect 2472 36874 2528 36876
rect 2472 36822 2474 36874
rect 2474 36822 2526 36874
rect 2526 36822 2528 36874
rect 2472 36820 2528 36822
rect 2576 36874 2632 36876
rect 2576 36822 2578 36874
rect 2578 36822 2630 36874
rect 2630 36822 2632 36874
rect 2576 36820 2632 36822
rect 17388 36316 17444 36372
rect 38056 40010 38112 40012
rect 38056 39958 38058 40010
rect 38058 39958 38110 40010
rect 38110 39958 38112 40010
rect 38056 39956 38112 39958
rect 38160 40010 38216 40012
rect 38160 39958 38162 40010
rect 38162 39958 38214 40010
rect 38214 39958 38216 40010
rect 38160 39956 38216 39958
rect 38264 40010 38320 40012
rect 38264 39958 38266 40010
rect 38266 39958 38318 40010
rect 38318 39958 38320 40010
rect 38264 39956 38320 39958
rect 38368 40010 38424 40012
rect 38368 39958 38370 40010
rect 38370 39958 38422 40010
rect 38422 39958 38424 40010
rect 38368 39956 38424 39958
rect 38472 40010 38528 40012
rect 38472 39958 38474 40010
rect 38474 39958 38526 40010
rect 38526 39958 38528 40010
rect 38472 39956 38528 39958
rect 38576 40010 38632 40012
rect 38576 39958 38578 40010
rect 38578 39958 38630 40010
rect 38630 39958 38632 40010
rect 38576 39956 38632 39958
rect 38056 38442 38112 38444
rect 38056 38390 38058 38442
rect 38058 38390 38110 38442
rect 38110 38390 38112 38442
rect 38056 38388 38112 38390
rect 38160 38442 38216 38444
rect 38160 38390 38162 38442
rect 38162 38390 38214 38442
rect 38214 38390 38216 38442
rect 38160 38388 38216 38390
rect 38264 38442 38320 38444
rect 38264 38390 38266 38442
rect 38266 38390 38318 38442
rect 38318 38390 38320 38442
rect 38264 38388 38320 38390
rect 38368 38442 38424 38444
rect 38368 38390 38370 38442
rect 38370 38390 38422 38442
rect 38422 38390 38424 38442
rect 38368 38388 38424 38390
rect 38472 38442 38528 38444
rect 38472 38390 38474 38442
rect 38474 38390 38526 38442
rect 38526 38390 38528 38442
rect 38472 38388 38528 38390
rect 38576 38442 38632 38444
rect 38576 38390 38578 38442
rect 38578 38390 38630 38442
rect 38630 38390 38632 38442
rect 38576 38388 38632 38390
rect 38056 36874 38112 36876
rect 38056 36822 38058 36874
rect 38058 36822 38110 36874
rect 38110 36822 38112 36874
rect 38056 36820 38112 36822
rect 38160 36874 38216 36876
rect 38160 36822 38162 36874
rect 38162 36822 38214 36874
rect 38214 36822 38216 36874
rect 38160 36820 38216 36822
rect 38264 36874 38320 36876
rect 38264 36822 38266 36874
rect 38266 36822 38318 36874
rect 38318 36822 38320 36874
rect 38264 36820 38320 36822
rect 38368 36874 38424 36876
rect 38368 36822 38370 36874
rect 38370 36822 38422 36874
rect 38422 36822 38424 36874
rect 38368 36820 38424 36822
rect 38472 36874 38528 36876
rect 38472 36822 38474 36874
rect 38474 36822 38526 36874
rect 38526 36822 38528 36874
rect 38472 36820 38528 36822
rect 38576 36874 38632 36876
rect 38576 36822 38578 36874
rect 38578 36822 38630 36874
rect 38630 36822 38632 36874
rect 38576 36820 38632 36822
rect 18284 36370 18340 36372
rect 18284 36318 18286 36370
rect 18286 36318 18338 36370
rect 18338 36318 18340 36370
rect 18284 36316 18340 36318
rect 5776 36090 5832 36092
rect 5776 36038 5778 36090
rect 5778 36038 5830 36090
rect 5830 36038 5832 36090
rect 5776 36036 5832 36038
rect 5880 36090 5936 36092
rect 5880 36038 5882 36090
rect 5882 36038 5934 36090
rect 5934 36038 5936 36090
rect 5880 36036 5936 36038
rect 5984 36090 6040 36092
rect 5984 36038 5986 36090
rect 5986 36038 6038 36090
rect 6038 36038 6040 36090
rect 5984 36036 6040 36038
rect 6088 36090 6144 36092
rect 6088 36038 6090 36090
rect 6090 36038 6142 36090
rect 6142 36038 6144 36090
rect 6088 36036 6144 36038
rect 6192 36090 6248 36092
rect 6192 36038 6194 36090
rect 6194 36038 6246 36090
rect 6246 36038 6248 36090
rect 6192 36036 6248 36038
rect 6296 36090 6352 36092
rect 6296 36038 6298 36090
rect 6298 36038 6350 36090
rect 6350 36038 6352 36090
rect 6296 36036 6352 36038
rect 2056 35306 2112 35308
rect 2056 35254 2058 35306
rect 2058 35254 2110 35306
rect 2110 35254 2112 35306
rect 2056 35252 2112 35254
rect 2160 35306 2216 35308
rect 2160 35254 2162 35306
rect 2162 35254 2214 35306
rect 2214 35254 2216 35306
rect 2160 35252 2216 35254
rect 2264 35306 2320 35308
rect 2264 35254 2266 35306
rect 2266 35254 2318 35306
rect 2318 35254 2320 35306
rect 2264 35252 2320 35254
rect 2368 35306 2424 35308
rect 2368 35254 2370 35306
rect 2370 35254 2422 35306
rect 2422 35254 2424 35306
rect 2368 35252 2424 35254
rect 2472 35306 2528 35308
rect 2472 35254 2474 35306
rect 2474 35254 2526 35306
rect 2526 35254 2528 35306
rect 2472 35252 2528 35254
rect 2576 35306 2632 35308
rect 2576 35254 2578 35306
rect 2578 35254 2630 35306
rect 2630 35254 2632 35306
rect 2576 35252 2632 35254
rect 5776 34522 5832 34524
rect 5776 34470 5778 34522
rect 5778 34470 5830 34522
rect 5830 34470 5832 34522
rect 5776 34468 5832 34470
rect 5880 34522 5936 34524
rect 5880 34470 5882 34522
rect 5882 34470 5934 34522
rect 5934 34470 5936 34522
rect 5880 34468 5936 34470
rect 5984 34522 6040 34524
rect 5984 34470 5986 34522
rect 5986 34470 6038 34522
rect 6038 34470 6040 34522
rect 5984 34468 6040 34470
rect 6088 34522 6144 34524
rect 6088 34470 6090 34522
rect 6090 34470 6142 34522
rect 6142 34470 6144 34522
rect 6088 34468 6144 34470
rect 6192 34522 6248 34524
rect 6192 34470 6194 34522
rect 6194 34470 6246 34522
rect 6246 34470 6248 34522
rect 6192 34468 6248 34470
rect 6296 34522 6352 34524
rect 6296 34470 6298 34522
rect 6298 34470 6350 34522
rect 6350 34470 6352 34522
rect 6296 34468 6352 34470
rect 1820 34300 1876 34356
rect 2056 33738 2112 33740
rect 2056 33686 2058 33738
rect 2058 33686 2110 33738
rect 2110 33686 2112 33738
rect 2056 33684 2112 33686
rect 2160 33738 2216 33740
rect 2160 33686 2162 33738
rect 2162 33686 2214 33738
rect 2214 33686 2216 33738
rect 2160 33684 2216 33686
rect 2264 33738 2320 33740
rect 2264 33686 2266 33738
rect 2266 33686 2318 33738
rect 2318 33686 2320 33738
rect 2264 33684 2320 33686
rect 2368 33738 2424 33740
rect 2368 33686 2370 33738
rect 2370 33686 2422 33738
rect 2422 33686 2424 33738
rect 2368 33684 2424 33686
rect 2472 33738 2528 33740
rect 2472 33686 2474 33738
rect 2474 33686 2526 33738
rect 2526 33686 2528 33738
rect 2472 33684 2528 33686
rect 2576 33738 2632 33740
rect 2576 33686 2578 33738
rect 2578 33686 2630 33738
rect 2630 33686 2632 33738
rect 2576 33684 2632 33686
rect 5776 32954 5832 32956
rect 5776 32902 5778 32954
rect 5778 32902 5830 32954
rect 5830 32902 5832 32954
rect 5776 32900 5832 32902
rect 5880 32954 5936 32956
rect 5880 32902 5882 32954
rect 5882 32902 5934 32954
rect 5934 32902 5936 32954
rect 5880 32900 5936 32902
rect 5984 32954 6040 32956
rect 5984 32902 5986 32954
rect 5986 32902 6038 32954
rect 6038 32902 6040 32954
rect 5984 32900 6040 32902
rect 6088 32954 6144 32956
rect 6088 32902 6090 32954
rect 6090 32902 6142 32954
rect 6142 32902 6144 32954
rect 6088 32900 6144 32902
rect 6192 32954 6248 32956
rect 6192 32902 6194 32954
rect 6194 32902 6246 32954
rect 6246 32902 6248 32954
rect 6192 32900 6248 32902
rect 6296 32954 6352 32956
rect 6296 32902 6298 32954
rect 6298 32902 6350 32954
rect 6350 32902 6352 32954
rect 6296 32900 6352 32902
rect 2056 32170 2112 32172
rect 2056 32118 2058 32170
rect 2058 32118 2110 32170
rect 2110 32118 2112 32170
rect 2056 32116 2112 32118
rect 2160 32170 2216 32172
rect 2160 32118 2162 32170
rect 2162 32118 2214 32170
rect 2214 32118 2216 32170
rect 2160 32116 2216 32118
rect 2264 32170 2320 32172
rect 2264 32118 2266 32170
rect 2266 32118 2318 32170
rect 2318 32118 2320 32170
rect 2264 32116 2320 32118
rect 2368 32170 2424 32172
rect 2368 32118 2370 32170
rect 2370 32118 2422 32170
rect 2422 32118 2424 32170
rect 2368 32116 2424 32118
rect 2472 32170 2528 32172
rect 2472 32118 2474 32170
rect 2474 32118 2526 32170
rect 2526 32118 2528 32170
rect 2472 32116 2528 32118
rect 2576 32170 2632 32172
rect 2576 32118 2578 32170
rect 2578 32118 2630 32170
rect 2630 32118 2632 32170
rect 2576 32116 2632 32118
rect 5776 31386 5832 31388
rect 5776 31334 5778 31386
rect 5778 31334 5830 31386
rect 5830 31334 5832 31386
rect 5776 31332 5832 31334
rect 5880 31386 5936 31388
rect 5880 31334 5882 31386
rect 5882 31334 5934 31386
rect 5934 31334 5936 31386
rect 5880 31332 5936 31334
rect 5984 31386 6040 31388
rect 5984 31334 5986 31386
rect 5986 31334 6038 31386
rect 6038 31334 6040 31386
rect 5984 31332 6040 31334
rect 6088 31386 6144 31388
rect 6088 31334 6090 31386
rect 6090 31334 6142 31386
rect 6142 31334 6144 31386
rect 6088 31332 6144 31334
rect 6192 31386 6248 31388
rect 6192 31334 6194 31386
rect 6194 31334 6246 31386
rect 6246 31334 6248 31386
rect 6192 31332 6248 31334
rect 6296 31386 6352 31388
rect 6296 31334 6298 31386
rect 6298 31334 6350 31386
rect 6350 31334 6352 31386
rect 6296 31332 6352 31334
rect 2056 30602 2112 30604
rect 2056 30550 2058 30602
rect 2058 30550 2110 30602
rect 2110 30550 2112 30602
rect 2056 30548 2112 30550
rect 2160 30602 2216 30604
rect 2160 30550 2162 30602
rect 2162 30550 2214 30602
rect 2214 30550 2216 30602
rect 2160 30548 2216 30550
rect 2264 30602 2320 30604
rect 2264 30550 2266 30602
rect 2266 30550 2318 30602
rect 2318 30550 2320 30602
rect 2264 30548 2320 30550
rect 2368 30602 2424 30604
rect 2368 30550 2370 30602
rect 2370 30550 2422 30602
rect 2422 30550 2424 30602
rect 2368 30548 2424 30550
rect 2472 30602 2528 30604
rect 2472 30550 2474 30602
rect 2474 30550 2526 30602
rect 2526 30550 2528 30602
rect 2472 30548 2528 30550
rect 2576 30602 2632 30604
rect 2576 30550 2578 30602
rect 2578 30550 2630 30602
rect 2630 30550 2632 30602
rect 2576 30548 2632 30550
rect 5776 29818 5832 29820
rect 5776 29766 5778 29818
rect 5778 29766 5830 29818
rect 5830 29766 5832 29818
rect 5776 29764 5832 29766
rect 5880 29818 5936 29820
rect 5880 29766 5882 29818
rect 5882 29766 5934 29818
rect 5934 29766 5936 29818
rect 5880 29764 5936 29766
rect 5984 29818 6040 29820
rect 5984 29766 5986 29818
rect 5986 29766 6038 29818
rect 6038 29766 6040 29818
rect 5984 29764 6040 29766
rect 6088 29818 6144 29820
rect 6088 29766 6090 29818
rect 6090 29766 6142 29818
rect 6142 29766 6144 29818
rect 6088 29764 6144 29766
rect 6192 29818 6248 29820
rect 6192 29766 6194 29818
rect 6194 29766 6246 29818
rect 6246 29766 6248 29818
rect 6192 29764 6248 29766
rect 6296 29818 6352 29820
rect 6296 29766 6298 29818
rect 6298 29766 6350 29818
rect 6350 29766 6352 29818
rect 6296 29764 6352 29766
rect 2056 29034 2112 29036
rect 2056 28982 2058 29034
rect 2058 28982 2110 29034
rect 2110 28982 2112 29034
rect 2056 28980 2112 28982
rect 2160 29034 2216 29036
rect 2160 28982 2162 29034
rect 2162 28982 2214 29034
rect 2214 28982 2216 29034
rect 2160 28980 2216 28982
rect 2264 29034 2320 29036
rect 2264 28982 2266 29034
rect 2266 28982 2318 29034
rect 2318 28982 2320 29034
rect 2264 28980 2320 28982
rect 2368 29034 2424 29036
rect 2368 28982 2370 29034
rect 2370 28982 2422 29034
rect 2422 28982 2424 29034
rect 2368 28980 2424 28982
rect 2472 29034 2528 29036
rect 2472 28982 2474 29034
rect 2474 28982 2526 29034
rect 2526 28982 2528 29034
rect 2472 28980 2528 28982
rect 2576 29034 2632 29036
rect 2576 28982 2578 29034
rect 2578 28982 2630 29034
rect 2630 28982 2632 29034
rect 2576 28980 2632 28982
rect 1820 28082 1876 28084
rect 1820 28030 1822 28082
rect 1822 28030 1874 28082
rect 1874 28030 1876 28082
rect 1820 28028 1876 28030
rect 2056 27466 2112 27468
rect 2056 27414 2058 27466
rect 2058 27414 2110 27466
rect 2110 27414 2112 27466
rect 2056 27412 2112 27414
rect 2160 27466 2216 27468
rect 2160 27414 2162 27466
rect 2162 27414 2214 27466
rect 2214 27414 2216 27466
rect 2160 27412 2216 27414
rect 2264 27466 2320 27468
rect 2264 27414 2266 27466
rect 2266 27414 2318 27466
rect 2318 27414 2320 27466
rect 2264 27412 2320 27414
rect 2368 27466 2424 27468
rect 2368 27414 2370 27466
rect 2370 27414 2422 27466
rect 2422 27414 2424 27466
rect 2368 27412 2424 27414
rect 2472 27466 2528 27468
rect 2472 27414 2474 27466
rect 2474 27414 2526 27466
rect 2526 27414 2528 27466
rect 2472 27412 2528 27414
rect 2576 27466 2632 27468
rect 2576 27414 2578 27466
rect 2578 27414 2630 27466
rect 2630 27414 2632 27466
rect 2576 27412 2632 27414
rect 2056 25898 2112 25900
rect 2056 25846 2058 25898
rect 2058 25846 2110 25898
rect 2110 25846 2112 25898
rect 2056 25844 2112 25846
rect 2160 25898 2216 25900
rect 2160 25846 2162 25898
rect 2162 25846 2214 25898
rect 2214 25846 2216 25898
rect 2160 25844 2216 25846
rect 2264 25898 2320 25900
rect 2264 25846 2266 25898
rect 2266 25846 2318 25898
rect 2318 25846 2320 25898
rect 2264 25844 2320 25846
rect 2368 25898 2424 25900
rect 2368 25846 2370 25898
rect 2370 25846 2422 25898
rect 2422 25846 2424 25898
rect 2368 25844 2424 25846
rect 2472 25898 2528 25900
rect 2472 25846 2474 25898
rect 2474 25846 2526 25898
rect 2526 25846 2528 25898
rect 2472 25844 2528 25846
rect 2576 25898 2632 25900
rect 2576 25846 2578 25898
rect 2578 25846 2630 25898
rect 2630 25846 2632 25898
rect 2576 25844 2632 25846
rect 2056 24330 2112 24332
rect 2056 24278 2058 24330
rect 2058 24278 2110 24330
rect 2110 24278 2112 24330
rect 2056 24276 2112 24278
rect 2160 24330 2216 24332
rect 2160 24278 2162 24330
rect 2162 24278 2214 24330
rect 2214 24278 2216 24330
rect 2160 24276 2216 24278
rect 2264 24330 2320 24332
rect 2264 24278 2266 24330
rect 2266 24278 2318 24330
rect 2318 24278 2320 24330
rect 2264 24276 2320 24278
rect 2368 24330 2424 24332
rect 2368 24278 2370 24330
rect 2370 24278 2422 24330
rect 2422 24278 2424 24330
rect 2368 24276 2424 24278
rect 2472 24330 2528 24332
rect 2472 24278 2474 24330
rect 2474 24278 2526 24330
rect 2526 24278 2528 24330
rect 2472 24276 2528 24278
rect 2576 24330 2632 24332
rect 2576 24278 2578 24330
rect 2578 24278 2630 24330
rect 2630 24278 2632 24330
rect 2576 24276 2632 24278
rect 2056 22762 2112 22764
rect 2056 22710 2058 22762
rect 2058 22710 2110 22762
rect 2110 22710 2112 22762
rect 2056 22708 2112 22710
rect 2160 22762 2216 22764
rect 2160 22710 2162 22762
rect 2162 22710 2214 22762
rect 2214 22710 2216 22762
rect 2160 22708 2216 22710
rect 2264 22762 2320 22764
rect 2264 22710 2266 22762
rect 2266 22710 2318 22762
rect 2318 22710 2320 22762
rect 2264 22708 2320 22710
rect 2368 22762 2424 22764
rect 2368 22710 2370 22762
rect 2370 22710 2422 22762
rect 2422 22710 2424 22762
rect 2368 22708 2424 22710
rect 2472 22762 2528 22764
rect 2472 22710 2474 22762
rect 2474 22710 2526 22762
rect 2526 22710 2528 22762
rect 2472 22708 2528 22710
rect 2576 22762 2632 22764
rect 2576 22710 2578 22762
rect 2578 22710 2630 22762
rect 2630 22710 2632 22762
rect 2576 22708 2632 22710
rect 1820 21980 1876 22036
rect 2056 21194 2112 21196
rect 2056 21142 2058 21194
rect 2058 21142 2110 21194
rect 2110 21142 2112 21194
rect 2056 21140 2112 21142
rect 2160 21194 2216 21196
rect 2160 21142 2162 21194
rect 2162 21142 2214 21194
rect 2214 21142 2216 21194
rect 2160 21140 2216 21142
rect 2264 21194 2320 21196
rect 2264 21142 2266 21194
rect 2266 21142 2318 21194
rect 2318 21142 2320 21194
rect 2264 21140 2320 21142
rect 2368 21194 2424 21196
rect 2368 21142 2370 21194
rect 2370 21142 2422 21194
rect 2422 21142 2424 21194
rect 2368 21140 2424 21142
rect 2472 21194 2528 21196
rect 2472 21142 2474 21194
rect 2474 21142 2526 21194
rect 2526 21142 2528 21194
rect 2472 21140 2528 21142
rect 2576 21194 2632 21196
rect 2576 21142 2578 21194
rect 2578 21142 2630 21194
rect 2630 21142 2632 21194
rect 2576 21140 2632 21142
rect 2056 19626 2112 19628
rect 2056 19574 2058 19626
rect 2058 19574 2110 19626
rect 2110 19574 2112 19626
rect 2056 19572 2112 19574
rect 2160 19626 2216 19628
rect 2160 19574 2162 19626
rect 2162 19574 2214 19626
rect 2214 19574 2216 19626
rect 2160 19572 2216 19574
rect 2264 19626 2320 19628
rect 2264 19574 2266 19626
rect 2266 19574 2318 19626
rect 2318 19574 2320 19626
rect 2264 19572 2320 19574
rect 2368 19626 2424 19628
rect 2368 19574 2370 19626
rect 2370 19574 2422 19626
rect 2422 19574 2424 19626
rect 2368 19572 2424 19574
rect 2472 19626 2528 19628
rect 2472 19574 2474 19626
rect 2474 19574 2526 19626
rect 2526 19574 2528 19626
rect 2472 19572 2528 19574
rect 2576 19626 2632 19628
rect 2576 19574 2578 19626
rect 2578 19574 2630 19626
rect 2630 19574 2632 19626
rect 2576 19572 2632 19574
rect 2056 18058 2112 18060
rect 2056 18006 2058 18058
rect 2058 18006 2110 18058
rect 2110 18006 2112 18058
rect 2056 18004 2112 18006
rect 2160 18058 2216 18060
rect 2160 18006 2162 18058
rect 2162 18006 2214 18058
rect 2214 18006 2216 18058
rect 2160 18004 2216 18006
rect 2264 18058 2320 18060
rect 2264 18006 2266 18058
rect 2266 18006 2318 18058
rect 2318 18006 2320 18058
rect 2264 18004 2320 18006
rect 2368 18058 2424 18060
rect 2368 18006 2370 18058
rect 2370 18006 2422 18058
rect 2422 18006 2424 18058
rect 2368 18004 2424 18006
rect 2472 18058 2528 18060
rect 2472 18006 2474 18058
rect 2474 18006 2526 18058
rect 2526 18006 2528 18058
rect 2472 18004 2528 18006
rect 2576 18058 2632 18060
rect 2576 18006 2578 18058
rect 2578 18006 2630 18058
rect 2630 18006 2632 18058
rect 2576 18004 2632 18006
rect 2056 16490 2112 16492
rect 2056 16438 2058 16490
rect 2058 16438 2110 16490
rect 2110 16438 2112 16490
rect 2056 16436 2112 16438
rect 2160 16490 2216 16492
rect 2160 16438 2162 16490
rect 2162 16438 2214 16490
rect 2214 16438 2216 16490
rect 2160 16436 2216 16438
rect 2264 16490 2320 16492
rect 2264 16438 2266 16490
rect 2266 16438 2318 16490
rect 2318 16438 2320 16490
rect 2264 16436 2320 16438
rect 2368 16490 2424 16492
rect 2368 16438 2370 16490
rect 2370 16438 2422 16490
rect 2422 16438 2424 16490
rect 2368 16436 2424 16438
rect 2472 16490 2528 16492
rect 2472 16438 2474 16490
rect 2474 16438 2526 16490
rect 2526 16438 2528 16490
rect 2472 16436 2528 16438
rect 2576 16490 2632 16492
rect 2576 16438 2578 16490
rect 2578 16438 2630 16490
rect 2630 16438 2632 16490
rect 2576 16436 2632 16438
rect 1820 15596 1876 15652
rect 2056 14922 2112 14924
rect 2056 14870 2058 14922
rect 2058 14870 2110 14922
rect 2110 14870 2112 14922
rect 2056 14868 2112 14870
rect 2160 14922 2216 14924
rect 2160 14870 2162 14922
rect 2162 14870 2214 14922
rect 2214 14870 2216 14922
rect 2160 14868 2216 14870
rect 2264 14922 2320 14924
rect 2264 14870 2266 14922
rect 2266 14870 2318 14922
rect 2318 14870 2320 14922
rect 2264 14868 2320 14870
rect 2368 14922 2424 14924
rect 2368 14870 2370 14922
rect 2370 14870 2422 14922
rect 2422 14870 2424 14922
rect 2368 14868 2424 14870
rect 2472 14922 2528 14924
rect 2472 14870 2474 14922
rect 2474 14870 2526 14922
rect 2526 14870 2528 14922
rect 2472 14868 2528 14870
rect 2576 14922 2632 14924
rect 2576 14870 2578 14922
rect 2578 14870 2630 14922
rect 2630 14870 2632 14922
rect 2576 14868 2632 14870
rect 2056 13354 2112 13356
rect 2056 13302 2058 13354
rect 2058 13302 2110 13354
rect 2110 13302 2112 13354
rect 2056 13300 2112 13302
rect 2160 13354 2216 13356
rect 2160 13302 2162 13354
rect 2162 13302 2214 13354
rect 2214 13302 2216 13354
rect 2160 13300 2216 13302
rect 2264 13354 2320 13356
rect 2264 13302 2266 13354
rect 2266 13302 2318 13354
rect 2318 13302 2320 13354
rect 2264 13300 2320 13302
rect 2368 13354 2424 13356
rect 2368 13302 2370 13354
rect 2370 13302 2422 13354
rect 2422 13302 2424 13354
rect 2368 13300 2424 13302
rect 2472 13354 2528 13356
rect 2472 13302 2474 13354
rect 2474 13302 2526 13354
rect 2526 13302 2528 13354
rect 2472 13300 2528 13302
rect 2576 13354 2632 13356
rect 2576 13302 2578 13354
rect 2578 13302 2630 13354
rect 2630 13302 2632 13354
rect 2576 13300 2632 13302
rect 2056 11786 2112 11788
rect 2056 11734 2058 11786
rect 2058 11734 2110 11786
rect 2110 11734 2112 11786
rect 2056 11732 2112 11734
rect 2160 11786 2216 11788
rect 2160 11734 2162 11786
rect 2162 11734 2214 11786
rect 2214 11734 2216 11786
rect 2160 11732 2216 11734
rect 2264 11786 2320 11788
rect 2264 11734 2266 11786
rect 2266 11734 2318 11786
rect 2318 11734 2320 11786
rect 2264 11732 2320 11734
rect 2368 11786 2424 11788
rect 2368 11734 2370 11786
rect 2370 11734 2422 11786
rect 2422 11734 2424 11786
rect 2368 11732 2424 11734
rect 2472 11786 2528 11788
rect 2472 11734 2474 11786
rect 2474 11734 2526 11786
rect 2526 11734 2528 11786
rect 2472 11732 2528 11734
rect 2576 11786 2632 11788
rect 2576 11734 2578 11786
rect 2578 11734 2630 11786
rect 2630 11734 2632 11786
rect 2576 11732 2632 11734
rect 5776 28250 5832 28252
rect 5776 28198 5778 28250
rect 5778 28198 5830 28250
rect 5830 28198 5832 28250
rect 5776 28196 5832 28198
rect 5880 28250 5936 28252
rect 5880 28198 5882 28250
rect 5882 28198 5934 28250
rect 5934 28198 5936 28250
rect 5880 28196 5936 28198
rect 5984 28250 6040 28252
rect 5984 28198 5986 28250
rect 5986 28198 6038 28250
rect 6038 28198 6040 28250
rect 5984 28196 6040 28198
rect 6088 28250 6144 28252
rect 6088 28198 6090 28250
rect 6090 28198 6142 28250
rect 6142 28198 6144 28250
rect 6088 28196 6144 28198
rect 6192 28250 6248 28252
rect 6192 28198 6194 28250
rect 6194 28198 6246 28250
rect 6246 28198 6248 28250
rect 6192 28196 6248 28198
rect 6296 28250 6352 28252
rect 6296 28198 6298 28250
rect 6298 28198 6350 28250
rect 6350 28198 6352 28250
rect 6296 28196 6352 28198
rect 5776 26682 5832 26684
rect 5776 26630 5778 26682
rect 5778 26630 5830 26682
rect 5830 26630 5832 26682
rect 5776 26628 5832 26630
rect 5880 26682 5936 26684
rect 5880 26630 5882 26682
rect 5882 26630 5934 26682
rect 5934 26630 5936 26682
rect 5880 26628 5936 26630
rect 5984 26682 6040 26684
rect 5984 26630 5986 26682
rect 5986 26630 6038 26682
rect 6038 26630 6040 26682
rect 5984 26628 6040 26630
rect 6088 26682 6144 26684
rect 6088 26630 6090 26682
rect 6090 26630 6142 26682
rect 6142 26630 6144 26682
rect 6088 26628 6144 26630
rect 6192 26682 6248 26684
rect 6192 26630 6194 26682
rect 6194 26630 6246 26682
rect 6246 26630 6248 26682
rect 6192 26628 6248 26630
rect 6296 26682 6352 26684
rect 6296 26630 6298 26682
rect 6298 26630 6350 26682
rect 6350 26630 6352 26682
rect 6296 26628 6352 26630
rect 5776 25114 5832 25116
rect 5776 25062 5778 25114
rect 5778 25062 5830 25114
rect 5830 25062 5832 25114
rect 5776 25060 5832 25062
rect 5880 25114 5936 25116
rect 5880 25062 5882 25114
rect 5882 25062 5934 25114
rect 5934 25062 5936 25114
rect 5880 25060 5936 25062
rect 5984 25114 6040 25116
rect 5984 25062 5986 25114
rect 5986 25062 6038 25114
rect 6038 25062 6040 25114
rect 5984 25060 6040 25062
rect 6088 25114 6144 25116
rect 6088 25062 6090 25114
rect 6090 25062 6142 25114
rect 6142 25062 6144 25114
rect 6088 25060 6144 25062
rect 6192 25114 6248 25116
rect 6192 25062 6194 25114
rect 6194 25062 6246 25114
rect 6246 25062 6248 25114
rect 6192 25060 6248 25062
rect 6296 25114 6352 25116
rect 6296 25062 6298 25114
rect 6298 25062 6350 25114
rect 6350 25062 6352 25114
rect 6296 25060 6352 25062
rect 5776 23546 5832 23548
rect 5776 23494 5778 23546
rect 5778 23494 5830 23546
rect 5830 23494 5832 23546
rect 5776 23492 5832 23494
rect 5880 23546 5936 23548
rect 5880 23494 5882 23546
rect 5882 23494 5934 23546
rect 5934 23494 5936 23546
rect 5880 23492 5936 23494
rect 5984 23546 6040 23548
rect 5984 23494 5986 23546
rect 5986 23494 6038 23546
rect 6038 23494 6040 23546
rect 5984 23492 6040 23494
rect 6088 23546 6144 23548
rect 6088 23494 6090 23546
rect 6090 23494 6142 23546
rect 6142 23494 6144 23546
rect 6088 23492 6144 23494
rect 6192 23546 6248 23548
rect 6192 23494 6194 23546
rect 6194 23494 6246 23546
rect 6246 23494 6248 23546
rect 6192 23492 6248 23494
rect 6296 23546 6352 23548
rect 6296 23494 6298 23546
rect 6298 23494 6350 23546
rect 6350 23494 6352 23546
rect 6296 23492 6352 23494
rect 12908 22204 12964 22260
rect 5776 21978 5832 21980
rect 5776 21926 5778 21978
rect 5778 21926 5830 21978
rect 5830 21926 5832 21978
rect 5776 21924 5832 21926
rect 5880 21978 5936 21980
rect 5880 21926 5882 21978
rect 5882 21926 5934 21978
rect 5934 21926 5936 21978
rect 5880 21924 5936 21926
rect 5984 21978 6040 21980
rect 5984 21926 5986 21978
rect 5986 21926 6038 21978
rect 6038 21926 6040 21978
rect 5984 21924 6040 21926
rect 6088 21978 6144 21980
rect 6088 21926 6090 21978
rect 6090 21926 6142 21978
rect 6142 21926 6144 21978
rect 6088 21924 6144 21926
rect 6192 21978 6248 21980
rect 6192 21926 6194 21978
rect 6194 21926 6246 21978
rect 6246 21926 6248 21978
rect 6192 21924 6248 21926
rect 6296 21978 6352 21980
rect 6296 21926 6298 21978
rect 6298 21926 6350 21978
rect 6350 21926 6352 21978
rect 6296 21924 6352 21926
rect 5776 20410 5832 20412
rect 5776 20358 5778 20410
rect 5778 20358 5830 20410
rect 5830 20358 5832 20410
rect 5776 20356 5832 20358
rect 5880 20410 5936 20412
rect 5880 20358 5882 20410
rect 5882 20358 5934 20410
rect 5934 20358 5936 20410
rect 5880 20356 5936 20358
rect 5984 20410 6040 20412
rect 5984 20358 5986 20410
rect 5986 20358 6038 20410
rect 6038 20358 6040 20410
rect 5984 20356 6040 20358
rect 6088 20410 6144 20412
rect 6088 20358 6090 20410
rect 6090 20358 6142 20410
rect 6142 20358 6144 20410
rect 6088 20356 6144 20358
rect 6192 20410 6248 20412
rect 6192 20358 6194 20410
rect 6194 20358 6246 20410
rect 6246 20358 6248 20410
rect 6192 20356 6248 20358
rect 6296 20410 6352 20412
rect 6296 20358 6298 20410
rect 6298 20358 6350 20410
rect 6350 20358 6352 20410
rect 6296 20356 6352 20358
rect 5776 18842 5832 18844
rect 5776 18790 5778 18842
rect 5778 18790 5830 18842
rect 5830 18790 5832 18842
rect 5776 18788 5832 18790
rect 5880 18842 5936 18844
rect 5880 18790 5882 18842
rect 5882 18790 5934 18842
rect 5934 18790 5936 18842
rect 5880 18788 5936 18790
rect 5984 18842 6040 18844
rect 5984 18790 5986 18842
rect 5986 18790 6038 18842
rect 6038 18790 6040 18842
rect 5984 18788 6040 18790
rect 6088 18842 6144 18844
rect 6088 18790 6090 18842
rect 6090 18790 6142 18842
rect 6142 18790 6144 18842
rect 6088 18788 6144 18790
rect 6192 18842 6248 18844
rect 6192 18790 6194 18842
rect 6194 18790 6246 18842
rect 6246 18790 6248 18842
rect 6192 18788 6248 18790
rect 6296 18842 6352 18844
rect 6296 18790 6298 18842
rect 6298 18790 6350 18842
rect 6350 18790 6352 18842
rect 6296 18788 6352 18790
rect 5776 17274 5832 17276
rect 5776 17222 5778 17274
rect 5778 17222 5830 17274
rect 5830 17222 5832 17274
rect 5776 17220 5832 17222
rect 5880 17274 5936 17276
rect 5880 17222 5882 17274
rect 5882 17222 5934 17274
rect 5934 17222 5936 17274
rect 5880 17220 5936 17222
rect 5984 17274 6040 17276
rect 5984 17222 5986 17274
rect 5986 17222 6038 17274
rect 6038 17222 6040 17274
rect 5984 17220 6040 17222
rect 6088 17274 6144 17276
rect 6088 17222 6090 17274
rect 6090 17222 6142 17274
rect 6142 17222 6144 17274
rect 6088 17220 6144 17222
rect 6192 17274 6248 17276
rect 6192 17222 6194 17274
rect 6194 17222 6246 17274
rect 6246 17222 6248 17274
rect 6192 17220 6248 17222
rect 6296 17274 6352 17276
rect 6296 17222 6298 17274
rect 6298 17222 6350 17274
rect 6350 17222 6352 17274
rect 6296 17220 6352 17222
rect 5776 15706 5832 15708
rect 5776 15654 5778 15706
rect 5778 15654 5830 15706
rect 5830 15654 5832 15706
rect 5776 15652 5832 15654
rect 5880 15706 5936 15708
rect 5880 15654 5882 15706
rect 5882 15654 5934 15706
rect 5934 15654 5936 15706
rect 5880 15652 5936 15654
rect 5984 15706 6040 15708
rect 5984 15654 5986 15706
rect 5986 15654 6038 15706
rect 6038 15654 6040 15706
rect 5984 15652 6040 15654
rect 6088 15706 6144 15708
rect 6088 15654 6090 15706
rect 6090 15654 6142 15706
rect 6142 15654 6144 15706
rect 6088 15652 6144 15654
rect 6192 15706 6248 15708
rect 6192 15654 6194 15706
rect 6194 15654 6246 15706
rect 6246 15654 6248 15706
rect 6192 15652 6248 15654
rect 6296 15706 6352 15708
rect 6296 15654 6298 15706
rect 6298 15654 6350 15706
rect 6350 15654 6352 15706
rect 6296 15652 6352 15654
rect 5776 14138 5832 14140
rect 5776 14086 5778 14138
rect 5778 14086 5830 14138
rect 5830 14086 5832 14138
rect 5776 14084 5832 14086
rect 5880 14138 5936 14140
rect 5880 14086 5882 14138
rect 5882 14086 5934 14138
rect 5934 14086 5936 14138
rect 5880 14084 5936 14086
rect 5984 14138 6040 14140
rect 5984 14086 5986 14138
rect 5986 14086 6038 14138
rect 6038 14086 6040 14138
rect 5984 14084 6040 14086
rect 6088 14138 6144 14140
rect 6088 14086 6090 14138
rect 6090 14086 6142 14138
rect 6142 14086 6144 14138
rect 6088 14084 6144 14086
rect 6192 14138 6248 14140
rect 6192 14086 6194 14138
rect 6194 14086 6246 14138
rect 6246 14086 6248 14138
rect 6192 14084 6248 14086
rect 6296 14138 6352 14140
rect 6296 14086 6298 14138
rect 6298 14086 6350 14138
rect 6350 14086 6352 14138
rect 6296 14084 6352 14086
rect 5776 12570 5832 12572
rect 5776 12518 5778 12570
rect 5778 12518 5830 12570
rect 5830 12518 5832 12570
rect 5776 12516 5832 12518
rect 5880 12570 5936 12572
rect 5880 12518 5882 12570
rect 5882 12518 5934 12570
rect 5934 12518 5936 12570
rect 5880 12516 5936 12518
rect 5984 12570 6040 12572
rect 5984 12518 5986 12570
rect 5986 12518 6038 12570
rect 6038 12518 6040 12570
rect 5984 12516 6040 12518
rect 6088 12570 6144 12572
rect 6088 12518 6090 12570
rect 6090 12518 6142 12570
rect 6142 12518 6144 12570
rect 6088 12516 6144 12518
rect 6192 12570 6248 12572
rect 6192 12518 6194 12570
rect 6194 12518 6246 12570
rect 6246 12518 6248 12570
rect 6192 12516 6248 12518
rect 6296 12570 6352 12572
rect 6296 12518 6298 12570
rect 6298 12518 6350 12570
rect 6350 12518 6352 12570
rect 6296 12516 6352 12518
rect 5776 11002 5832 11004
rect 5776 10950 5778 11002
rect 5778 10950 5830 11002
rect 5830 10950 5832 11002
rect 5776 10948 5832 10950
rect 5880 11002 5936 11004
rect 5880 10950 5882 11002
rect 5882 10950 5934 11002
rect 5934 10950 5936 11002
rect 5880 10948 5936 10950
rect 5984 11002 6040 11004
rect 5984 10950 5986 11002
rect 5986 10950 6038 11002
rect 6038 10950 6040 11002
rect 5984 10948 6040 10950
rect 6088 11002 6144 11004
rect 6088 10950 6090 11002
rect 6090 10950 6142 11002
rect 6142 10950 6144 11002
rect 6088 10948 6144 10950
rect 6192 11002 6248 11004
rect 6192 10950 6194 11002
rect 6194 10950 6246 11002
rect 6246 10950 6248 11002
rect 6192 10948 6248 10950
rect 6296 11002 6352 11004
rect 6296 10950 6298 11002
rect 6298 10950 6350 11002
rect 6350 10950 6352 11002
rect 6296 10948 6352 10950
rect 2828 10668 2884 10724
rect 4172 10722 4228 10724
rect 4172 10670 4174 10722
rect 4174 10670 4226 10722
rect 4226 10670 4228 10722
rect 4172 10668 4228 10670
rect 2056 10218 2112 10220
rect 2056 10166 2058 10218
rect 2058 10166 2110 10218
rect 2110 10166 2112 10218
rect 2056 10164 2112 10166
rect 2160 10218 2216 10220
rect 2160 10166 2162 10218
rect 2162 10166 2214 10218
rect 2214 10166 2216 10218
rect 2160 10164 2216 10166
rect 2264 10218 2320 10220
rect 2264 10166 2266 10218
rect 2266 10166 2318 10218
rect 2318 10166 2320 10218
rect 2264 10164 2320 10166
rect 2368 10218 2424 10220
rect 2368 10166 2370 10218
rect 2370 10166 2422 10218
rect 2422 10166 2424 10218
rect 2368 10164 2424 10166
rect 2472 10218 2528 10220
rect 2472 10166 2474 10218
rect 2474 10166 2526 10218
rect 2526 10166 2528 10218
rect 2472 10164 2528 10166
rect 2576 10218 2632 10220
rect 2576 10166 2578 10218
rect 2578 10166 2630 10218
rect 2630 10166 2632 10218
rect 2576 10164 2632 10166
rect 2156 9548 2212 9604
rect 1820 9436 1876 9492
rect 2056 8650 2112 8652
rect 2056 8598 2058 8650
rect 2058 8598 2110 8650
rect 2110 8598 2112 8650
rect 2056 8596 2112 8598
rect 2160 8650 2216 8652
rect 2160 8598 2162 8650
rect 2162 8598 2214 8650
rect 2214 8598 2216 8650
rect 2160 8596 2216 8598
rect 2264 8650 2320 8652
rect 2264 8598 2266 8650
rect 2266 8598 2318 8650
rect 2318 8598 2320 8650
rect 2264 8596 2320 8598
rect 2368 8650 2424 8652
rect 2368 8598 2370 8650
rect 2370 8598 2422 8650
rect 2422 8598 2424 8650
rect 2368 8596 2424 8598
rect 2472 8650 2528 8652
rect 2472 8598 2474 8650
rect 2474 8598 2526 8650
rect 2526 8598 2528 8650
rect 2472 8596 2528 8598
rect 2576 8650 2632 8652
rect 2576 8598 2578 8650
rect 2578 8598 2630 8650
rect 2630 8598 2632 8650
rect 2576 8596 2632 8598
rect 2044 8092 2100 8148
rect 2056 7082 2112 7084
rect 2056 7030 2058 7082
rect 2058 7030 2110 7082
rect 2110 7030 2112 7082
rect 2056 7028 2112 7030
rect 2160 7082 2216 7084
rect 2160 7030 2162 7082
rect 2162 7030 2214 7082
rect 2214 7030 2216 7082
rect 2160 7028 2216 7030
rect 2264 7082 2320 7084
rect 2264 7030 2266 7082
rect 2266 7030 2318 7082
rect 2318 7030 2320 7082
rect 2264 7028 2320 7030
rect 2368 7082 2424 7084
rect 2368 7030 2370 7082
rect 2370 7030 2422 7082
rect 2422 7030 2424 7082
rect 2368 7028 2424 7030
rect 2472 7082 2528 7084
rect 2472 7030 2474 7082
rect 2474 7030 2526 7082
rect 2526 7030 2528 7082
rect 2472 7028 2528 7030
rect 2576 7082 2632 7084
rect 2576 7030 2578 7082
rect 2578 7030 2630 7082
rect 2630 7030 2632 7082
rect 2576 7028 2632 7030
rect 2056 5514 2112 5516
rect 2056 5462 2058 5514
rect 2058 5462 2110 5514
rect 2110 5462 2112 5514
rect 2056 5460 2112 5462
rect 2160 5514 2216 5516
rect 2160 5462 2162 5514
rect 2162 5462 2214 5514
rect 2214 5462 2216 5514
rect 2160 5460 2216 5462
rect 2264 5514 2320 5516
rect 2264 5462 2266 5514
rect 2266 5462 2318 5514
rect 2318 5462 2320 5514
rect 2264 5460 2320 5462
rect 2368 5514 2424 5516
rect 2368 5462 2370 5514
rect 2370 5462 2422 5514
rect 2422 5462 2424 5514
rect 2368 5460 2424 5462
rect 2472 5514 2528 5516
rect 2472 5462 2474 5514
rect 2474 5462 2526 5514
rect 2526 5462 2528 5514
rect 2472 5460 2528 5462
rect 2576 5514 2632 5516
rect 2576 5462 2578 5514
rect 2578 5462 2630 5514
rect 2630 5462 2632 5514
rect 2576 5460 2632 5462
rect 2056 3946 2112 3948
rect 2056 3894 2058 3946
rect 2058 3894 2110 3946
rect 2110 3894 2112 3946
rect 2056 3892 2112 3894
rect 2160 3946 2216 3948
rect 2160 3894 2162 3946
rect 2162 3894 2214 3946
rect 2214 3894 2216 3946
rect 2160 3892 2216 3894
rect 2264 3946 2320 3948
rect 2264 3894 2266 3946
rect 2266 3894 2318 3946
rect 2318 3894 2320 3946
rect 2264 3892 2320 3894
rect 2368 3946 2424 3948
rect 2368 3894 2370 3946
rect 2370 3894 2422 3946
rect 2422 3894 2424 3946
rect 2368 3892 2424 3894
rect 2472 3946 2528 3948
rect 2472 3894 2474 3946
rect 2474 3894 2526 3946
rect 2526 3894 2528 3946
rect 2472 3892 2528 3894
rect 2576 3946 2632 3948
rect 2576 3894 2578 3946
rect 2578 3894 2630 3946
rect 2630 3894 2632 3946
rect 2576 3892 2632 3894
rect 1820 3554 1876 3556
rect 1820 3502 1822 3554
rect 1822 3502 1874 3554
rect 1874 3502 1876 3554
rect 1820 3500 1876 3502
rect 2940 9100 2996 9156
rect 3612 9548 3668 9604
rect 3052 8988 3108 9044
rect 4284 9154 4340 9156
rect 4284 9102 4286 9154
rect 4286 9102 4338 9154
rect 4338 9102 4340 9154
rect 4284 9100 4340 9102
rect 5628 9602 5684 9604
rect 5628 9550 5630 9602
rect 5630 9550 5682 9602
rect 5682 9550 5684 9602
rect 5628 9548 5684 9550
rect 5776 9434 5832 9436
rect 5776 9382 5778 9434
rect 5778 9382 5830 9434
rect 5830 9382 5832 9434
rect 5776 9380 5832 9382
rect 5880 9434 5936 9436
rect 5880 9382 5882 9434
rect 5882 9382 5934 9434
rect 5934 9382 5936 9434
rect 5880 9380 5936 9382
rect 5984 9434 6040 9436
rect 5984 9382 5986 9434
rect 5986 9382 6038 9434
rect 6038 9382 6040 9434
rect 5984 9380 6040 9382
rect 6088 9434 6144 9436
rect 6088 9382 6090 9434
rect 6090 9382 6142 9434
rect 6142 9382 6144 9434
rect 6088 9380 6144 9382
rect 6192 9434 6248 9436
rect 6192 9382 6194 9434
rect 6194 9382 6246 9434
rect 6246 9382 6248 9434
rect 6192 9380 6248 9382
rect 6296 9434 6352 9436
rect 6296 9382 6298 9434
rect 6298 9382 6350 9434
rect 6350 9382 6352 9434
rect 6296 9380 6352 9382
rect 4956 8258 5012 8260
rect 4956 8206 4958 8258
rect 4958 8206 5010 8258
rect 5010 8206 5012 8258
rect 4956 8204 5012 8206
rect 5628 8204 5684 8260
rect 5180 7362 5236 7364
rect 5180 7310 5182 7362
rect 5182 7310 5234 7362
rect 5234 7310 5236 7362
rect 5180 7308 5236 7310
rect 5776 7866 5832 7868
rect 5776 7814 5778 7866
rect 5778 7814 5830 7866
rect 5830 7814 5832 7866
rect 5776 7812 5832 7814
rect 5880 7866 5936 7868
rect 5880 7814 5882 7866
rect 5882 7814 5934 7866
rect 5934 7814 5936 7866
rect 5880 7812 5936 7814
rect 5984 7866 6040 7868
rect 5984 7814 5986 7866
rect 5986 7814 6038 7866
rect 6038 7814 6040 7866
rect 5984 7812 6040 7814
rect 6088 7866 6144 7868
rect 6088 7814 6090 7866
rect 6090 7814 6142 7866
rect 6142 7814 6144 7866
rect 6088 7812 6144 7814
rect 6192 7866 6248 7868
rect 6192 7814 6194 7866
rect 6194 7814 6246 7866
rect 6246 7814 6248 7866
rect 6192 7812 6248 7814
rect 6296 7866 6352 7868
rect 6296 7814 6298 7866
rect 6298 7814 6350 7866
rect 6350 7814 6352 7866
rect 6296 7812 6352 7814
rect 6860 9548 6916 9604
rect 6860 8930 6916 8932
rect 6860 8878 6862 8930
rect 6862 8878 6914 8930
rect 6914 8878 6916 8930
rect 6860 8876 6916 8878
rect 8652 8370 8708 8372
rect 8652 8318 8654 8370
rect 8654 8318 8706 8370
rect 8706 8318 8708 8370
rect 8652 8316 8708 8318
rect 11788 8930 11844 8932
rect 11788 8878 11790 8930
rect 11790 8878 11842 8930
rect 11842 8878 11844 8930
rect 11788 8876 11844 8878
rect 12572 8876 12628 8932
rect 8988 8204 9044 8260
rect 9660 8204 9716 8260
rect 9548 8146 9604 8148
rect 9548 8094 9550 8146
rect 9550 8094 9602 8146
rect 9602 8094 9604 8146
rect 9548 8092 9604 8094
rect 9996 8258 10052 8260
rect 9996 8206 9998 8258
rect 9998 8206 10050 8258
rect 10050 8206 10052 8258
rect 9996 8204 10052 8206
rect 10780 8146 10836 8148
rect 10780 8094 10782 8146
rect 10782 8094 10834 8146
rect 10834 8094 10836 8146
rect 10780 8092 10836 8094
rect 6412 7532 6468 7588
rect 6860 7586 6916 7588
rect 6860 7534 6862 7586
rect 6862 7534 6914 7586
rect 6914 7534 6916 7586
rect 6860 7532 6916 7534
rect 5628 7308 5684 7364
rect 6188 7308 6244 7364
rect 5776 6298 5832 6300
rect 5776 6246 5778 6298
rect 5778 6246 5830 6298
rect 5830 6246 5832 6298
rect 5776 6244 5832 6246
rect 5880 6298 5936 6300
rect 5880 6246 5882 6298
rect 5882 6246 5934 6298
rect 5934 6246 5936 6298
rect 5880 6244 5936 6246
rect 5984 6298 6040 6300
rect 5984 6246 5986 6298
rect 5986 6246 6038 6298
rect 6038 6246 6040 6298
rect 5984 6244 6040 6246
rect 6088 6298 6144 6300
rect 6088 6246 6090 6298
rect 6090 6246 6142 6298
rect 6142 6246 6144 6298
rect 6088 6244 6144 6246
rect 6192 6298 6248 6300
rect 6192 6246 6194 6298
rect 6194 6246 6246 6298
rect 6246 6246 6248 6298
rect 6192 6244 6248 6246
rect 6296 6298 6352 6300
rect 6296 6246 6298 6298
rect 6298 6246 6350 6298
rect 6350 6246 6352 6298
rect 6296 6244 6352 6246
rect 9660 7308 9716 7364
rect 11788 7362 11844 7364
rect 11788 7310 11790 7362
rect 11790 7310 11842 7362
rect 11842 7310 11844 7362
rect 11788 7308 11844 7310
rect 16380 22092 16436 22148
rect 14476 18956 14532 19012
rect 13468 9884 13524 9940
rect 13468 8876 13524 8932
rect 13020 8316 13076 8372
rect 13580 8034 13636 8036
rect 13580 7982 13582 8034
rect 13582 7982 13634 8034
rect 13634 7982 13636 8034
rect 13580 7980 13636 7982
rect 13580 7308 13636 7364
rect 13020 6690 13076 6692
rect 13020 6638 13022 6690
rect 13022 6638 13074 6690
rect 13074 6638 13076 6690
rect 13020 6636 13076 6638
rect 12684 6076 12740 6132
rect 15484 16828 15540 16884
rect 14812 10722 14868 10724
rect 14812 10670 14814 10722
rect 14814 10670 14866 10722
rect 14866 10670 14868 10722
rect 14812 10668 14868 10670
rect 14476 6690 14532 6692
rect 14476 6638 14478 6690
rect 14478 6638 14530 6690
rect 14530 6638 14532 6690
rect 14476 6636 14532 6638
rect 13804 6076 13860 6132
rect 13356 6018 13412 6020
rect 13356 5966 13358 6018
rect 13358 5966 13410 6018
rect 13410 5966 13412 6018
rect 13356 5964 13412 5966
rect 15596 9884 15652 9940
rect 16044 9938 16100 9940
rect 16044 9886 16046 9938
rect 16046 9886 16098 9938
rect 16098 9886 16100 9938
rect 16044 9884 16100 9886
rect 15932 6130 15988 6132
rect 15932 6078 15934 6130
rect 15934 6078 15986 6130
rect 15986 6078 15988 6130
rect 15932 6076 15988 6078
rect 38056 35306 38112 35308
rect 38056 35254 38058 35306
rect 38058 35254 38110 35306
rect 38110 35254 38112 35306
rect 38056 35252 38112 35254
rect 38160 35306 38216 35308
rect 38160 35254 38162 35306
rect 38162 35254 38214 35306
rect 38214 35254 38216 35306
rect 38160 35252 38216 35254
rect 38264 35306 38320 35308
rect 38264 35254 38266 35306
rect 38266 35254 38318 35306
rect 38318 35254 38320 35306
rect 38264 35252 38320 35254
rect 38368 35306 38424 35308
rect 38368 35254 38370 35306
rect 38370 35254 38422 35306
rect 38422 35254 38424 35306
rect 38368 35252 38424 35254
rect 38472 35306 38528 35308
rect 38472 35254 38474 35306
rect 38474 35254 38526 35306
rect 38526 35254 38528 35306
rect 38472 35252 38528 35254
rect 38576 35306 38632 35308
rect 38576 35254 38578 35306
rect 38578 35254 38630 35306
rect 38630 35254 38632 35306
rect 38576 35252 38632 35254
rect 38056 33738 38112 33740
rect 38056 33686 38058 33738
rect 38058 33686 38110 33738
rect 38110 33686 38112 33738
rect 38056 33684 38112 33686
rect 38160 33738 38216 33740
rect 38160 33686 38162 33738
rect 38162 33686 38214 33738
rect 38214 33686 38216 33738
rect 38160 33684 38216 33686
rect 38264 33738 38320 33740
rect 38264 33686 38266 33738
rect 38266 33686 38318 33738
rect 38318 33686 38320 33738
rect 38264 33684 38320 33686
rect 38368 33738 38424 33740
rect 38368 33686 38370 33738
rect 38370 33686 38422 33738
rect 38422 33686 38424 33738
rect 38368 33684 38424 33686
rect 38472 33738 38528 33740
rect 38472 33686 38474 33738
rect 38474 33686 38526 33738
rect 38526 33686 38528 33738
rect 38472 33684 38528 33686
rect 38576 33738 38632 33740
rect 38576 33686 38578 33738
rect 38578 33686 38630 33738
rect 38630 33686 38632 33738
rect 38576 33684 38632 33686
rect 38056 32170 38112 32172
rect 38056 32118 38058 32170
rect 38058 32118 38110 32170
rect 38110 32118 38112 32170
rect 38056 32116 38112 32118
rect 38160 32170 38216 32172
rect 38160 32118 38162 32170
rect 38162 32118 38214 32170
rect 38214 32118 38216 32170
rect 38160 32116 38216 32118
rect 38264 32170 38320 32172
rect 38264 32118 38266 32170
rect 38266 32118 38318 32170
rect 38318 32118 38320 32170
rect 38264 32116 38320 32118
rect 38368 32170 38424 32172
rect 38368 32118 38370 32170
rect 38370 32118 38422 32170
rect 38422 32118 38424 32170
rect 38368 32116 38424 32118
rect 38472 32170 38528 32172
rect 38472 32118 38474 32170
rect 38474 32118 38526 32170
rect 38526 32118 38528 32170
rect 38472 32116 38528 32118
rect 38576 32170 38632 32172
rect 38576 32118 38578 32170
rect 38578 32118 38630 32170
rect 38630 32118 38632 32170
rect 38576 32116 38632 32118
rect 38056 30602 38112 30604
rect 38056 30550 38058 30602
rect 38058 30550 38110 30602
rect 38110 30550 38112 30602
rect 38056 30548 38112 30550
rect 38160 30602 38216 30604
rect 38160 30550 38162 30602
rect 38162 30550 38214 30602
rect 38214 30550 38216 30602
rect 38160 30548 38216 30550
rect 38264 30602 38320 30604
rect 38264 30550 38266 30602
rect 38266 30550 38318 30602
rect 38318 30550 38320 30602
rect 38264 30548 38320 30550
rect 38368 30602 38424 30604
rect 38368 30550 38370 30602
rect 38370 30550 38422 30602
rect 38422 30550 38424 30602
rect 38368 30548 38424 30550
rect 38472 30602 38528 30604
rect 38472 30550 38474 30602
rect 38474 30550 38526 30602
rect 38526 30550 38528 30602
rect 38472 30548 38528 30550
rect 38576 30602 38632 30604
rect 38576 30550 38578 30602
rect 38578 30550 38630 30602
rect 38630 30550 38632 30602
rect 38576 30548 38632 30550
rect 39004 29538 39060 29540
rect 39004 29486 39006 29538
rect 39006 29486 39058 29538
rect 39058 29486 39060 29538
rect 39004 29484 39060 29486
rect 32956 28700 33012 28756
rect 30380 28588 30436 28644
rect 29484 27916 29540 27972
rect 27916 25340 27972 25396
rect 17388 20524 17444 20580
rect 20524 21420 20580 21476
rect 17388 16828 17444 16884
rect 19740 19292 19796 19348
rect 19068 13074 19124 13076
rect 19068 13022 19070 13074
rect 19070 13022 19122 13074
rect 19122 13022 19124 13074
rect 19068 13020 19124 13022
rect 16940 12850 16996 12852
rect 16940 12798 16942 12850
rect 16942 12798 16994 12850
rect 16994 12798 16996 12850
rect 16940 12796 16996 12798
rect 19628 12850 19684 12852
rect 19628 12798 19630 12850
rect 19630 12798 19682 12850
rect 19682 12798 19684 12850
rect 19628 12796 19684 12798
rect 18396 12348 18452 12404
rect 16940 11004 16996 11060
rect 16604 9884 16660 9940
rect 17612 10722 17668 10724
rect 17612 10670 17614 10722
rect 17614 10670 17666 10722
rect 17666 10670 17668 10722
rect 17612 10668 17668 10670
rect 17052 9884 17108 9940
rect 22428 21308 22484 21364
rect 20860 18284 20916 18340
rect 20748 12402 20804 12404
rect 20748 12350 20750 12402
rect 20750 12350 20802 12402
rect 20802 12350 20804 12402
rect 20748 12348 20804 12350
rect 20300 10780 20356 10836
rect 18956 9884 19012 9940
rect 17388 9714 17444 9716
rect 17388 9662 17390 9714
rect 17390 9662 17442 9714
rect 17442 9662 17444 9714
rect 17388 9660 17444 9662
rect 20076 9714 20132 9716
rect 20076 9662 20078 9714
rect 20078 9662 20130 9714
rect 20130 9662 20132 9714
rect 20076 9660 20132 9662
rect 19964 9212 20020 9268
rect 19180 9042 19236 9044
rect 19180 8990 19182 9042
rect 19182 8990 19234 9042
rect 19234 8990 19236 9042
rect 19180 8988 19236 8990
rect 19628 9042 19684 9044
rect 19628 8990 19630 9042
rect 19630 8990 19682 9042
rect 19682 8990 19684 9042
rect 19628 8988 19684 8990
rect 16716 8876 16772 8932
rect 16492 8034 16548 8036
rect 16492 7982 16494 8034
rect 16494 7982 16546 8034
rect 16546 7982 16548 8034
rect 16492 7980 16548 7982
rect 17724 8930 17780 8932
rect 17724 8878 17726 8930
rect 17726 8878 17778 8930
rect 17778 8878 17780 8930
rect 17724 8876 17780 8878
rect 17052 7980 17108 8036
rect 17388 7980 17444 8036
rect 16604 6636 16660 6692
rect 17836 7980 17892 8036
rect 20524 8034 20580 8036
rect 20524 7982 20526 8034
rect 20526 7982 20578 8034
rect 20578 7982 20580 8034
rect 20524 7980 20580 7982
rect 20300 6860 20356 6916
rect 17388 6802 17444 6804
rect 17388 6750 17390 6802
rect 17390 6750 17442 6802
rect 17442 6750 17444 6802
rect 17388 6748 17444 6750
rect 16380 5964 16436 6020
rect 8988 5180 9044 5236
rect 17948 6748 18004 6804
rect 18732 6578 18788 6580
rect 18732 6526 18734 6578
rect 18734 6526 18786 6578
rect 18786 6526 18788 6578
rect 18732 6524 18788 6526
rect 16940 5234 16996 5236
rect 16940 5182 16942 5234
rect 16942 5182 16994 5234
rect 16994 5182 16996 5234
rect 16940 5180 16996 5182
rect 18172 5234 18228 5236
rect 18172 5182 18174 5234
rect 18174 5182 18226 5234
rect 18226 5182 18228 5234
rect 18172 5180 18228 5182
rect 21644 11506 21700 11508
rect 21644 11454 21646 11506
rect 21646 11454 21698 11506
rect 21698 11454 21700 11506
rect 21644 11452 21700 11454
rect 22652 20188 22708 20244
rect 21644 9996 21700 10052
rect 25676 19852 25732 19908
rect 23660 19740 23716 19796
rect 23660 13020 23716 13076
rect 23772 15820 23828 15876
rect 25004 15596 25060 15652
rect 24556 11394 24612 11396
rect 24556 11342 24558 11394
rect 24558 11342 24610 11394
rect 24610 11342 24612 11394
rect 24556 11340 24612 11342
rect 24780 11340 24836 11396
rect 22876 10834 22932 10836
rect 22876 10782 22878 10834
rect 22878 10782 22930 10834
rect 22930 10782 22932 10834
rect 22876 10780 22932 10782
rect 22652 9996 22708 10052
rect 28028 22146 28084 22148
rect 28028 22094 28030 22146
rect 28030 22094 28082 22146
rect 28082 22094 28084 22146
rect 28028 22092 28084 22094
rect 28028 21868 28084 21924
rect 27132 15874 27188 15876
rect 27132 15822 27134 15874
rect 27134 15822 27186 15874
rect 27186 15822 27188 15874
rect 27132 15820 27188 15822
rect 25676 11452 25732 11508
rect 25900 11506 25956 11508
rect 25900 11454 25902 11506
rect 25902 11454 25954 11506
rect 25954 11454 25956 11506
rect 25900 11452 25956 11454
rect 25116 11394 25172 11396
rect 25116 11342 25118 11394
rect 25118 11342 25170 11394
rect 25170 11342 25172 11394
rect 25116 11340 25172 11342
rect 27468 11340 27524 11396
rect 28364 20972 28420 21028
rect 28812 20578 28868 20580
rect 28812 20526 28814 20578
rect 28814 20526 28866 20578
rect 28866 20526 28868 20578
rect 28812 20524 28868 20526
rect 29372 20130 29428 20132
rect 29372 20078 29374 20130
rect 29374 20078 29426 20130
rect 29426 20078 29428 20130
rect 29372 20076 29428 20078
rect 30044 26012 30100 26068
rect 29820 21026 29876 21028
rect 29820 20974 29822 21026
rect 29822 20974 29874 21026
rect 29874 20974 29876 21026
rect 29820 20972 29876 20974
rect 30156 20524 30212 20580
rect 28476 16044 28532 16100
rect 28252 15820 28308 15876
rect 27916 11340 27972 11396
rect 28924 15708 28980 15764
rect 28812 13692 28868 13748
rect 28364 11340 28420 11396
rect 25004 9212 25060 9268
rect 23436 8930 23492 8932
rect 23436 8878 23438 8930
rect 23438 8878 23490 8930
rect 23490 8878 23492 8930
rect 23436 8876 23492 8878
rect 23436 7420 23492 7476
rect 24444 7420 24500 7476
rect 21644 6578 21700 6580
rect 21644 6526 21646 6578
rect 21646 6526 21698 6578
rect 21698 6526 21700 6578
rect 21644 6524 21700 6526
rect 22876 7196 22932 7252
rect 22876 5180 22932 5236
rect 26236 7474 26292 7476
rect 26236 7422 26238 7474
rect 26238 7422 26290 7474
rect 26290 7422 26292 7474
rect 26236 7420 26292 7422
rect 28252 7474 28308 7476
rect 28252 7422 28254 7474
rect 28254 7422 28306 7474
rect 28306 7422 28308 7474
rect 28252 7420 28308 7422
rect 26684 6578 26740 6580
rect 26684 6526 26686 6578
rect 26686 6526 26738 6578
rect 26738 6526 26740 6578
rect 26684 6524 26740 6526
rect 26460 5906 26516 5908
rect 26460 5854 26462 5906
rect 26462 5854 26514 5906
rect 26514 5854 26516 5906
rect 26460 5852 26516 5854
rect 26012 4956 26068 5012
rect 5776 4730 5832 4732
rect 5776 4678 5778 4730
rect 5778 4678 5830 4730
rect 5830 4678 5832 4730
rect 5776 4676 5832 4678
rect 5880 4730 5936 4732
rect 5880 4678 5882 4730
rect 5882 4678 5934 4730
rect 5934 4678 5936 4730
rect 5880 4676 5936 4678
rect 5984 4730 6040 4732
rect 5984 4678 5986 4730
rect 5986 4678 6038 4730
rect 6038 4678 6040 4730
rect 5984 4676 6040 4678
rect 6088 4730 6144 4732
rect 6088 4678 6090 4730
rect 6090 4678 6142 4730
rect 6142 4678 6144 4730
rect 6088 4676 6144 4678
rect 6192 4730 6248 4732
rect 6192 4678 6194 4730
rect 6194 4678 6246 4730
rect 6246 4678 6248 4730
rect 6192 4676 6248 4678
rect 6296 4730 6352 4732
rect 6296 4678 6298 4730
rect 6298 4678 6350 4730
rect 6350 4678 6352 4730
rect 6296 4676 6352 4678
rect 22540 4620 22596 4676
rect 20412 4396 20468 4452
rect 24220 4620 24276 4676
rect 23324 4338 23380 4340
rect 23324 4286 23326 4338
rect 23326 4286 23378 4338
rect 23378 4286 23380 4338
rect 23324 4284 23380 4286
rect 23772 4338 23828 4340
rect 23772 4286 23774 4338
rect 23774 4286 23826 4338
rect 23826 4286 23828 4338
rect 23772 4284 23828 4286
rect 28028 5010 28084 5012
rect 28028 4958 28030 5010
rect 28030 4958 28082 5010
rect 28082 4958 28084 5010
rect 28028 4956 28084 4958
rect 26460 4508 26516 4564
rect 25676 4284 25732 4340
rect 28588 11506 28644 11508
rect 28588 11454 28590 11506
rect 28590 11454 28642 11506
rect 28642 11454 28644 11506
rect 28588 11452 28644 11454
rect 29148 15426 29204 15428
rect 29148 15374 29150 15426
rect 29150 15374 29202 15426
rect 29202 15374 29204 15426
rect 29148 15372 29204 15374
rect 29708 17666 29764 17668
rect 29708 17614 29710 17666
rect 29710 17614 29762 17666
rect 29762 17614 29764 17666
rect 29708 17612 29764 17614
rect 31500 27804 31556 27860
rect 30828 25228 30884 25284
rect 30380 17612 30436 17668
rect 30492 23324 30548 23380
rect 29932 16268 29988 16324
rect 30380 16268 30436 16324
rect 30044 15372 30100 15428
rect 29484 13468 29540 13524
rect 30044 14588 30100 14644
rect 29596 11394 29652 11396
rect 29596 11342 29598 11394
rect 29598 11342 29650 11394
rect 29650 11342 29652 11394
rect 29596 11340 29652 11342
rect 29932 9772 29988 9828
rect 29148 7420 29204 7476
rect 29036 5906 29092 5908
rect 29036 5854 29038 5906
rect 29038 5854 29090 5906
rect 29090 5854 29092 5906
rect 29036 5852 29092 5854
rect 29596 6578 29652 6580
rect 29596 6526 29598 6578
rect 29598 6526 29650 6578
rect 29650 6526 29652 6578
rect 29596 6524 29652 6526
rect 29260 4956 29316 5012
rect 29484 4956 29540 5012
rect 29708 4956 29764 5012
rect 29932 4956 29988 5012
rect 29708 4562 29764 4564
rect 29708 4510 29710 4562
rect 29710 4510 29762 4562
rect 29762 4510 29764 4562
rect 29708 4508 29764 4510
rect 31612 27692 31668 27748
rect 32396 26124 32452 26180
rect 30828 20076 30884 20132
rect 31836 23100 31892 23156
rect 31276 19122 31332 19124
rect 31276 19070 31278 19122
rect 31278 19070 31330 19122
rect 31330 19070 31332 19122
rect 31276 19068 31332 19070
rect 30940 16380 30996 16436
rect 31276 18562 31332 18564
rect 31276 18510 31278 18562
rect 31278 18510 31330 18562
rect 31330 18510 31332 18562
rect 31276 18508 31332 18510
rect 30492 13468 30548 13524
rect 30380 10556 30436 10612
rect 31052 15874 31108 15876
rect 31052 15822 31054 15874
rect 31054 15822 31106 15874
rect 31106 15822 31108 15874
rect 31052 15820 31108 15822
rect 30940 12684 30996 12740
rect 31052 15484 31108 15540
rect 30828 9772 30884 9828
rect 30716 8930 30772 8932
rect 30716 8878 30718 8930
rect 30718 8878 30770 8930
rect 30770 8878 30772 8930
rect 30716 8876 30772 8878
rect 31164 11452 31220 11508
rect 32172 20524 32228 20580
rect 31612 17724 31668 17780
rect 31500 17052 31556 17108
rect 31388 15986 31444 15988
rect 31388 15934 31390 15986
rect 31390 15934 31442 15986
rect 31442 15934 31444 15986
rect 31388 15932 31444 15934
rect 32060 17778 32116 17780
rect 32060 17726 32062 17778
rect 32062 17726 32114 17778
rect 32114 17726 32116 17778
rect 32060 17724 32116 17726
rect 32060 17106 32116 17108
rect 32060 17054 32062 17106
rect 32062 17054 32114 17106
rect 32114 17054 32116 17106
rect 32060 17052 32116 17054
rect 31836 15932 31892 15988
rect 31836 12348 31892 12404
rect 31836 12124 31892 12180
rect 31276 10780 31332 10836
rect 32284 10668 32340 10724
rect 32620 18284 32676 18340
rect 32844 16098 32900 16100
rect 32844 16046 32846 16098
rect 32846 16046 32898 16098
rect 32898 16046 32900 16098
rect 32844 16044 32900 16046
rect 36764 28754 36820 28756
rect 36764 28702 36766 28754
rect 36766 28702 36818 28754
rect 36818 28702 36820 28754
rect 36764 28700 36820 28702
rect 35196 28028 35252 28084
rect 34636 27580 34692 27636
rect 34636 25340 34692 25396
rect 36652 28082 36708 28084
rect 36652 28030 36654 28082
rect 36654 28030 36706 28082
rect 36706 28030 36708 28082
rect 36652 28028 36708 28030
rect 36204 27746 36260 27748
rect 36204 27694 36206 27746
rect 36206 27694 36258 27746
rect 36258 27694 36260 27746
rect 36204 27692 36260 27694
rect 37660 28028 37716 28084
rect 38056 29034 38112 29036
rect 38056 28982 38058 29034
rect 38058 28982 38110 29034
rect 38110 28982 38112 29034
rect 38056 28980 38112 28982
rect 38160 29034 38216 29036
rect 38160 28982 38162 29034
rect 38162 28982 38214 29034
rect 38214 28982 38216 29034
rect 38160 28980 38216 28982
rect 38264 29034 38320 29036
rect 38264 28982 38266 29034
rect 38266 28982 38318 29034
rect 38318 28982 38320 29034
rect 38264 28980 38320 28982
rect 38368 29034 38424 29036
rect 38368 28982 38370 29034
rect 38370 28982 38422 29034
rect 38422 28982 38424 29034
rect 38368 28980 38424 28982
rect 38472 29034 38528 29036
rect 38472 28982 38474 29034
rect 38474 28982 38526 29034
rect 38526 28982 38528 29034
rect 38472 28980 38528 28982
rect 38576 29034 38632 29036
rect 38576 28982 38578 29034
rect 38578 28982 38630 29034
rect 38630 28982 38632 29034
rect 38576 28980 38632 28982
rect 38332 28754 38388 28756
rect 38332 28702 38334 28754
rect 38334 28702 38386 28754
rect 38386 28702 38388 28754
rect 38332 28700 38388 28702
rect 37996 28642 38052 28644
rect 37996 28590 37998 28642
rect 37998 28590 38050 28642
rect 38050 28590 38052 28642
rect 37996 28588 38052 28590
rect 37884 27916 37940 27972
rect 38220 27970 38276 27972
rect 38220 27918 38222 27970
rect 38222 27918 38274 27970
rect 38274 27918 38276 27970
rect 38220 27916 38276 27918
rect 38108 27858 38164 27860
rect 38108 27806 38110 27858
rect 38110 27806 38162 27858
rect 38162 27806 38164 27858
rect 38108 27804 38164 27806
rect 37436 27692 37492 27748
rect 38556 27804 38612 27860
rect 39004 28588 39060 28644
rect 38780 28476 38836 28532
rect 38780 27804 38836 27860
rect 38220 27692 38276 27748
rect 37324 27634 37380 27636
rect 37324 27582 37326 27634
rect 37326 27582 37378 27634
rect 37378 27582 37380 27634
rect 37324 27580 37380 27582
rect 38056 27466 38112 27468
rect 38056 27414 38058 27466
rect 38058 27414 38110 27466
rect 38110 27414 38112 27466
rect 38056 27412 38112 27414
rect 38160 27466 38216 27468
rect 38160 27414 38162 27466
rect 38162 27414 38214 27466
rect 38214 27414 38216 27466
rect 38160 27412 38216 27414
rect 38264 27466 38320 27468
rect 38264 27414 38266 27466
rect 38266 27414 38318 27466
rect 38318 27414 38320 27466
rect 38264 27412 38320 27414
rect 38368 27466 38424 27468
rect 38368 27414 38370 27466
rect 38370 27414 38422 27466
rect 38422 27414 38424 27466
rect 38368 27412 38424 27414
rect 38472 27466 38528 27468
rect 38472 27414 38474 27466
rect 38474 27414 38526 27466
rect 38526 27414 38528 27466
rect 38472 27412 38528 27414
rect 38576 27466 38632 27468
rect 38576 27414 38578 27466
rect 38578 27414 38630 27466
rect 38630 27414 38632 27466
rect 38576 27412 38632 27414
rect 41776 40794 41832 40796
rect 41776 40742 41778 40794
rect 41778 40742 41830 40794
rect 41830 40742 41832 40794
rect 41776 40740 41832 40742
rect 41880 40794 41936 40796
rect 41880 40742 41882 40794
rect 41882 40742 41934 40794
rect 41934 40742 41936 40794
rect 41880 40740 41936 40742
rect 41984 40794 42040 40796
rect 41984 40742 41986 40794
rect 41986 40742 42038 40794
rect 42038 40742 42040 40794
rect 41984 40740 42040 40742
rect 42088 40794 42144 40796
rect 42088 40742 42090 40794
rect 42090 40742 42142 40794
rect 42142 40742 42144 40794
rect 42088 40740 42144 40742
rect 42192 40794 42248 40796
rect 42192 40742 42194 40794
rect 42194 40742 42246 40794
rect 42246 40742 42248 40794
rect 42192 40740 42248 40742
rect 42296 40794 42352 40796
rect 42296 40742 42298 40794
rect 42298 40742 42350 40794
rect 42350 40742 42352 40794
rect 42296 40740 42352 40742
rect 41776 39226 41832 39228
rect 41776 39174 41778 39226
rect 41778 39174 41830 39226
rect 41830 39174 41832 39226
rect 41776 39172 41832 39174
rect 41880 39226 41936 39228
rect 41880 39174 41882 39226
rect 41882 39174 41934 39226
rect 41934 39174 41936 39226
rect 41880 39172 41936 39174
rect 41984 39226 42040 39228
rect 41984 39174 41986 39226
rect 41986 39174 42038 39226
rect 42038 39174 42040 39226
rect 41984 39172 42040 39174
rect 42088 39226 42144 39228
rect 42088 39174 42090 39226
rect 42090 39174 42142 39226
rect 42142 39174 42144 39226
rect 42088 39172 42144 39174
rect 42192 39226 42248 39228
rect 42192 39174 42194 39226
rect 42194 39174 42246 39226
rect 42246 39174 42248 39226
rect 42192 39172 42248 39174
rect 42296 39226 42352 39228
rect 42296 39174 42298 39226
rect 42298 39174 42350 39226
rect 42350 39174 42352 39226
rect 42296 39172 42352 39174
rect 41132 38668 41188 38724
rect 39788 28476 39844 28532
rect 40124 28530 40180 28532
rect 40124 28478 40126 28530
rect 40126 28478 40178 28530
rect 40178 28478 40180 28530
rect 40124 28476 40180 28478
rect 35196 25228 35252 25284
rect 37100 26348 37156 26404
rect 37548 26178 37604 26180
rect 37548 26126 37550 26178
rect 37550 26126 37602 26178
rect 37602 26126 37604 26178
rect 37548 26124 37604 26126
rect 38556 26178 38612 26180
rect 38556 26126 38558 26178
rect 38558 26126 38610 26178
rect 38610 26126 38612 26178
rect 38556 26124 38612 26126
rect 39116 27858 39172 27860
rect 39116 27806 39118 27858
rect 39118 27806 39170 27858
rect 39170 27806 39172 27858
rect 39116 27804 39172 27806
rect 39116 26402 39172 26404
rect 39116 26350 39118 26402
rect 39118 26350 39170 26402
rect 39170 26350 39172 26402
rect 39116 26348 39172 26350
rect 39788 26796 39844 26852
rect 40236 26850 40292 26852
rect 40236 26798 40238 26850
rect 40238 26798 40290 26850
rect 40290 26798 40292 26850
rect 40236 26796 40292 26798
rect 40796 26796 40852 26852
rect 38892 26124 38948 26180
rect 38220 26066 38276 26068
rect 38220 26014 38222 26066
rect 38222 26014 38274 26066
rect 38274 26014 38276 26066
rect 38220 26012 38276 26014
rect 38056 25898 38112 25900
rect 38056 25846 38058 25898
rect 38058 25846 38110 25898
rect 38110 25846 38112 25898
rect 38056 25844 38112 25846
rect 38160 25898 38216 25900
rect 38160 25846 38162 25898
rect 38162 25846 38214 25898
rect 38214 25846 38216 25898
rect 38160 25844 38216 25846
rect 38264 25898 38320 25900
rect 38264 25846 38266 25898
rect 38266 25846 38318 25898
rect 38318 25846 38320 25898
rect 38264 25844 38320 25846
rect 38368 25898 38424 25900
rect 38368 25846 38370 25898
rect 38370 25846 38422 25898
rect 38422 25846 38424 25898
rect 38368 25844 38424 25846
rect 38472 25898 38528 25900
rect 38472 25846 38474 25898
rect 38474 25846 38526 25898
rect 38526 25846 38528 25898
rect 38472 25844 38528 25846
rect 38576 25898 38632 25900
rect 38576 25846 38578 25898
rect 38578 25846 38630 25898
rect 38630 25846 38632 25898
rect 38576 25844 38632 25846
rect 39116 24834 39172 24836
rect 39116 24782 39118 24834
rect 39118 24782 39170 24834
rect 39170 24782 39172 24834
rect 39116 24780 39172 24782
rect 36988 23884 37044 23940
rect 34972 22092 35028 22148
rect 33404 21756 33460 21812
rect 32620 13468 32676 13524
rect 32508 11676 32564 11732
rect 31836 9772 31892 9828
rect 31052 9660 31108 9716
rect 32732 12124 32788 12180
rect 33292 15708 33348 15764
rect 33292 14700 33348 14756
rect 34300 20636 34356 20692
rect 33628 20242 33684 20244
rect 33628 20190 33630 20242
rect 33630 20190 33682 20242
rect 33682 20190 33684 20242
rect 33628 20188 33684 20190
rect 33516 18620 33572 18676
rect 33516 16044 33572 16100
rect 33740 18844 33796 18900
rect 34188 18956 34244 19012
rect 34300 18844 34356 18900
rect 33964 17948 34020 18004
rect 33964 16828 34020 16884
rect 34860 19010 34916 19012
rect 34860 18958 34862 19010
rect 34862 18958 34914 19010
rect 34914 18958 34916 19010
rect 34860 18956 34916 18958
rect 34748 17836 34804 17892
rect 34860 18450 34916 18452
rect 34860 18398 34862 18450
rect 34862 18398 34914 18450
rect 34914 18398 34916 18450
rect 34860 18396 34916 18398
rect 34300 16940 34356 16996
rect 34188 16044 34244 16100
rect 34300 15708 34356 15764
rect 34300 15484 34356 15540
rect 33740 14700 33796 14756
rect 33404 11676 33460 11732
rect 33180 11228 33236 11284
rect 32956 9938 33012 9940
rect 32956 9886 32958 9938
rect 32958 9886 33010 9938
rect 33010 9886 33012 9938
rect 32956 9884 33012 9886
rect 33516 9938 33572 9940
rect 33516 9886 33518 9938
rect 33518 9886 33570 9938
rect 33570 9886 33572 9938
rect 33516 9884 33572 9886
rect 33516 9324 33572 9380
rect 33516 8876 33572 8932
rect 34412 15260 34468 15316
rect 34860 17612 34916 17668
rect 34300 14700 34356 14756
rect 34076 13634 34132 13636
rect 34076 13582 34078 13634
rect 34078 13582 34130 13634
rect 34130 13582 34132 13634
rect 34076 13580 34132 13582
rect 34860 16828 34916 16884
rect 36428 21474 36484 21476
rect 36428 21422 36430 21474
rect 36430 21422 36482 21474
rect 36482 21422 36484 21474
rect 36428 21420 36484 21422
rect 36876 23212 36932 23268
rect 36764 21420 36820 21476
rect 37324 22876 37380 22932
rect 37324 21868 37380 21924
rect 38056 24330 38112 24332
rect 38056 24278 38058 24330
rect 38058 24278 38110 24330
rect 38110 24278 38112 24330
rect 38056 24276 38112 24278
rect 38160 24330 38216 24332
rect 38160 24278 38162 24330
rect 38162 24278 38214 24330
rect 38214 24278 38216 24330
rect 38160 24276 38216 24278
rect 38264 24330 38320 24332
rect 38264 24278 38266 24330
rect 38266 24278 38318 24330
rect 38318 24278 38320 24330
rect 38264 24276 38320 24278
rect 38368 24330 38424 24332
rect 38368 24278 38370 24330
rect 38370 24278 38422 24330
rect 38422 24278 38424 24330
rect 38368 24276 38424 24278
rect 38472 24330 38528 24332
rect 38472 24278 38474 24330
rect 38474 24278 38526 24330
rect 38526 24278 38528 24330
rect 38472 24276 38528 24278
rect 38576 24330 38632 24332
rect 38576 24278 38578 24330
rect 38578 24278 38630 24330
rect 38630 24278 38632 24330
rect 38576 24276 38632 24278
rect 39116 24108 39172 24164
rect 38332 23938 38388 23940
rect 38332 23886 38334 23938
rect 38334 23886 38386 23938
rect 38386 23886 38388 23938
rect 38332 23884 38388 23886
rect 39676 25228 39732 25284
rect 37884 23324 37940 23380
rect 37996 23100 38052 23156
rect 38332 23436 38388 23492
rect 37436 21756 37492 21812
rect 36876 21308 36932 21364
rect 36764 20972 36820 21028
rect 36428 20188 36484 20244
rect 35980 19740 36036 19796
rect 36428 19292 36484 19348
rect 36764 19740 36820 19796
rect 36764 19404 36820 19460
rect 36204 19010 36260 19012
rect 36204 18958 36206 19010
rect 36206 18958 36258 19010
rect 36258 18958 36260 19010
rect 36204 18956 36260 18958
rect 35756 18732 35812 18788
rect 35084 18396 35140 18452
rect 35644 18450 35700 18452
rect 35644 18398 35646 18450
rect 35646 18398 35698 18450
rect 35698 18398 35700 18450
rect 35644 18396 35700 18398
rect 35420 18060 35476 18116
rect 35532 17948 35588 18004
rect 35420 17836 35476 17892
rect 34748 15708 34804 15764
rect 35308 17500 35364 17556
rect 34860 15484 34916 15540
rect 34972 16044 35028 16100
rect 34748 15260 34804 15316
rect 36764 18732 36820 18788
rect 36652 18396 36708 18452
rect 36428 18338 36484 18340
rect 36428 18286 36430 18338
rect 36430 18286 36482 18338
rect 36482 18286 36484 18338
rect 36428 18284 36484 18286
rect 36204 18060 36260 18116
rect 35868 17666 35924 17668
rect 35868 17614 35870 17666
rect 35870 17614 35922 17666
rect 35922 17614 35924 17666
rect 35868 17612 35924 17614
rect 35644 17388 35700 17444
rect 34860 14754 34916 14756
rect 34860 14702 34862 14754
rect 34862 14702 34914 14754
rect 34914 14702 34916 14754
rect 34860 14700 34916 14702
rect 33852 11506 33908 11508
rect 33852 11454 33854 11506
rect 33854 11454 33906 11506
rect 33906 11454 33908 11506
rect 33852 11452 33908 11454
rect 34076 11340 34132 11396
rect 33964 9266 34020 9268
rect 33964 9214 33966 9266
rect 33966 9214 34018 9266
rect 34018 9214 34020 9266
rect 33964 9212 34020 9214
rect 33180 7980 33236 8036
rect 33628 6636 33684 6692
rect 33068 5964 33124 6020
rect 30380 5122 30436 5124
rect 30380 5070 30382 5122
rect 30382 5070 30434 5122
rect 30434 5070 30436 5122
rect 30380 5068 30436 5070
rect 33068 5068 33124 5124
rect 32508 4732 32564 4788
rect 33516 4956 33572 5012
rect 33852 4956 33908 5012
rect 35308 11340 35364 11396
rect 35868 17164 35924 17220
rect 35756 16882 35812 16884
rect 35756 16830 35758 16882
rect 35758 16830 35810 16882
rect 35810 16830 35812 16882
rect 35756 16828 35812 16830
rect 35644 15260 35700 15316
rect 35532 15036 35588 15092
rect 35756 15036 35812 15092
rect 37436 20188 37492 20244
rect 37324 18956 37380 19012
rect 37100 18508 37156 18564
rect 37212 18620 37268 18676
rect 36428 17612 36484 17668
rect 36316 16994 36372 16996
rect 36316 16942 36318 16994
rect 36318 16942 36370 16994
rect 36370 16942 36372 16994
rect 36316 16940 36372 16942
rect 36428 16828 36484 16884
rect 36204 14924 36260 14980
rect 36092 14700 36148 14756
rect 35532 13580 35588 13636
rect 35420 11004 35476 11060
rect 34636 10722 34692 10724
rect 34636 10670 34638 10722
rect 34638 10670 34690 10722
rect 34690 10670 34692 10722
rect 34636 10668 34692 10670
rect 35196 9266 35252 9268
rect 35196 9214 35198 9266
rect 35198 9214 35250 9266
rect 35250 9214 35252 9266
rect 35196 9212 35252 9214
rect 35756 9212 35812 9268
rect 35980 14252 36036 14308
rect 36204 13468 36260 13524
rect 36092 12684 36148 12740
rect 36428 15090 36484 15092
rect 36428 15038 36430 15090
rect 36430 15038 36482 15090
rect 36482 15038 36484 15090
rect 36428 15036 36484 15038
rect 36428 13468 36484 13524
rect 37660 20578 37716 20580
rect 37660 20526 37662 20578
rect 37662 20526 37714 20578
rect 37714 20526 37716 20578
rect 37660 20524 37716 20526
rect 37660 19122 37716 19124
rect 37660 19070 37662 19122
rect 37662 19070 37714 19122
rect 37714 19070 37716 19122
rect 37660 19068 37716 19070
rect 37324 18562 37380 18564
rect 37324 18510 37326 18562
rect 37326 18510 37378 18562
rect 37378 18510 37380 18562
rect 37324 18508 37380 18510
rect 37660 18508 37716 18564
rect 37548 18450 37604 18452
rect 37548 18398 37550 18450
rect 37550 18398 37602 18450
rect 37602 18398 37604 18450
rect 37548 18396 37604 18398
rect 37436 17724 37492 17780
rect 37436 17164 37492 17220
rect 37436 15596 37492 15652
rect 36876 15314 36932 15316
rect 36876 15262 36878 15314
rect 36878 15262 36930 15314
rect 36930 15262 36932 15314
rect 36876 15260 36932 15262
rect 36764 14700 36820 14756
rect 36652 12738 36708 12740
rect 36652 12686 36654 12738
rect 36654 12686 36706 12738
rect 36706 12686 36708 12738
rect 36652 12684 36708 12686
rect 36540 11506 36596 11508
rect 36540 11454 36542 11506
rect 36542 11454 36594 11506
rect 36594 11454 36596 11506
rect 36540 11452 36596 11454
rect 36540 11228 36596 11284
rect 34636 4844 34692 4900
rect 34860 4956 34916 5012
rect 34412 4620 34468 4676
rect 34188 4508 34244 4564
rect 34076 4284 34132 4340
rect 36428 7644 36484 7700
rect 36204 6524 36260 6580
rect 36204 6076 36260 6132
rect 36988 14924 37044 14980
rect 36988 14588 37044 14644
rect 37324 14700 37380 14756
rect 39004 23436 39060 23492
rect 39004 23266 39060 23268
rect 39004 23214 39006 23266
rect 39006 23214 39058 23266
rect 39058 23214 39060 23266
rect 39004 23212 39060 23214
rect 41776 37658 41832 37660
rect 41776 37606 41778 37658
rect 41778 37606 41830 37658
rect 41830 37606 41832 37658
rect 41776 37604 41832 37606
rect 41880 37658 41936 37660
rect 41880 37606 41882 37658
rect 41882 37606 41934 37658
rect 41934 37606 41936 37658
rect 41880 37604 41936 37606
rect 41984 37658 42040 37660
rect 41984 37606 41986 37658
rect 41986 37606 42038 37658
rect 42038 37606 42040 37658
rect 41984 37604 42040 37606
rect 42088 37658 42144 37660
rect 42088 37606 42090 37658
rect 42090 37606 42142 37658
rect 42142 37606 42144 37658
rect 42088 37604 42144 37606
rect 42192 37658 42248 37660
rect 42192 37606 42194 37658
rect 42194 37606 42246 37658
rect 42246 37606 42248 37658
rect 42192 37604 42248 37606
rect 42296 37658 42352 37660
rect 42296 37606 42298 37658
rect 42298 37606 42350 37658
rect 42350 37606 42352 37658
rect 42296 37604 42352 37606
rect 44156 36204 44212 36260
rect 45612 37100 45668 37156
rect 41776 36090 41832 36092
rect 41776 36038 41778 36090
rect 41778 36038 41830 36090
rect 41830 36038 41832 36090
rect 41776 36036 41832 36038
rect 41880 36090 41936 36092
rect 41880 36038 41882 36090
rect 41882 36038 41934 36090
rect 41934 36038 41936 36090
rect 41880 36036 41936 36038
rect 41984 36090 42040 36092
rect 41984 36038 41986 36090
rect 41986 36038 42038 36090
rect 42038 36038 42040 36090
rect 41984 36036 42040 36038
rect 42088 36090 42144 36092
rect 42088 36038 42090 36090
rect 42090 36038 42142 36090
rect 42142 36038 42144 36090
rect 42088 36036 42144 36038
rect 42192 36090 42248 36092
rect 42192 36038 42194 36090
rect 42194 36038 42246 36090
rect 42246 36038 42248 36090
rect 42192 36036 42248 36038
rect 42296 36090 42352 36092
rect 42296 36038 42298 36090
rect 42298 36038 42350 36090
rect 42350 36038 42352 36090
rect 42296 36036 42352 36038
rect 41776 34522 41832 34524
rect 41776 34470 41778 34522
rect 41778 34470 41830 34522
rect 41830 34470 41832 34522
rect 41776 34468 41832 34470
rect 41880 34522 41936 34524
rect 41880 34470 41882 34522
rect 41882 34470 41934 34522
rect 41934 34470 41936 34522
rect 41880 34468 41936 34470
rect 41984 34522 42040 34524
rect 41984 34470 41986 34522
rect 41986 34470 42038 34522
rect 42038 34470 42040 34522
rect 41984 34468 42040 34470
rect 42088 34522 42144 34524
rect 42088 34470 42090 34522
rect 42090 34470 42142 34522
rect 42142 34470 42144 34522
rect 42088 34468 42144 34470
rect 42192 34522 42248 34524
rect 42192 34470 42194 34522
rect 42194 34470 42246 34522
rect 42246 34470 42248 34522
rect 42192 34468 42248 34470
rect 42296 34522 42352 34524
rect 42296 34470 42298 34522
rect 42298 34470 42350 34522
rect 42350 34470 42352 34522
rect 42296 34468 42352 34470
rect 41776 32954 41832 32956
rect 41776 32902 41778 32954
rect 41778 32902 41830 32954
rect 41830 32902 41832 32954
rect 41776 32900 41832 32902
rect 41880 32954 41936 32956
rect 41880 32902 41882 32954
rect 41882 32902 41934 32954
rect 41934 32902 41936 32954
rect 41880 32900 41936 32902
rect 41984 32954 42040 32956
rect 41984 32902 41986 32954
rect 41986 32902 42038 32954
rect 42038 32902 42040 32954
rect 41984 32900 42040 32902
rect 42088 32954 42144 32956
rect 42088 32902 42090 32954
rect 42090 32902 42142 32954
rect 42142 32902 42144 32954
rect 42088 32900 42144 32902
rect 42192 32954 42248 32956
rect 42192 32902 42194 32954
rect 42194 32902 42246 32954
rect 42246 32902 42248 32954
rect 42192 32900 42248 32902
rect 42296 32954 42352 32956
rect 42296 32902 42298 32954
rect 42298 32902 42350 32954
rect 42350 32902 42352 32954
rect 42296 32900 42352 32902
rect 44492 32396 44548 32452
rect 41776 31386 41832 31388
rect 41776 31334 41778 31386
rect 41778 31334 41830 31386
rect 41830 31334 41832 31386
rect 41776 31332 41832 31334
rect 41880 31386 41936 31388
rect 41880 31334 41882 31386
rect 41882 31334 41934 31386
rect 41934 31334 41936 31386
rect 41880 31332 41936 31334
rect 41984 31386 42040 31388
rect 41984 31334 41986 31386
rect 41986 31334 42038 31386
rect 42038 31334 42040 31386
rect 41984 31332 42040 31334
rect 42088 31386 42144 31388
rect 42088 31334 42090 31386
rect 42090 31334 42142 31386
rect 42142 31334 42144 31386
rect 42088 31332 42144 31334
rect 42192 31386 42248 31388
rect 42192 31334 42194 31386
rect 42194 31334 42246 31386
rect 42246 31334 42248 31386
rect 42192 31332 42248 31334
rect 42296 31386 42352 31388
rect 42296 31334 42298 31386
rect 42298 31334 42350 31386
rect 42350 31334 42352 31386
rect 42296 31332 42352 31334
rect 41776 29818 41832 29820
rect 41776 29766 41778 29818
rect 41778 29766 41830 29818
rect 41830 29766 41832 29818
rect 41776 29764 41832 29766
rect 41880 29818 41936 29820
rect 41880 29766 41882 29818
rect 41882 29766 41934 29818
rect 41934 29766 41936 29818
rect 41880 29764 41936 29766
rect 41984 29818 42040 29820
rect 41984 29766 41986 29818
rect 41986 29766 42038 29818
rect 42038 29766 42040 29818
rect 41984 29764 42040 29766
rect 42088 29818 42144 29820
rect 42088 29766 42090 29818
rect 42090 29766 42142 29818
rect 42142 29766 42144 29818
rect 42088 29764 42144 29766
rect 42192 29818 42248 29820
rect 42192 29766 42194 29818
rect 42194 29766 42246 29818
rect 42246 29766 42248 29818
rect 42192 29764 42248 29766
rect 42296 29818 42352 29820
rect 42296 29766 42298 29818
rect 42298 29766 42350 29818
rect 42350 29766 42352 29818
rect 42296 29764 42352 29766
rect 41132 25228 41188 25284
rect 41244 29260 41300 29316
rect 39676 23436 39732 23492
rect 38332 22930 38388 22932
rect 38332 22878 38334 22930
rect 38334 22878 38386 22930
rect 38386 22878 38388 22930
rect 38332 22876 38388 22878
rect 38056 22762 38112 22764
rect 38056 22710 38058 22762
rect 38058 22710 38110 22762
rect 38110 22710 38112 22762
rect 38056 22708 38112 22710
rect 38160 22762 38216 22764
rect 38160 22710 38162 22762
rect 38162 22710 38214 22762
rect 38214 22710 38216 22762
rect 38160 22708 38216 22710
rect 38264 22762 38320 22764
rect 38264 22710 38266 22762
rect 38266 22710 38318 22762
rect 38318 22710 38320 22762
rect 38264 22708 38320 22710
rect 38368 22762 38424 22764
rect 38368 22710 38370 22762
rect 38370 22710 38422 22762
rect 38422 22710 38424 22762
rect 38368 22708 38424 22710
rect 38472 22762 38528 22764
rect 38472 22710 38474 22762
rect 38474 22710 38526 22762
rect 38526 22710 38528 22762
rect 38472 22708 38528 22710
rect 38576 22762 38632 22764
rect 38576 22710 38578 22762
rect 38578 22710 38630 22762
rect 38630 22710 38632 22762
rect 38576 22708 38632 22710
rect 38108 22258 38164 22260
rect 38108 22206 38110 22258
rect 38110 22206 38162 22258
rect 38162 22206 38164 22258
rect 38108 22204 38164 22206
rect 38668 22258 38724 22260
rect 38668 22206 38670 22258
rect 38670 22206 38722 22258
rect 38722 22206 38724 22258
rect 38668 22204 38724 22206
rect 37884 21362 37940 21364
rect 37884 21310 37886 21362
rect 37886 21310 37938 21362
rect 37938 21310 37940 21362
rect 37884 21308 37940 21310
rect 38668 21586 38724 21588
rect 38668 21534 38670 21586
rect 38670 21534 38722 21586
rect 38722 21534 38724 21586
rect 38668 21532 38724 21534
rect 38444 21420 38500 21476
rect 38220 21308 38276 21364
rect 38056 21194 38112 21196
rect 38056 21142 38058 21194
rect 38058 21142 38110 21194
rect 38110 21142 38112 21194
rect 38056 21140 38112 21142
rect 38160 21194 38216 21196
rect 38160 21142 38162 21194
rect 38162 21142 38214 21194
rect 38214 21142 38216 21194
rect 38160 21140 38216 21142
rect 38264 21194 38320 21196
rect 38264 21142 38266 21194
rect 38266 21142 38318 21194
rect 38318 21142 38320 21194
rect 38264 21140 38320 21142
rect 38368 21194 38424 21196
rect 38368 21142 38370 21194
rect 38370 21142 38422 21194
rect 38422 21142 38424 21194
rect 38368 21140 38424 21142
rect 38472 21194 38528 21196
rect 38472 21142 38474 21194
rect 38474 21142 38526 21194
rect 38526 21142 38528 21194
rect 38472 21140 38528 21142
rect 38576 21194 38632 21196
rect 38576 21142 38578 21194
rect 38578 21142 38630 21194
rect 38630 21142 38632 21194
rect 38576 21140 38632 21142
rect 37996 21026 38052 21028
rect 37996 20974 37998 21026
rect 37998 20974 38050 21026
rect 38050 20974 38052 21026
rect 37996 20972 38052 20974
rect 38332 20972 38388 21028
rect 38668 20972 38724 21028
rect 40348 21532 40404 21588
rect 38332 20188 38388 20244
rect 37996 20130 38052 20132
rect 37996 20078 37998 20130
rect 37998 20078 38050 20130
rect 38050 20078 38052 20130
rect 37996 20076 38052 20078
rect 38220 20018 38276 20020
rect 38220 19966 38222 20018
rect 38222 19966 38274 20018
rect 38274 19966 38276 20018
rect 38220 19964 38276 19966
rect 39900 21308 39956 21364
rect 39452 20690 39508 20692
rect 39452 20638 39454 20690
rect 39454 20638 39506 20690
rect 39506 20638 39508 20690
rect 39452 20636 39508 20638
rect 40012 20690 40068 20692
rect 40012 20638 40014 20690
rect 40014 20638 40066 20690
rect 40066 20638 40068 20690
rect 40012 20636 40068 20638
rect 38780 19964 38836 20020
rect 38056 19626 38112 19628
rect 38056 19574 38058 19626
rect 38058 19574 38110 19626
rect 38110 19574 38112 19626
rect 38056 19572 38112 19574
rect 38160 19626 38216 19628
rect 38160 19574 38162 19626
rect 38162 19574 38214 19626
rect 38214 19574 38216 19626
rect 38160 19572 38216 19574
rect 38264 19626 38320 19628
rect 38264 19574 38266 19626
rect 38266 19574 38318 19626
rect 38318 19574 38320 19626
rect 38264 19572 38320 19574
rect 38368 19626 38424 19628
rect 38368 19574 38370 19626
rect 38370 19574 38422 19626
rect 38422 19574 38424 19626
rect 38368 19572 38424 19574
rect 38472 19626 38528 19628
rect 38472 19574 38474 19626
rect 38474 19574 38526 19626
rect 38526 19574 38528 19626
rect 38472 19572 38528 19574
rect 38576 19626 38632 19628
rect 38576 19574 38578 19626
rect 38578 19574 38630 19626
rect 38630 19574 38632 19626
rect 38576 19572 38632 19574
rect 39116 20524 39172 20580
rect 39676 20578 39732 20580
rect 39676 20526 39678 20578
rect 39678 20526 39730 20578
rect 39730 20526 39732 20578
rect 39676 20524 39732 20526
rect 37996 19458 38052 19460
rect 37996 19406 37998 19458
rect 37998 19406 38050 19458
rect 38050 19406 38052 19458
rect 37996 19404 38052 19406
rect 38780 19122 38836 19124
rect 38780 19070 38782 19122
rect 38782 19070 38834 19122
rect 38834 19070 38836 19122
rect 38780 19068 38836 19070
rect 38108 18732 38164 18788
rect 38780 18732 38836 18788
rect 38556 18450 38612 18452
rect 38556 18398 38558 18450
rect 38558 18398 38610 18450
rect 38610 18398 38612 18450
rect 38556 18396 38612 18398
rect 38780 18396 38836 18452
rect 38056 18058 38112 18060
rect 38056 18006 38058 18058
rect 38058 18006 38110 18058
rect 38110 18006 38112 18058
rect 38056 18004 38112 18006
rect 38160 18058 38216 18060
rect 38160 18006 38162 18058
rect 38162 18006 38214 18058
rect 38214 18006 38216 18058
rect 38160 18004 38216 18006
rect 38264 18058 38320 18060
rect 38264 18006 38266 18058
rect 38266 18006 38318 18058
rect 38318 18006 38320 18058
rect 38264 18004 38320 18006
rect 38368 18058 38424 18060
rect 38368 18006 38370 18058
rect 38370 18006 38422 18058
rect 38422 18006 38424 18058
rect 38368 18004 38424 18006
rect 38472 18058 38528 18060
rect 38472 18006 38474 18058
rect 38474 18006 38526 18058
rect 38526 18006 38528 18058
rect 38472 18004 38528 18006
rect 38576 18058 38632 18060
rect 38576 18006 38578 18058
rect 38578 18006 38630 18058
rect 38630 18006 38632 18058
rect 38576 18004 38632 18006
rect 37884 17554 37940 17556
rect 37884 17502 37886 17554
rect 37886 17502 37938 17554
rect 37938 17502 37940 17554
rect 37884 17500 37940 17502
rect 37772 17052 37828 17108
rect 38220 17164 38276 17220
rect 38056 16490 38112 16492
rect 38056 16438 38058 16490
rect 38058 16438 38110 16490
rect 38110 16438 38112 16490
rect 38056 16436 38112 16438
rect 38160 16490 38216 16492
rect 38160 16438 38162 16490
rect 38162 16438 38214 16490
rect 38214 16438 38216 16490
rect 38160 16436 38216 16438
rect 38264 16490 38320 16492
rect 38264 16438 38266 16490
rect 38266 16438 38318 16490
rect 38318 16438 38320 16490
rect 38264 16436 38320 16438
rect 38368 16490 38424 16492
rect 38368 16438 38370 16490
rect 38370 16438 38422 16490
rect 38422 16438 38424 16490
rect 38368 16436 38424 16438
rect 38472 16490 38528 16492
rect 38472 16438 38474 16490
rect 38474 16438 38526 16490
rect 38526 16438 38528 16490
rect 38472 16436 38528 16438
rect 38576 16490 38632 16492
rect 38576 16438 38578 16490
rect 38578 16438 38630 16490
rect 38630 16438 38632 16490
rect 38576 16436 38632 16438
rect 40796 20690 40852 20692
rect 40796 20638 40798 20690
rect 40798 20638 40850 20690
rect 40850 20638 40852 20690
rect 40796 20636 40852 20638
rect 41776 28250 41832 28252
rect 41776 28198 41778 28250
rect 41778 28198 41830 28250
rect 41830 28198 41832 28250
rect 41776 28196 41832 28198
rect 41880 28250 41936 28252
rect 41880 28198 41882 28250
rect 41882 28198 41934 28250
rect 41934 28198 41936 28250
rect 41880 28196 41936 28198
rect 41984 28250 42040 28252
rect 41984 28198 41986 28250
rect 41986 28198 42038 28250
rect 42038 28198 42040 28250
rect 41984 28196 42040 28198
rect 42088 28250 42144 28252
rect 42088 28198 42090 28250
rect 42090 28198 42142 28250
rect 42142 28198 42144 28250
rect 42088 28196 42144 28198
rect 42192 28250 42248 28252
rect 42192 28198 42194 28250
rect 42194 28198 42246 28250
rect 42246 28198 42248 28250
rect 42192 28196 42248 28198
rect 42296 28250 42352 28252
rect 42296 28198 42298 28250
rect 42298 28198 42350 28250
rect 42350 28198 42352 28250
rect 42296 28196 42352 28198
rect 42812 26908 42868 26964
rect 41776 26682 41832 26684
rect 41776 26630 41778 26682
rect 41778 26630 41830 26682
rect 41830 26630 41832 26682
rect 41776 26628 41832 26630
rect 41880 26682 41936 26684
rect 41880 26630 41882 26682
rect 41882 26630 41934 26682
rect 41934 26630 41936 26682
rect 41880 26628 41936 26630
rect 41984 26682 42040 26684
rect 41984 26630 41986 26682
rect 41986 26630 42038 26682
rect 42038 26630 42040 26682
rect 41984 26628 42040 26630
rect 42088 26682 42144 26684
rect 42088 26630 42090 26682
rect 42090 26630 42142 26682
rect 42142 26630 42144 26682
rect 42088 26628 42144 26630
rect 42192 26682 42248 26684
rect 42192 26630 42194 26682
rect 42194 26630 42246 26682
rect 42246 26630 42248 26682
rect 42192 26628 42248 26630
rect 42296 26682 42352 26684
rect 42296 26630 42298 26682
rect 42298 26630 42350 26682
rect 42350 26630 42352 26682
rect 42296 26628 42352 26630
rect 41776 25114 41832 25116
rect 41776 25062 41778 25114
rect 41778 25062 41830 25114
rect 41830 25062 41832 25114
rect 41776 25060 41832 25062
rect 41880 25114 41936 25116
rect 41880 25062 41882 25114
rect 41882 25062 41934 25114
rect 41934 25062 41936 25114
rect 41880 25060 41936 25062
rect 41984 25114 42040 25116
rect 41984 25062 41986 25114
rect 41986 25062 42038 25114
rect 42038 25062 42040 25114
rect 41984 25060 42040 25062
rect 42088 25114 42144 25116
rect 42088 25062 42090 25114
rect 42090 25062 42142 25114
rect 42142 25062 42144 25114
rect 42088 25060 42144 25062
rect 42192 25114 42248 25116
rect 42192 25062 42194 25114
rect 42194 25062 42246 25114
rect 42246 25062 42248 25114
rect 42192 25060 42248 25062
rect 42296 25114 42352 25116
rect 42296 25062 42298 25114
rect 42298 25062 42350 25114
rect 42350 25062 42352 25114
rect 42296 25060 42352 25062
rect 41776 23546 41832 23548
rect 41776 23494 41778 23546
rect 41778 23494 41830 23546
rect 41830 23494 41832 23546
rect 41776 23492 41832 23494
rect 41880 23546 41936 23548
rect 41880 23494 41882 23546
rect 41882 23494 41934 23546
rect 41934 23494 41936 23546
rect 41880 23492 41936 23494
rect 41984 23546 42040 23548
rect 41984 23494 41986 23546
rect 41986 23494 42038 23546
rect 42038 23494 42040 23546
rect 41984 23492 42040 23494
rect 42088 23546 42144 23548
rect 42088 23494 42090 23546
rect 42090 23494 42142 23546
rect 42142 23494 42144 23546
rect 42088 23492 42144 23494
rect 42192 23546 42248 23548
rect 42192 23494 42194 23546
rect 42194 23494 42246 23546
rect 42246 23494 42248 23546
rect 42192 23492 42248 23494
rect 42296 23546 42352 23548
rect 42296 23494 42298 23546
rect 42298 23494 42350 23546
rect 42350 23494 42352 23546
rect 42296 23492 42352 23494
rect 41776 21978 41832 21980
rect 41776 21926 41778 21978
rect 41778 21926 41830 21978
rect 41830 21926 41832 21978
rect 41776 21924 41832 21926
rect 41880 21978 41936 21980
rect 41880 21926 41882 21978
rect 41882 21926 41934 21978
rect 41934 21926 41936 21978
rect 41880 21924 41936 21926
rect 41984 21978 42040 21980
rect 41984 21926 41986 21978
rect 41986 21926 42038 21978
rect 42038 21926 42040 21978
rect 41984 21924 42040 21926
rect 42088 21978 42144 21980
rect 42088 21926 42090 21978
rect 42090 21926 42142 21978
rect 42142 21926 42144 21978
rect 42088 21924 42144 21926
rect 42192 21978 42248 21980
rect 42192 21926 42194 21978
rect 42194 21926 42246 21978
rect 42246 21926 42248 21978
rect 42192 21924 42248 21926
rect 42296 21978 42352 21980
rect 42296 21926 42298 21978
rect 42298 21926 42350 21978
rect 42350 21926 42352 21978
rect 42296 21924 42352 21926
rect 41244 18956 41300 19012
rect 41580 20636 41636 20692
rect 40348 18396 40404 18452
rect 37660 15596 37716 15652
rect 37884 15932 37940 15988
rect 37660 15036 37716 15092
rect 39116 15538 39172 15540
rect 39116 15486 39118 15538
rect 39118 15486 39170 15538
rect 39170 15486 39172 15538
rect 39116 15484 39172 15486
rect 38892 15372 38948 15428
rect 38220 15148 38276 15204
rect 37996 15036 38052 15092
rect 38780 15036 38836 15092
rect 38056 14922 38112 14924
rect 38056 14870 38058 14922
rect 38058 14870 38110 14922
rect 38110 14870 38112 14922
rect 38056 14868 38112 14870
rect 38160 14922 38216 14924
rect 38160 14870 38162 14922
rect 38162 14870 38214 14922
rect 38214 14870 38216 14922
rect 38160 14868 38216 14870
rect 38264 14922 38320 14924
rect 38264 14870 38266 14922
rect 38266 14870 38318 14922
rect 38318 14870 38320 14922
rect 38264 14868 38320 14870
rect 38368 14922 38424 14924
rect 38368 14870 38370 14922
rect 38370 14870 38422 14922
rect 38422 14870 38424 14922
rect 38368 14868 38424 14870
rect 38472 14922 38528 14924
rect 38472 14870 38474 14922
rect 38474 14870 38526 14922
rect 38526 14870 38528 14922
rect 38472 14868 38528 14870
rect 38576 14922 38632 14924
rect 38576 14870 38578 14922
rect 38578 14870 38630 14922
rect 38630 14870 38632 14922
rect 38576 14868 38632 14870
rect 37660 14364 37716 14420
rect 38108 14418 38164 14420
rect 38108 14366 38110 14418
rect 38110 14366 38162 14418
rect 38162 14366 38164 14418
rect 38108 14364 38164 14366
rect 37884 14140 37940 14196
rect 36876 10556 36932 10612
rect 38444 14642 38500 14644
rect 38444 14590 38446 14642
rect 38446 14590 38498 14642
rect 38498 14590 38500 14642
rect 38444 14588 38500 14590
rect 39004 13970 39060 13972
rect 39004 13918 39006 13970
rect 39006 13918 39058 13970
rect 39058 13918 39060 13970
rect 39004 13916 39060 13918
rect 36652 5852 36708 5908
rect 36764 6524 36820 6580
rect 35756 4396 35812 4452
rect 34636 4338 34692 4340
rect 34636 4286 34638 4338
rect 34638 4286 34690 4338
rect 34690 4286 34692 4338
rect 34636 4284 34692 4286
rect 29260 3666 29316 3668
rect 29260 3614 29262 3666
rect 29262 3614 29314 3666
rect 29314 3614 29316 3666
rect 29260 3612 29316 3614
rect 30156 3666 30212 3668
rect 30156 3614 30158 3666
rect 30158 3614 30210 3666
rect 30210 3614 30212 3666
rect 30156 3612 30212 3614
rect 35420 3612 35476 3668
rect 26348 3442 26404 3444
rect 26348 3390 26350 3442
rect 26350 3390 26402 3442
rect 26402 3390 26404 3442
rect 26348 3388 26404 3390
rect 29708 3442 29764 3444
rect 29708 3390 29710 3442
rect 29710 3390 29762 3442
rect 29762 3390 29764 3442
rect 29708 3388 29764 3390
rect 38056 13354 38112 13356
rect 38056 13302 38058 13354
rect 38058 13302 38110 13354
rect 38110 13302 38112 13354
rect 38056 13300 38112 13302
rect 38160 13354 38216 13356
rect 38160 13302 38162 13354
rect 38162 13302 38214 13354
rect 38214 13302 38216 13354
rect 38160 13300 38216 13302
rect 38264 13354 38320 13356
rect 38264 13302 38266 13354
rect 38266 13302 38318 13354
rect 38318 13302 38320 13354
rect 38264 13300 38320 13302
rect 38368 13354 38424 13356
rect 38368 13302 38370 13354
rect 38370 13302 38422 13354
rect 38422 13302 38424 13354
rect 38368 13300 38424 13302
rect 38472 13354 38528 13356
rect 38472 13302 38474 13354
rect 38474 13302 38526 13354
rect 38526 13302 38528 13354
rect 38472 13300 38528 13302
rect 38576 13354 38632 13356
rect 38576 13302 38578 13354
rect 38578 13302 38630 13354
rect 38630 13302 38632 13354
rect 38576 13300 38632 13302
rect 38556 13132 38612 13188
rect 37436 12738 37492 12740
rect 37436 12686 37438 12738
rect 37438 12686 37490 12738
rect 37490 12686 37492 12738
rect 37436 12684 37492 12686
rect 39340 15372 39396 15428
rect 39452 16828 39508 16884
rect 39340 15148 39396 15204
rect 39452 15036 39508 15092
rect 39340 13132 39396 13188
rect 38056 11786 38112 11788
rect 38056 11734 38058 11786
rect 38058 11734 38110 11786
rect 38110 11734 38112 11786
rect 38056 11732 38112 11734
rect 38160 11786 38216 11788
rect 38160 11734 38162 11786
rect 38162 11734 38214 11786
rect 38214 11734 38216 11786
rect 38160 11732 38216 11734
rect 38264 11786 38320 11788
rect 38264 11734 38266 11786
rect 38266 11734 38318 11786
rect 38318 11734 38320 11786
rect 38264 11732 38320 11734
rect 38368 11786 38424 11788
rect 38368 11734 38370 11786
rect 38370 11734 38422 11786
rect 38422 11734 38424 11786
rect 38368 11732 38424 11734
rect 38472 11786 38528 11788
rect 38472 11734 38474 11786
rect 38474 11734 38526 11786
rect 38526 11734 38528 11786
rect 38472 11732 38528 11734
rect 38576 11786 38632 11788
rect 38576 11734 38578 11786
rect 38578 11734 38630 11786
rect 38630 11734 38632 11786
rect 38576 11732 38632 11734
rect 38332 11564 38388 11620
rect 37212 11340 37268 11396
rect 37660 11340 37716 11396
rect 37660 10668 37716 10724
rect 38780 10444 38836 10500
rect 38056 10218 38112 10220
rect 38056 10166 38058 10218
rect 38058 10166 38110 10218
rect 38110 10166 38112 10218
rect 38056 10164 38112 10166
rect 38160 10218 38216 10220
rect 38160 10166 38162 10218
rect 38162 10166 38214 10218
rect 38214 10166 38216 10218
rect 38160 10164 38216 10166
rect 38264 10218 38320 10220
rect 38264 10166 38266 10218
rect 38266 10166 38318 10218
rect 38318 10166 38320 10218
rect 38264 10164 38320 10166
rect 38368 10218 38424 10220
rect 38368 10166 38370 10218
rect 38370 10166 38422 10218
rect 38422 10166 38424 10218
rect 38368 10164 38424 10166
rect 38472 10218 38528 10220
rect 38472 10166 38474 10218
rect 38474 10166 38526 10218
rect 38526 10166 38528 10218
rect 38472 10164 38528 10166
rect 38576 10218 38632 10220
rect 38576 10166 38578 10218
rect 38578 10166 38630 10218
rect 38630 10166 38632 10218
rect 38576 10164 38632 10166
rect 37548 9548 37604 9604
rect 38056 8650 38112 8652
rect 38056 8598 38058 8650
rect 38058 8598 38110 8650
rect 38110 8598 38112 8650
rect 38056 8596 38112 8598
rect 38160 8650 38216 8652
rect 38160 8598 38162 8650
rect 38162 8598 38214 8650
rect 38214 8598 38216 8650
rect 38160 8596 38216 8598
rect 38264 8650 38320 8652
rect 38264 8598 38266 8650
rect 38266 8598 38318 8650
rect 38318 8598 38320 8650
rect 38264 8596 38320 8598
rect 38368 8650 38424 8652
rect 38368 8598 38370 8650
rect 38370 8598 38422 8650
rect 38422 8598 38424 8650
rect 38368 8596 38424 8598
rect 38472 8650 38528 8652
rect 38472 8598 38474 8650
rect 38474 8598 38526 8650
rect 38526 8598 38528 8650
rect 38472 8596 38528 8598
rect 38576 8650 38632 8652
rect 38576 8598 38578 8650
rect 38578 8598 38630 8650
rect 38630 8598 38632 8650
rect 38576 8596 38632 8598
rect 38556 8428 38612 8484
rect 39676 14306 39732 14308
rect 39676 14254 39678 14306
rect 39678 14254 39730 14306
rect 39730 14254 39732 14306
rect 39676 14252 39732 14254
rect 39564 11452 39620 11508
rect 41776 20410 41832 20412
rect 41776 20358 41778 20410
rect 41778 20358 41830 20410
rect 41830 20358 41832 20410
rect 41776 20356 41832 20358
rect 41880 20410 41936 20412
rect 41880 20358 41882 20410
rect 41882 20358 41934 20410
rect 41934 20358 41936 20410
rect 41880 20356 41936 20358
rect 41984 20410 42040 20412
rect 41984 20358 41986 20410
rect 41986 20358 42038 20410
rect 42038 20358 42040 20410
rect 41984 20356 42040 20358
rect 42088 20410 42144 20412
rect 42088 20358 42090 20410
rect 42090 20358 42142 20410
rect 42142 20358 42144 20410
rect 42088 20356 42144 20358
rect 42192 20410 42248 20412
rect 42192 20358 42194 20410
rect 42194 20358 42246 20410
rect 42246 20358 42248 20410
rect 42192 20356 42248 20358
rect 42296 20410 42352 20412
rect 42296 20358 42298 20410
rect 42298 20358 42350 20410
rect 42350 20358 42352 20410
rect 42296 20356 42352 20358
rect 41776 18842 41832 18844
rect 41776 18790 41778 18842
rect 41778 18790 41830 18842
rect 41830 18790 41832 18842
rect 41776 18788 41832 18790
rect 41880 18842 41936 18844
rect 41880 18790 41882 18842
rect 41882 18790 41934 18842
rect 41934 18790 41936 18842
rect 41880 18788 41936 18790
rect 41984 18842 42040 18844
rect 41984 18790 41986 18842
rect 41986 18790 42038 18842
rect 42038 18790 42040 18842
rect 41984 18788 42040 18790
rect 42088 18842 42144 18844
rect 42088 18790 42090 18842
rect 42090 18790 42142 18842
rect 42142 18790 42144 18842
rect 42088 18788 42144 18790
rect 42192 18842 42248 18844
rect 42192 18790 42194 18842
rect 42194 18790 42246 18842
rect 42246 18790 42248 18842
rect 42192 18788 42248 18790
rect 42296 18842 42352 18844
rect 42296 18790 42298 18842
rect 42298 18790 42350 18842
rect 42350 18790 42352 18842
rect 42296 18788 42352 18790
rect 45500 31052 45556 31108
rect 45500 24780 45556 24836
rect 45612 23212 45668 23268
rect 45724 28588 45780 28644
rect 44492 20076 44548 20132
rect 42812 17612 42868 17668
rect 41776 17274 41832 17276
rect 41776 17222 41778 17274
rect 41778 17222 41830 17274
rect 41830 17222 41832 17274
rect 41776 17220 41832 17222
rect 41880 17274 41936 17276
rect 41880 17222 41882 17274
rect 41882 17222 41934 17274
rect 41934 17222 41936 17274
rect 41880 17220 41936 17222
rect 41984 17274 42040 17276
rect 41984 17222 41986 17274
rect 41986 17222 42038 17274
rect 42038 17222 42040 17274
rect 41984 17220 42040 17222
rect 42088 17274 42144 17276
rect 42088 17222 42090 17274
rect 42090 17222 42142 17274
rect 42142 17222 42144 17274
rect 42088 17220 42144 17222
rect 42192 17274 42248 17276
rect 42192 17222 42194 17274
rect 42194 17222 42246 17274
rect 42246 17222 42248 17274
rect 42192 17220 42248 17222
rect 42296 17274 42352 17276
rect 42296 17222 42298 17274
rect 42298 17222 42350 17274
rect 42350 17222 42352 17274
rect 42296 17220 42352 17222
rect 47740 45276 47796 45332
rect 47740 43820 47796 43876
rect 46284 41916 46340 41972
rect 47740 42364 47796 42420
rect 46844 41916 46900 41972
rect 47740 40908 47796 40964
rect 47740 39506 47796 39508
rect 47740 39454 47742 39506
rect 47742 39454 47794 39506
rect 47794 39454 47796 39506
rect 47740 39452 47796 39454
rect 46396 38722 46452 38724
rect 46396 38670 46398 38722
rect 46398 38670 46450 38722
rect 46450 38670 46452 38722
rect 46396 38668 46452 38670
rect 46396 37154 46452 37156
rect 46396 37102 46398 37154
rect 46398 37102 46450 37154
rect 46450 37102 46452 37154
rect 46396 37100 46452 37102
rect 46396 35698 46452 35700
rect 46396 35646 46398 35698
rect 46398 35646 46450 35698
rect 46450 35646 46452 35698
rect 46396 35644 46452 35646
rect 46396 32450 46452 32452
rect 46396 32398 46398 32450
rect 46398 32398 46450 32450
rect 46450 32398 46452 32450
rect 46396 32396 46452 32398
rect 46060 29484 46116 29540
rect 45948 28028 46004 28084
rect 45836 27916 45892 27972
rect 46396 29314 46452 29316
rect 46396 29262 46398 29314
rect 46398 29262 46450 29314
rect 46450 29262 46452 29314
rect 46396 29260 46452 29262
rect 46284 28642 46340 28644
rect 46284 28590 46286 28642
rect 46286 28590 46338 28642
rect 46338 28590 46340 28642
rect 46284 28588 46340 28590
rect 46284 26962 46340 26964
rect 46284 26910 46286 26962
rect 46286 26910 46338 26962
rect 46338 26910 46340 26962
rect 46284 26908 46340 26910
rect 45836 25676 45892 25732
rect 46844 38668 46900 38724
rect 47852 38722 47908 38724
rect 47852 38670 47854 38722
rect 47854 38670 47906 38722
rect 47906 38670 47908 38722
rect 47852 38668 47908 38670
rect 46844 37100 46900 37156
rect 47852 36540 47908 36596
rect 46956 35698 47012 35700
rect 46956 35646 46958 35698
rect 46958 35646 47010 35698
rect 47010 35646 47012 35698
rect 46956 35644 47012 35646
rect 46844 32396 46900 32452
rect 46732 31052 46788 31108
rect 46844 29260 46900 29316
rect 46844 28642 46900 28644
rect 46844 28590 46846 28642
rect 46846 28590 46898 28642
rect 46898 28590 46900 28642
rect 46844 28588 46900 28590
rect 46844 26908 46900 26964
rect 46620 26348 46676 26404
rect 46956 25676 47012 25732
rect 46060 20972 46116 21028
rect 46284 22146 46340 22148
rect 46284 22094 46286 22146
rect 46286 22094 46338 22146
rect 46338 22094 46340 22146
rect 46284 22092 46340 22094
rect 46844 22092 46900 22148
rect 45836 19068 45892 19124
rect 45724 17052 45780 17108
rect 40012 15986 40068 15988
rect 40012 15934 40014 15986
rect 40014 15934 40066 15986
rect 40066 15934 40068 15986
rect 40012 15932 40068 15934
rect 40012 15314 40068 15316
rect 40012 15262 40014 15314
rect 40014 15262 40066 15314
rect 40066 15262 40068 15314
rect 40012 15260 40068 15262
rect 39900 13916 39956 13972
rect 40012 14364 40068 14420
rect 40124 13692 40180 13748
rect 46060 17388 46116 17444
rect 45948 16044 46004 16100
rect 40796 15484 40852 15540
rect 41776 15706 41832 15708
rect 41776 15654 41778 15706
rect 41778 15654 41830 15706
rect 41830 15654 41832 15706
rect 41776 15652 41832 15654
rect 41880 15706 41936 15708
rect 41880 15654 41882 15706
rect 41882 15654 41934 15706
rect 41934 15654 41936 15706
rect 41880 15652 41936 15654
rect 41984 15706 42040 15708
rect 41984 15654 41986 15706
rect 41986 15654 42038 15706
rect 42038 15654 42040 15706
rect 41984 15652 42040 15654
rect 42088 15706 42144 15708
rect 42088 15654 42090 15706
rect 42090 15654 42142 15706
rect 42142 15654 42144 15706
rect 42088 15652 42144 15654
rect 42192 15706 42248 15708
rect 42192 15654 42194 15706
rect 42194 15654 42246 15706
rect 42246 15654 42248 15706
rect 42192 15652 42248 15654
rect 42296 15706 42352 15708
rect 42296 15654 42298 15706
rect 42298 15654 42350 15706
rect 42350 15654 42352 15706
rect 42296 15652 42352 15654
rect 41468 15314 41524 15316
rect 41468 15262 41470 15314
rect 41470 15262 41522 15314
rect 41522 15262 41524 15314
rect 41468 15260 41524 15262
rect 40572 14418 40628 14420
rect 40572 14366 40574 14418
rect 40574 14366 40626 14418
rect 40626 14366 40628 14418
rect 40572 14364 40628 14366
rect 46396 16882 46452 16884
rect 46396 16830 46398 16882
rect 46398 16830 46450 16882
rect 46450 16830 46452 16882
rect 46396 16828 46452 16830
rect 46284 15314 46340 15316
rect 46284 15262 46286 15314
rect 46286 15262 46338 15314
rect 46338 15262 46340 15314
rect 46284 15260 46340 15262
rect 46172 14588 46228 14644
rect 40684 13746 40740 13748
rect 40684 13694 40686 13746
rect 40686 13694 40738 13746
rect 40738 13694 40740 13746
rect 40684 13692 40740 13694
rect 47852 35308 47908 35364
rect 47852 33628 47908 33684
rect 47852 32172 47908 32228
rect 47852 30716 47908 30772
rect 47852 29314 47908 29316
rect 47852 29262 47854 29314
rect 47854 29262 47906 29314
rect 47906 29262 47908 29314
rect 47852 29260 47908 29262
rect 47852 27804 47908 27860
rect 47740 26348 47796 26404
rect 47740 24892 47796 24948
rect 47740 23436 47796 23492
rect 47740 21980 47796 22036
rect 47068 20860 47124 20916
rect 47740 20524 47796 20580
rect 47740 19122 47796 19124
rect 47740 19070 47742 19122
rect 47742 19070 47794 19122
rect 47794 19070 47796 19122
rect 47740 19068 47796 19070
rect 47852 17612 47908 17668
rect 46956 16940 47012 16996
rect 46844 16882 46900 16884
rect 46844 16830 46846 16882
rect 46846 16830 46898 16882
rect 46898 16830 46900 16882
rect 46844 16828 46900 16830
rect 47740 16882 47796 16884
rect 47740 16830 47742 16882
rect 47742 16830 47794 16882
rect 47794 16830 47796 16882
rect 47740 16828 47796 16830
rect 46844 15314 46900 15316
rect 46844 15262 46846 15314
rect 46846 15262 46898 15314
rect 46898 15262 46900 15314
rect 46844 15260 46900 15262
rect 47852 14700 47908 14756
rect 46508 14252 46564 14308
rect 41776 14138 41832 14140
rect 41776 14086 41778 14138
rect 41778 14086 41830 14138
rect 41830 14086 41832 14138
rect 41776 14084 41832 14086
rect 41880 14138 41936 14140
rect 41880 14086 41882 14138
rect 41882 14086 41934 14138
rect 41934 14086 41936 14138
rect 41880 14084 41936 14086
rect 41984 14138 42040 14140
rect 41984 14086 41986 14138
rect 41986 14086 42038 14138
rect 42038 14086 42040 14138
rect 41984 14084 42040 14086
rect 42088 14138 42144 14140
rect 42088 14086 42090 14138
rect 42090 14086 42142 14138
rect 42142 14086 42144 14138
rect 42088 14084 42144 14086
rect 42192 14138 42248 14140
rect 42192 14086 42194 14138
rect 42194 14086 42246 14138
rect 42246 14086 42248 14138
rect 42192 14084 42248 14086
rect 42296 14138 42352 14140
rect 42296 14086 42298 14138
rect 42298 14086 42350 14138
rect 42350 14086 42352 14138
rect 42296 14084 42352 14086
rect 42476 13692 42532 13748
rect 40348 11788 40404 11844
rect 40460 11676 40516 11732
rect 40796 12348 40852 12404
rect 41916 12850 41972 12852
rect 41916 12798 41918 12850
rect 41918 12798 41970 12850
rect 41970 12798 41972 12850
rect 41916 12796 41972 12798
rect 41776 12570 41832 12572
rect 41776 12518 41778 12570
rect 41778 12518 41830 12570
rect 41830 12518 41832 12570
rect 41776 12516 41832 12518
rect 41880 12570 41936 12572
rect 41880 12518 41882 12570
rect 41882 12518 41934 12570
rect 41934 12518 41936 12570
rect 41880 12516 41936 12518
rect 41984 12570 42040 12572
rect 41984 12518 41986 12570
rect 41986 12518 42038 12570
rect 42038 12518 42040 12570
rect 41984 12516 42040 12518
rect 42088 12570 42144 12572
rect 42088 12518 42090 12570
rect 42090 12518 42142 12570
rect 42142 12518 42144 12570
rect 42088 12516 42144 12518
rect 42192 12570 42248 12572
rect 42192 12518 42194 12570
rect 42194 12518 42246 12570
rect 42246 12518 42248 12570
rect 42192 12516 42248 12518
rect 42296 12570 42352 12572
rect 42296 12518 42298 12570
rect 42298 12518 42350 12570
rect 42350 12518 42352 12570
rect 42296 12516 42352 12518
rect 46284 13746 46340 13748
rect 46284 13694 46286 13746
rect 46286 13694 46338 13746
rect 46338 13694 46340 13746
rect 46284 13692 46340 13694
rect 46844 13746 46900 13748
rect 46844 13694 46846 13746
rect 46846 13694 46898 13746
rect 46898 13694 46900 13746
rect 46844 13692 46900 13694
rect 47852 13468 47908 13524
rect 42700 12796 42756 12852
rect 41132 11788 41188 11844
rect 40684 11340 40740 11396
rect 40572 11228 40628 11284
rect 41468 11228 41524 11284
rect 40796 10498 40852 10500
rect 40796 10446 40798 10498
rect 40798 10446 40850 10498
rect 40850 10446 40852 10498
rect 40796 10444 40852 10446
rect 39788 9324 39844 9380
rect 41132 8428 41188 8484
rect 38892 8092 38948 8148
rect 40684 8146 40740 8148
rect 40684 8094 40686 8146
rect 40686 8094 40738 8146
rect 40738 8094 40740 8146
rect 40684 8092 40740 8094
rect 39004 7698 39060 7700
rect 39004 7646 39006 7698
rect 39006 7646 39058 7698
rect 39058 7646 39060 7698
rect 39004 7644 39060 7646
rect 41692 12066 41748 12068
rect 41692 12014 41694 12066
rect 41694 12014 41746 12066
rect 41746 12014 41748 12066
rect 41692 12012 41748 12014
rect 42028 11788 42084 11844
rect 42588 12290 42644 12292
rect 42588 12238 42590 12290
rect 42590 12238 42642 12290
rect 42642 12238 42644 12290
rect 42588 12236 42644 12238
rect 42364 11282 42420 11284
rect 42364 11230 42366 11282
rect 42366 11230 42418 11282
rect 42418 11230 42420 11282
rect 42364 11228 42420 11230
rect 41776 11002 41832 11004
rect 41776 10950 41778 11002
rect 41778 10950 41830 11002
rect 41830 10950 41832 11002
rect 41776 10948 41832 10950
rect 41880 11002 41936 11004
rect 41880 10950 41882 11002
rect 41882 10950 41934 11002
rect 41934 10950 41936 11002
rect 41880 10948 41936 10950
rect 41984 11002 42040 11004
rect 41984 10950 41986 11002
rect 41986 10950 42038 11002
rect 42038 10950 42040 11002
rect 41984 10948 42040 10950
rect 42088 11002 42144 11004
rect 42088 10950 42090 11002
rect 42090 10950 42142 11002
rect 42142 10950 42144 11002
rect 42088 10948 42144 10950
rect 42192 11002 42248 11004
rect 42192 10950 42194 11002
rect 42194 10950 42246 11002
rect 42246 10950 42248 11002
rect 42192 10948 42248 10950
rect 42296 11002 42352 11004
rect 42296 10950 42298 11002
rect 42298 10950 42350 11002
rect 42350 10950 42352 11002
rect 42296 10948 42352 10950
rect 42028 10498 42084 10500
rect 42028 10446 42030 10498
rect 42030 10446 42082 10498
rect 42082 10446 42084 10498
rect 42028 10444 42084 10446
rect 43372 12290 43428 12292
rect 43372 12238 43374 12290
rect 43374 12238 43426 12290
rect 43426 12238 43428 12290
rect 43372 12236 43428 12238
rect 46284 12290 46340 12292
rect 46284 12238 46286 12290
rect 46286 12238 46338 12290
rect 46338 12238 46340 12290
rect 46284 12236 46340 12238
rect 46844 12236 46900 12292
rect 42476 10444 42532 10500
rect 42588 9996 42644 10052
rect 42140 9602 42196 9604
rect 42140 9550 42142 9602
rect 42142 9550 42194 9602
rect 42194 9550 42196 9602
rect 42140 9548 42196 9550
rect 41776 9434 41832 9436
rect 41776 9382 41778 9434
rect 41778 9382 41830 9434
rect 41830 9382 41832 9434
rect 41776 9380 41832 9382
rect 41880 9434 41936 9436
rect 41880 9382 41882 9434
rect 41882 9382 41934 9434
rect 41934 9382 41936 9434
rect 41880 9380 41936 9382
rect 41984 9434 42040 9436
rect 41984 9382 41986 9434
rect 41986 9382 42038 9434
rect 42038 9382 42040 9434
rect 41984 9380 42040 9382
rect 42088 9434 42144 9436
rect 42088 9382 42090 9434
rect 42090 9382 42142 9434
rect 42142 9382 42144 9434
rect 42088 9380 42144 9382
rect 42192 9434 42248 9436
rect 42192 9382 42194 9434
rect 42194 9382 42246 9434
rect 42246 9382 42248 9434
rect 42192 9380 42248 9382
rect 42296 9434 42352 9436
rect 42296 9382 42298 9434
rect 42298 9382 42350 9434
rect 42350 9382 42352 9434
rect 42296 9380 42352 9382
rect 38056 7082 38112 7084
rect 38056 7030 38058 7082
rect 38058 7030 38110 7082
rect 38110 7030 38112 7082
rect 38056 7028 38112 7030
rect 38160 7082 38216 7084
rect 38160 7030 38162 7082
rect 38162 7030 38214 7082
rect 38214 7030 38216 7082
rect 38160 7028 38216 7030
rect 38264 7082 38320 7084
rect 38264 7030 38266 7082
rect 38266 7030 38318 7082
rect 38318 7030 38320 7082
rect 38264 7028 38320 7030
rect 38368 7082 38424 7084
rect 38368 7030 38370 7082
rect 38370 7030 38422 7082
rect 38422 7030 38424 7082
rect 38368 7028 38424 7030
rect 38472 7082 38528 7084
rect 38472 7030 38474 7082
rect 38474 7030 38526 7082
rect 38526 7030 38528 7082
rect 38472 7028 38528 7030
rect 38576 7082 38632 7084
rect 38576 7030 38578 7082
rect 38578 7030 38630 7082
rect 38630 7030 38632 7082
rect 38576 7028 38632 7030
rect 38332 6748 38388 6804
rect 38108 6578 38164 6580
rect 38108 6526 38110 6578
rect 38110 6526 38162 6578
rect 38162 6526 38164 6578
rect 38108 6524 38164 6526
rect 37548 6076 37604 6132
rect 37660 6300 37716 6356
rect 37324 4956 37380 5012
rect 37548 4956 37604 5012
rect 40796 6748 40852 6804
rect 38556 6578 38612 6580
rect 38556 6526 38558 6578
rect 38558 6526 38610 6578
rect 38610 6526 38612 6578
rect 38556 6524 38612 6526
rect 39788 6578 39844 6580
rect 39788 6526 39790 6578
rect 39790 6526 39842 6578
rect 39842 6526 39844 6578
rect 39788 6524 39844 6526
rect 38892 6300 38948 6356
rect 38892 6076 38948 6132
rect 39676 6412 39732 6468
rect 38056 5514 38112 5516
rect 38056 5462 38058 5514
rect 38058 5462 38110 5514
rect 38110 5462 38112 5514
rect 38056 5460 38112 5462
rect 38160 5514 38216 5516
rect 38160 5462 38162 5514
rect 38162 5462 38214 5514
rect 38214 5462 38216 5514
rect 38160 5460 38216 5462
rect 38264 5514 38320 5516
rect 38264 5462 38266 5514
rect 38266 5462 38318 5514
rect 38318 5462 38320 5514
rect 38264 5460 38320 5462
rect 38368 5514 38424 5516
rect 38368 5462 38370 5514
rect 38370 5462 38422 5514
rect 38422 5462 38424 5514
rect 38368 5460 38424 5462
rect 38472 5514 38528 5516
rect 38472 5462 38474 5514
rect 38474 5462 38526 5514
rect 38526 5462 38528 5514
rect 38472 5460 38528 5462
rect 38576 5514 38632 5516
rect 38576 5462 38578 5514
rect 38578 5462 38630 5514
rect 38630 5462 38632 5514
rect 38576 5460 38632 5462
rect 38332 5234 38388 5236
rect 38332 5182 38334 5234
rect 38334 5182 38386 5234
rect 38386 5182 38388 5234
rect 38332 5180 38388 5182
rect 38108 4956 38164 5012
rect 38892 4956 38948 5012
rect 38444 4562 38500 4564
rect 38444 4510 38446 4562
rect 38446 4510 38498 4562
rect 38498 4510 38500 4562
rect 38444 4508 38500 4510
rect 40124 6578 40180 6580
rect 40124 6526 40126 6578
rect 40126 6526 40178 6578
rect 40178 6526 40180 6578
rect 40124 6524 40180 6526
rect 40684 6690 40740 6692
rect 40684 6638 40686 6690
rect 40686 6638 40738 6690
rect 40738 6638 40740 6690
rect 40684 6636 40740 6638
rect 41580 8204 41636 8260
rect 42028 8258 42084 8260
rect 42028 8206 42030 8258
rect 42030 8206 42082 8258
rect 42082 8206 42084 8258
rect 42028 8204 42084 8206
rect 41916 8146 41972 8148
rect 41916 8094 41918 8146
rect 41918 8094 41970 8146
rect 41970 8094 41972 8146
rect 41916 8092 41972 8094
rect 41776 7866 41832 7868
rect 41776 7814 41778 7866
rect 41778 7814 41830 7866
rect 41830 7814 41832 7866
rect 41776 7812 41832 7814
rect 41880 7866 41936 7868
rect 41880 7814 41882 7866
rect 41882 7814 41934 7866
rect 41934 7814 41936 7866
rect 41880 7812 41936 7814
rect 41984 7866 42040 7868
rect 41984 7814 41986 7866
rect 41986 7814 42038 7866
rect 42038 7814 42040 7866
rect 41984 7812 42040 7814
rect 42088 7866 42144 7868
rect 42088 7814 42090 7866
rect 42090 7814 42142 7866
rect 42142 7814 42144 7866
rect 42088 7812 42144 7814
rect 42192 7866 42248 7868
rect 42192 7814 42194 7866
rect 42194 7814 42246 7866
rect 42246 7814 42248 7866
rect 42192 7812 42248 7814
rect 42296 7866 42352 7868
rect 42296 7814 42298 7866
rect 42298 7814 42350 7866
rect 42350 7814 42352 7866
rect 42296 7812 42352 7814
rect 41356 6524 41412 6580
rect 40348 6076 40404 6132
rect 41244 6076 41300 6132
rect 39900 5682 39956 5684
rect 39900 5630 39902 5682
rect 39902 5630 39954 5682
rect 39954 5630 39956 5682
rect 39900 5628 39956 5630
rect 40684 5404 40740 5460
rect 40460 5292 40516 5348
rect 40236 4956 40292 5012
rect 39340 4732 39396 4788
rect 39340 4396 39396 4452
rect 40124 4450 40180 4452
rect 40124 4398 40126 4450
rect 40126 4398 40178 4450
rect 40178 4398 40180 4450
rect 40124 4396 40180 4398
rect 40796 4396 40852 4452
rect 41692 6578 41748 6580
rect 41692 6526 41694 6578
rect 41694 6526 41746 6578
rect 41746 6526 41748 6578
rect 41692 6524 41748 6526
rect 42252 6972 42308 7028
rect 42588 8428 42644 8484
rect 47852 11788 47908 11844
rect 42700 8204 42756 8260
rect 42588 8092 42644 8148
rect 46284 9996 46340 10052
rect 47852 10332 47908 10388
rect 46844 9996 46900 10052
rect 47852 8930 47908 8932
rect 47852 8878 47854 8930
rect 47854 8878 47906 8930
rect 47906 8878 47908 8930
rect 47852 8876 47908 8878
rect 46396 8092 46452 8148
rect 42812 7644 42868 7700
rect 42812 7196 42868 7252
rect 42588 6972 42644 7028
rect 43932 7250 43988 7252
rect 43932 7198 43934 7250
rect 43934 7198 43986 7250
rect 43986 7198 43988 7250
rect 43932 7196 43988 7198
rect 43260 6860 43316 6916
rect 43484 6690 43540 6692
rect 43484 6638 43486 6690
rect 43486 6638 43538 6690
rect 43538 6638 43540 6690
rect 43484 6636 43540 6638
rect 41916 6524 41972 6580
rect 41356 5852 41412 5908
rect 42476 6412 42532 6468
rect 41776 6298 41832 6300
rect 41776 6246 41778 6298
rect 41778 6246 41830 6298
rect 41830 6246 41832 6298
rect 41776 6244 41832 6246
rect 41880 6298 41936 6300
rect 41880 6246 41882 6298
rect 41882 6246 41934 6298
rect 41934 6246 41936 6298
rect 41880 6244 41936 6246
rect 41984 6298 42040 6300
rect 41984 6246 41986 6298
rect 41986 6246 42038 6298
rect 42038 6246 42040 6298
rect 41984 6244 42040 6246
rect 42088 6298 42144 6300
rect 42088 6246 42090 6298
rect 42090 6246 42142 6298
rect 42142 6246 42144 6298
rect 42088 6244 42144 6246
rect 42192 6298 42248 6300
rect 42192 6246 42194 6298
rect 42194 6246 42246 6298
rect 42246 6246 42248 6298
rect 42192 6244 42248 6246
rect 42296 6298 42352 6300
rect 42296 6246 42298 6298
rect 42298 6246 42350 6298
rect 42350 6246 42352 6298
rect 42296 6244 42352 6246
rect 41916 6076 41972 6132
rect 41468 5292 41524 5348
rect 41356 5068 41412 5124
rect 41692 5906 41748 5908
rect 41692 5854 41694 5906
rect 41694 5854 41746 5906
rect 41746 5854 41748 5906
rect 41692 5852 41748 5854
rect 42812 5906 42868 5908
rect 42812 5854 42814 5906
rect 42814 5854 42866 5906
rect 42866 5854 42868 5906
rect 42812 5852 42868 5854
rect 41692 5404 41748 5460
rect 42700 5404 42756 5460
rect 42252 5346 42308 5348
rect 42252 5294 42254 5346
rect 42254 5294 42306 5346
rect 42306 5294 42308 5346
rect 42252 5292 42308 5294
rect 41776 4730 41832 4732
rect 41776 4678 41778 4730
rect 41778 4678 41830 4730
rect 41830 4678 41832 4730
rect 41776 4676 41832 4678
rect 41880 4730 41936 4732
rect 41880 4678 41882 4730
rect 41882 4678 41934 4730
rect 41934 4678 41936 4730
rect 41880 4676 41936 4678
rect 41984 4730 42040 4732
rect 41984 4678 41986 4730
rect 41986 4678 42038 4730
rect 42038 4678 42040 4730
rect 41984 4676 42040 4678
rect 42088 4730 42144 4732
rect 42088 4678 42090 4730
rect 42090 4678 42142 4730
rect 42142 4678 42144 4730
rect 42088 4676 42144 4678
rect 42192 4730 42248 4732
rect 42192 4678 42194 4730
rect 42194 4678 42246 4730
rect 42246 4678 42248 4730
rect 42192 4676 42248 4678
rect 42296 4730 42352 4732
rect 42296 4678 42298 4730
rect 42298 4678 42350 4730
rect 42350 4678 42352 4730
rect 42296 4676 42352 4678
rect 42476 4732 42532 4788
rect 42924 4898 42980 4900
rect 42924 4846 42926 4898
rect 42926 4846 42978 4898
rect 42978 4846 42980 4898
rect 42924 4844 42980 4846
rect 42476 4396 42532 4452
rect 38056 3946 38112 3948
rect 38056 3894 38058 3946
rect 38058 3894 38110 3946
rect 38110 3894 38112 3946
rect 38056 3892 38112 3894
rect 38160 3946 38216 3948
rect 38160 3894 38162 3946
rect 38162 3894 38214 3946
rect 38214 3894 38216 3946
rect 38160 3892 38216 3894
rect 38264 3946 38320 3948
rect 38264 3894 38266 3946
rect 38266 3894 38318 3946
rect 38318 3894 38320 3946
rect 38264 3892 38320 3894
rect 38368 3946 38424 3948
rect 38368 3894 38370 3946
rect 38370 3894 38422 3946
rect 38422 3894 38424 3946
rect 38368 3892 38424 3894
rect 38472 3946 38528 3948
rect 38472 3894 38474 3946
rect 38474 3894 38526 3946
rect 38526 3894 38528 3946
rect 38472 3892 38528 3894
rect 38576 3946 38632 3948
rect 38576 3894 38578 3946
rect 38578 3894 38630 3946
rect 38630 3894 38632 3946
rect 38576 3892 38632 3894
rect 37884 3666 37940 3668
rect 37884 3614 37886 3666
rect 37886 3614 37938 3666
rect 37938 3614 37940 3666
rect 37884 3612 37940 3614
rect 43484 6018 43540 6020
rect 43484 5966 43486 6018
rect 43486 5966 43538 6018
rect 43538 5966 43540 6018
rect 43484 5964 43540 5966
rect 43596 5404 43652 5460
rect 43708 5292 43764 5348
rect 46284 6690 46340 6692
rect 46284 6638 46286 6690
rect 46286 6638 46338 6690
rect 46338 6638 46340 6690
rect 46284 6636 46340 6638
rect 47740 7420 47796 7476
rect 46844 6690 46900 6692
rect 46844 6638 46846 6690
rect 46846 6638 46898 6690
rect 46898 6638 46900 6690
rect 46844 6636 46900 6638
rect 46396 6524 46452 6580
rect 46284 6076 46340 6132
rect 47740 5964 47796 6020
rect 44604 5906 44660 5908
rect 44604 5854 44606 5906
rect 44606 5854 44658 5906
rect 44658 5854 44660 5906
rect 44604 5852 44660 5854
rect 44380 5180 44436 5236
rect 46396 5628 46452 5684
rect 44268 5068 44324 5124
rect 43260 5010 43316 5012
rect 43260 4958 43262 5010
rect 43262 4958 43314 5010
rect 43314 4958 43316 5010
rect 43260 4956 43316 4958
rect 43148 3612 43204 3668
rect 46396 4732 46452 4788
rect 47852 4620 47908 4676
rect 47180 4562 47236 4564
rect 47180 4510 47182 4562
rect 47182 4510 47234 4562
rect 47234 4510 47236 4562
rect 47180 4508 47236 4510
rect 47740 4562 47796 4564
rect 47740 4510 47742 4562
rect 47742 4510 47794 4562
rect 47794 4510 47796 4562
rect 47740 4508 47796 4510
rect 37100 3388 37156 3444
rect 5776 3162 5832 3164
rect 5776 3110 5778 3162
rect 5778 3110 5830 3162
rect 5830 3110 5832 3162
rect 5776 3108 5832 3110
rect 5880 3162 5936 3164
rect 5880 3110 5882 3162
rect 5882 3110 5934 3162
rect 5934 3110 5936 3162
rect 5880 3108 5936 3110
rect 5984 3162 6040 3164
rect 5984 3110 5986 3162
rect 5986 3110 6038 3162
rect 6038 3110 6040 3162
rect 5984 3108 6040 3110
rect 6088 3162 6144 3164
rect 6088 3110 6090 3162
rect 6090 3110 6142 3162
rect 6142 3110 6144 3162
rect 6088 3108 6144 3110
rect 6192 3162 6248 3164
rect 6192 3110 6194 3162
rect 6194 3110 6246 3162
rect 6246 3110 6248 3162
rect 6192 3108 6248 3110
rect 6296 3162 6352 3164
rect 6296 3110 6298 3162
rect 6298 3110 6350 3162
rect 6350 3110 6352 3162
rect 6296 3108 6352 3110
rect 41776 3162 41832 3164
rect 41776 3110 41778 3162
rect 41778 3110 41830 3162
rect 41830 3110 41832 3162
rect 41776 3108 41832 3110
rect 41880 3162 41936 3164
rect 41880 3110 41882 3162
rect 41882 3110 41934 3162
rect 41934 3110 41936 3162
rect 41880 3108 41936 3110
rect 41984 3162 42040 3164
rect 41984 3110 41986 3162
rect 41986 3110 42038 3162
rect 42038 3110 42040 3162
rect 41984 3108 42040 3110
rect 42088 3162 42144 3164
rect 42088 3110 42090 3162
rect 42090 3110 42142 3162
rect 42142 3110 42144 3162
rect 42088 3108 42144 3110
rect 42192 3162 42248 3164
rect 42192 3110 42194 3162
rect 42194 3110 42246 3162
rect 42246 3110 42248 3162
rect 42192 3108 42248 3110
rect 42296 3162 42352 3164
rect 42296 3110 42298 3162
rect 42298 3110 42350 3162
rect 42350 3110 42352 3162
rect 42296 3108 42352 3110
rect 47740 3052 47796 3108
rect 48076 1596 48132 1652
<< metal3 >>
rect 49520 48244 50960 48328
rect 46050 48188 46060 48244
rect 46116 48188 50960 48244
rect 49520 48104 50960 48188
rect 49520 46788 50960 46872
rect 47842 46732 47852 46788
rect 47908 46732 50960 46788
rect 49520 46648 50960 46732
rect -960 46452 480 46648
rect -960 46424 1820 46452
rect 392 46396 1820 46424
rect 1876 46396 1886 46452
rect 2046 46228 2056 46284
rect 2112 46228 2160 46284
rect 2216 46228 2264 46284
rect 2320 46228 2368 46284
rect 2424 46228 2472 46284
rect 2528 46228 2576 46284
rect 2632 46228 2642 46284
rect 38046 46228 38056 46284
rect 38112 46228 38160 46284
rect 38216 46228 38264 46284
rect 38320 46228 38368 46284
rect 38424 46228 38472 46284
rect 38528 46228 38576 46284
rect 38632 46228 38642 46284
rect 5766 45444 5776 45500
rect 5832 45444 5880 45500
rect 5936 45444 5984 45500
rect 6040 45444 6088 45500
rect 6144 45444 6192 45500
rect 6248 45444 6296 45500
rect 6352 45444 6362 45500
rect 41766 45444 41776 45500
rect 41832 45444 41880 45500
rect 41936 45444 41984 45500
rect 42040 45444 42088 45500
rect 42144 45444 42192 45500
rect 42248 45444 42296 45500
rect 42352 45444 42362 45500
rect 49520 45332 50960 45416
rect 47730 45276 47740 45332
rect 47796 45276 50960 45332
rect 49520 45192 50960 45276
rect 2046 44660 2056 44716
rect 2112 44660 2160 44716
rect 2216 44660 2264 44716
rect 2320 44660 2368 44716
rect 2424 44660 2472 44716
rect 2528 44660 2576 44716
rect 2632 44660 2642 44716
rect 38046 44660 38056 44716
rect 38112 44660 38160 44716
rect 38216 44660 38264 44716
rect 38320 44660 38368 44716
rect 38424 44660 38472 44716
rect 38528 44660 38576 44716
rect 38632 44660 38642 44716
rect 5766 43876 5776 43932
rect 5832 43876 5880 43932
rect 5936 43876 5984 43932
rect 6040 43876 6088 43932
rect 6144 43876 6192 43932
rect 6248 43876 6296 43932
rect 6352 43876 6362 43932
rect 41766 43876 41776 43932
rect 41832 43876 41880 43932
rect 41936 43876 41984 43932
rect 42040 43876 42088 43932
rect 42144 43876 42192 43932
rect 42248 43876 42296 43932
rect 42352 43876 42362 43932
rect 49520 43876 50960 43960
rect 47730 43820 47740 43876
rect 47796 43820 50960 43876
rect 49520 43736 50960 43820
rect 2046 43092 2056 43148
rect 2112 43092 2160 43148
rect 2216 43092 2264 43148
rect 2320 43092 2368 43148
rect 2424 43092 2472 43148
rect 2528 43092 2576 43148
rect 2632 43092 2642 43148
rect 38046 43092 38056 43148
rect 38112 43092 38160 43148
rect 38216 43092 38264 43148
rect 38320 43092 38368 43148
rect 38424 43092 38472 43148
rect 38528 43092 38576 43148
rect 38632 43092 38642 43148
rect 49520 42420 50960 42504
rect 47730 42364 47740 42420
rect 47796 42364 50960 42420
rect 5766 42308 5776 42364
rect 5832 42308 5880 42364
rect 5936 42308 5984 42364
rect 6040 42308 6088 42364
rect 6144 42308 6192 42364
rect 6248 42308 6296 42364
rect 6352 42308 6362 42364
rect 41766 42308 41776 42364
rect 41832 42308 41880 42364
rect 41936 42308 41984 42364
rect 42040 42308 42088 42364
rect 42144 42308 42192 42364
rect 42248 42308 42296 42364
rect 42352 42308 42362 42364
rect 49520 42280 50960 42364
rect 40226 41916 40236 41972
rect 40292 41916 46284 41972
rect 46340 41916 46844 41972
rect 46900 41916 46910 41972
rect 2046 41524 2056 41580
rect 2112 41524 2160 41580
rect 2216 41524 2264 41580
rect 2320 41524 2368 41580
rect 2424 41524 2472 41580
rect 2528 41524 2576 41580
rect 2632 41524 2642 41580
rect 38046 41524 38056 41580
rect 38112 41524 38160 41580
rect 38216 41524 38264 41580
rect 38320 41524 38368 41580
rect 38424 41524 38472 41580
rect 38528 41524 38576 41580
rect 38632 41524 38642 41580
rect 49520 40964 50960 41048
rect 3042 40908 3052 40964
rect 3108 40908 3500 40964
rect 3556 40908 17948 40964
rect 18004 40908 18014 40964
rect 47730 40908 47740 40964
rect 47796 40908 50960 40964
rect 49520 40824 50960 40908
rect 5766 40740 5776 40796
rect 5832 40740 5880 40796
rect 5936 40740 5984 40796
rect 6040 40740 6088 40796
rect 6144 40740 6192 40796
rect 6248 40740 6296 40796
rect 6352 40740 6362 40796
rect 41766 40740 41776 40796
rect 41832 40740 41880 40796
rect 41936 40740 41984 40796
rect 42040 40740 42088 40796
rect 42144 40740 42192 40796
rect 42248 40740 42296 40796
rect 42352 40740 42362 40796
rect 392 40488 2156 40516
rect -960 40460 2156 40488
rect 2212 40460 2222 40516
rect -960 40264 480 40460
rect 2046 39956 2056 40012
rect 2112 39956 2160 40012
rect 2216 39956 2264 40012
rect 2320 39956 2368 40012
rect 2424 39956 2472 40012
rect 2528 39956 2576 40012
rect 2632 39956 2642 40012
rect 38046 39956 38056 40012
rect 38112 39956 38160 40012
rect 38216 39956 38264 40012
rect 38320 39956 38368 40012
rect 38424 39956 38472 40012
rect 38528 39956 38576 40012
rect 38632 39956 38642 40012
rect 49520 39508 50960 39592
rect 47730 39452 47740 39508
rect 47796 39452 50960 39508
rect 49520 39368 50960 39452
rect 5766 39172 5776 39228
rect 5832 39172 5880 39228
rect 5936 39172 5984 39228
rect 6040 39172 6088 39228
rect 6144 39172 6192 39228
rect 6248 39172 6296 39228
rect 6352 39172 6362 39228
rect 41766 39172 41776 39228
rect 41832 39172 41880 39228
rect 41936 39172 41984 39228
rect 42040 39172 42088 39228
rect 42144 39172 42192 39228
rect 42248 39172 42296 39228
rect 42352 39172 42362 39228
rect 41122 38668 41132 38724
rect 41188 38668 46396 38724
rect 46452 38668 46844 38724
rect 46900 38668 46910 38724
rect 47842 38668 47852 38724
rect 47908 38668 49588 38724
rect 2046 38388 2056 38444
rect 2112 38388 2160 38444
rect 2216 38388 2264 38444
rect 2320 38388 2368 38444
rect 2424 38388 2472 38444
rect 2528 38388 2576 38444
rect 2632 38388 2642 38444
rect 38046 38388 38056 38444
rect 38112 38388 38160 38444
rect 38216 38388 38264 38444
rect 38320 38388 38368 38444
rect 38424 38388 38472 38444
rect 38528 38388 38576 38444
rect 38632 38388 38642 38444
rect 49532 38276 49588 38668
rect 49308 38220 49588 38276
rect 49308 38052 49364 38220
rect 49520 38052 50960 38136
rect 49308 37996 50960 38052
rect 49520 37912 50960 37996
rect 5766 37604 5776 37660
rect 5832 37604 5880 37660
rect 5936 37604 5984 37660
rect 6040 37604 6088 37660
rect 6144 37604 6192 37660
rect 6248 37604 6296 37660
rect 6352 37604 6362 37660
rect 41766 37604 41776 37660
rect 41832 37604 41880 37660
rect 41936 37604 41984 37660
rect 42040 37604 42088 37660
rect 42144 37604 42192 37660
rect 42248 37604 42296 37660
rect 42352 37604 42362 37660
rect 45602 37100 45612 37156
rect 45668 37100 46396 37156
rect 46452 37100 46844 37156
rect 46900 37100 46910 37156
rect 2046 36820 2056 36876
rect 2112 36820 2160 36876
rect 2216 36820 2264 36876
rect 2320 36820 2368 36876
rect 2424 36820 2472 36876
rect 2528 36820 2576 36876
rect 2632 36820 2642 36876
rect 38046 36820 38056 36876
rect 38112 36820 38160 36876
rect 38216 36820 38264 36876
rect 38320 36820 38368 36876
rect 38424 36820 38472 36876
rect 38528 36820 38576 36876
rect 38632 36820 38642 36876
rect 49520 36596 50960 36680
rect 47842 36540 47852 36596
rect 47908 36540 50960 36596
rect 49520 36456 50960 36540
rect 17378 36316 17388 36372
rect 17444 36316 18284 36372
rect 18340 36316 20188 36372
rect 20132 36260 20188 36316
rect 20132 36204 44156 36260
rect 44212 36204 44222 36260
rect 5766 36036 5776 36092
rect 5832 36036 5880 36092
rect 5936 36036 5984 36092
rect 6040 36036 6088 36092
rect 6144 36036 6192 36092
rect 6248 36036 6296 36092
rect 6352 36036 6362 36092
rect 41766 36036 41776 36092
rect 41832 36036 41880 36092
rect 41936 36036 41984 36092
rect 42040 36036 42088 36092
rect 42144 36036 42192 36092
rect 42248 36036 42296 36092
rect 42352 36036 42362 36092
rect 46386 35644 46396 35700
rect 46452 35644 46956 35700
rect 47012 35644 47022 35700
rect 47842 35308 47852 35364
rect 47908 35308 47918 35364
rect 2046 35252 2056 35308
rect 2112 35252 2160 35308
rect 2216 35252 2264 35308
rect 2320 35252 2368 35308
rect 2424 35252 2472 35308
rect 2528 35252 2576 35308
rect 2632 35252 2642 35308
rect 38046 35252 38056 35308
rect 38112 35252 38160 35308
rect 38216 35252 38264 35308
rect 38320 35252 38368 35308
rect 38424 35252 38472 35308
rect 38528 35252 38576 35308
rect 38632 35252 38642 35308
rect 47852 35140 47908 35308
rect 49520 35140 50960 35224
rect 47852 35084 50960 35140
rect 49520 35000 50960 35084
rect 5766 34468 5776 34524
rect 5832 34468 5880 34524
rect 5936 34468 5984 34524
rect 6040 34468 6088 34524
rect 6144 34468 6192 34524
rect 6248 34468 6296 34524
rect 6352 34468 6362 34524
rect 41766 34468 41776 34524
rect 41832 34468 41880 34524
rect 41936 34468 41984 34524
rect 42040 34468 42088 34524
rect 42144 34468 42192 34524
rect 42248 34468 42296 34524
rect 42352 34468 42362 34524
rect 392 34328 1820 34356
rect -960 34300 1820 34328
rect 1876 34300 1886 34356
rect -960 34104 480 34300
rect 2046 33684 2056 33740
rect 2112 33684 2160 33740
rect 2216 33684 2264 33740
rect 2320 33684 2368 33740
rect 2424 33684 2472 33740
rect 2528 33684 2576 33740
rect 2632 33684 2642 33740
rect 38046 33684 38056 33740
rect 38112 33684 38160 33740
rect 38216 33684 38264 33740
rect 38320 33684 38368 33740
rect 38424 33684 38472 33740
rect 38528 33684 38576 33740
rect 38632 33684 38642 33740
rect 49520 33684 50960 33768
rect 47842 33628 47852 33684
rect 47908 33628 50960 33684
rect 49520 33544 50960 33628
rect 5766 32900 5776 32956
rect 5832 32900 5880 32956
rect 5936 32900 5984 32956
rect 6040 32900 6088 32956
rect 6144 32900 6192 32956
rect 6248 32900 6296 32956
rect 6352 32900 6362 32956
rect 41766 32900 41776 32956
rect 41832 32900 41880 32956
rect 41936 32900 41984 32956
rect 42040 32900 42088 32956
rect 42144 32900 42192 32956
rect 42248 32900 42296 32956
rect 42352 32900 42362 32956
rect 44482 32396 44492 32452
rect 44548 32396 46396 32452
rect 46452 32396 46844 32452
rect 46900 32396 46910 32452
rect 49520 32228 50960 32312
rect 47842 32172 47852 32228
rect 47908 32172 50960 32228
rect 2046 32116 2056 32172
rect 2112 32116 2160 32172
rect 2216 32116 2264 32172
rect 2320 32116 2368 32172
rect 2424 32116 2472 32172
rect 2528 32116 2576 32172
rect 2632 32116 2642 32172
rect 38046 32116 38056 32172
rect 38112 32116 38160 32172
rect 38216 32116 38264 32172
rect 38320 32116 38368 32172
rect 38424 32116 38472 32172
rect 38528 32116 38576 32172
rect 38632 32116 38642 32172
rect 49520 32088 50960 32172
rect 5766 31332 5776 31388
rect 5832 31332 5880 31388
rect 5936 31332 5984 31388
rect 6040 31332 6088 31388
rect 6144 31332 6192 31388
rect 6248 31332 6296 31388
rect 6352 31332 6362 31388
rect 41766 31332 41776 31388
rect 41832 31332 41880 31388
rect 41936 31332 41984 31388
rect 42040 31332 42088 31388
rect 42144 31332 42192 31388
rect 42248 31332 42296 31388
rect 42352 31332 42362 31388
rect 45490 31052 45500 31108
rect 45556 31052 46732 31108
rect 46788 31052 46798 31108
rect 49520 30772 50960 30856
rect 47842 30716 47852 30772
rect 47908 30716 50960 30772
rect 49520 30632 50960 30716
rect 2046 30548 2056 30604
rect 2112 30548 2160 30604
rect 2216 30548 2264 30604
rect 2320 30548 2368 30604
rect 2424 30548 2472 30604
rect 2528 30548 2576 30604
rect 2632 30548 2642 30604
rect 38046 30548 38056 30604
rect 38112 30548 38160 30604
rect 38216 30548 38264 30604
rect 38320 30548 38368 30604
rect 38424 30548 38472 30604
rect 38528 30548 38576 30604
rect 38632 30548 38642 30604
rect 5766 29764 5776 29820
rect 5832 29764 5880 29820
rect 5936 29764 5984 29820
rect 6040 29764 6088 29820
rect 6144 29764 6192 29820
rect 6248 29764 6296 29820
rect 6352 29764 6362 29820
rect 41766 29764 41776 29820
rect 41832 29764 41880 29820
rect 41936 29764 41984 29820
rect 42040 29764 42088 29820
rect 42144 29764 42192 29820
rect 42248 29764 42296 29820
rect 42352 29764 42362 29820
rect 38994 29484 39004 29540
rect 39060 29484 46060 29540
rect 46116 29484 46126 29540
rect 49520 29316 50960 29400
rect 41234 29260 41244 29316
rect 41300 29260 46396 29316
rect 46452 29260 46844 29316
rect 46900 29260 46910 29316
rect 47842 29260 47852 29316
rect 47908 29260 50960 29316
rect 49520 29176 50960 29260
rect 2046 28980 2056 29036
rect 2112 28980 2160 29036
rect 2216 28980 2264 29036
rect 2320 28980 2368 29036
rect 2424 28980 2472 29036
rect 2528 28980 2576 29036
rect 2632 28980 2642 29036
rect 38046 28980 38056 29036
rect 38112 28980 38160 29036
rect 38216 28980 38264 29036
rect 38320 28980 38368 29036
rect 38424 28980 38472 29036
rect 38528 28980 38576 29036
rect 38632 28980 38642 29036
rect 32946 28700 32956 28756
rect 33012 28700 36764 28756
rect 36820 28700 38332 28756
rect 38388 28700 38668 28756
rect 38612 28644 38668 28700
rect 30370 28588 30380 28644
rect 30436 28588 37996 28644
rect 38052 28588 38062 28644
rect 38612 28588 39004 28644
rect 39060 28588 39070 28644
rect 45714 28588 45724 28644
rect 45780 28588 46284 28644
rect 46340 28588 46844 28644
rect 46900 28588 46910 28644
rect 38770 28476 38780 28532
rect 38836 28476 39788 28532
rect 39844 28476 40124 28532
rect 40180 28476 40190 28532
rect 5766 28196 5776 28252
rect 5832 28196 5880 28252
rect 5936 28196 5984 28252
rect 6040 28196 6088 28252
rect 6144 28196 6192 28252
rect 6248 28196 6296 28252
rect 6352 28196 6362 28252
rect 41766 28196 41776 28252
rect 41832 28196 41880 28252
rect 41936 28196 41984 28252
rect 42040 28196 42088 28252
rect 42144 28196 42192 28252
rect 42248 28196 42296 28252
rect 42352 28196 42362 28252
rect -960 28084 480 28168
rect -960 28028 1820 28084
rect 1876 28028 1886 28084
rect 35186 28028 35196 28084
rect 35252 28028 36652 28084
rect 36708 28028 37660 28084
rect 37716 28028 45948 28084
rect 46004 28028 46014 28084
rect -960 27944 480 28028
rect 29474 27916 29484 27972
rect 29540 27916 37884 27972
rect 37940 27916 37950 27972
rect 38210 27916 38220 27972
rect 38276 27916 45836 27972
rect 45892 27916 45902 27972
rect 49520 27860 50960 27944
rect 31490 27804 31500 27860
rect 31556 27804 38108 27860
rect 38164 27804 38556 27860
rect 38612 27804 38780 27860
rect 38836 27804 39116 27860
rect 39172 27804 39182 27860
rect 47842 27804 47852 27860
rect 47908 27804 50960 27860
rect 31602 27692 31612 27748
rect 31668 27692 36204 27748
rect 36260 27692 37436 27748
rect 37492 27692 38220 27748
rect 38276 27692 38286 27748
rect 49520 27720 50960 27804
rect 34626 27580 34636 27636
rect 34692 27580 37324 27636
rect 37380 27580 37390 27636
rect 2046 27412 2056 27468
rect 2112 27412 2160 27468
rect 2216 27412 2264 27468
rect 2320 27412 2368 27468
rect 2424 27412 2472 27468
rect 2528 27412 2576 27468
rect 2632 27412 2642 27468
rect 38046 27412 38056 27468
rect 38112 27412 38160 27468
rect 38216 27412 38264 27468
rect 38320 27412 38368 27468
rect 38424 27412 38472 27468
rect 38528 27412 38576 27468
rect 38632 27412 38642 27468
rect 42802 26908 42812 26964
rect 42868 26908 46284 26964
rect 46340 26908 46844 26964
rect 46900 26908 46910 26964
rect 39778 26796 39788 26852
rect 39844 26796 40236 26852
rect 40292 26796 40796 26852
rect 40852 26796 40862 26852
rect 5766 26628 5776 26684
rect 5832 26628 5880 26684
rect 5936 26628 5984 26684
rect 6040 26628 6088 26684
rect 6144 26628 6192 26684
rect 6248 26628 6296 26684
rect 6352 26628 6362 26684
rect 41766 26628 41776 26684
rect 41832 26628 41880 26684
rect 41936 26628 41984 26684
rect 42040 26628 42088 26684
rect 42144 26628 42192 26684
rect 42248 26628 42296 26684
rect 42352 26628 42362 26684
rect 49520 26404 50960 26488
rect 37090 26348 37100 26404
rect 37156 26348 39116 26404
rect 39172 26348 46620 26404
rect 46676 26348 46686 26404
rect 47730 26348 47740 26404
rect 47796 26348 50960 26404
rect 49520 26264 50960 26348
rect 32386 26124 32396 26180
rect 32452 26124 37548 26180
rect 37604 26124 38556 26180
rect 38612 26124 38892 26180
rect 38948 26124 38958 26180
rect 30034 26012 30044 26068
rect 30100 26012 38220 26068
rect 38276 26012 38286 26068
rect 2046 25844 2056 25900
rect 2112 25844 2160 25900
rect 2216 25844 2264 25900
rect 2320 25844 2368 25900
rect 2424 25844 2472 25900
rect 2528 25844 2576 25900
rect 2632 25844 2642 25900
rect 38046 25844 38056 25900
rect 38112 25844 38160 25900
rect 38216 25844 38264 25900
rect 38320 25844 38368 25900
rect 38424 25844 38472 25900
rect 38528 25844 38576 25900
rect 38632 25844 38642 25900
rect 45826 25676 45836 25732
rect 45892 25676 46956 25732
rect 47012 25676 47022 25732
rect 27906 25340 27916 25396
rect 27972 25340 34636 25396
rect 34692 25340 34702 25396
rect 30818 25228 30828 25284
rect 30884 25228 35196 25284
rect 35252 25228 35262 25284
rect 39666 25228 39676 25284
rect 39732 25228 41132 25284
rect 41188 25228 41198 25284
rect 5766 25060 5776 25116
rect 5832 25060 5880 25116
rect 5936 25060 5984 25116
rect 6040 25060 6088 25116
rect 6144 25060 6192 25116
rect 6248 25060 6296 25116
rect 6352 25060 6362 25116
rect 41766 25060 41776 25116
rect 41832 25060 41880 25116
rect 41936 25060 41984 25116
rect 42040 25060 42088 25116
rect 42144 25060 42192 25116
rect 42248 25060 42296 25116
rect 42352 25060 42362 25116
rect 49520 24948 50960 25032
rect 47730 24892 47740 24948
rect 47796 24892 50960 24948
rect 39106 24780 39116 24836
rect 39172 24780 45500 24836
rect 45556 24780 45566 24836
rect 49520 24808 50960 24892
rect 2046 24276 2056 24332
rect 2112 24276 2160 24332
rect 2216 24276 2264 24332
rect 2320 24276 2368 24332
rect 2424 24276 2472 24332
rect 2528 24276 2576 24332
rect 2632 24276 2642 24332
rect 38046 24276 38056 24332
rect 38112 24276 38160 24332
rect 38216 24276 38264 24332
rect 38320 24276 38368 24332
rect 38424 24276 38472 24332
rect 38528 24276 38576 24332
rect 38632 24276 38642 24332
rect 38612 24108 39116 24164
rect 39172 24108 39182 24164
rect 38612 23940 38668 24108
rect 36978 23884 36988 23940
rect 37044 23884 38332 23940
rect 38388 23884 38668 23940
rect 5766 23492 5776 23548
rect 5832 23492 5880 23548
rect 5936 23492 5984 23548
rect 6040 23492 6088 23548
rect 6144 23492 6192 23548
rect 6248 23492 6296 23548
rect 6352 23492 6362 23548
rect 41766 23492 41776 23548
rect 41832 23492 41880 23548
rect 41936 23492 41984 23548
rect 42040 23492 42088 23548
rect 42144 23492 42192 23548
rect 42248 23492 42296 23548
rect 42352 23492 42362 23548
rect 49520 23492 50960 23576
rect 38322 23436 38332 23492
rect 38388 23436 39004 23492
rect 39060 23436 39676 23492
rect 39732 23436 39742 23492
rect 47730 23436 47740 23492
rect 47796 23436 50960 23492
rect 30482 23324 30492 23380
rect 30548 23324 37884 23380
rect 37940 23324 37950 23380
rect 49520 23352 50960 23436
rect 36866 23212 36876 23268
rect 36932 23212 39004 23268
rect 39060 23212 45612 23268
rect 45668 23212 45678 23268
rect 31826 23100 31836 23156
rect 31892 23100 37996 23156
rect 38052 23100 38062 23156
rect 37314 22876 37324 22932
rect 37380 22876 38332 22932
rect 38388 22876 38398 22932
rect 2046 22708 2056 22764
rect 2112 22708 2160 22764
rect 2216 22708 2264 22764
rect 2320 22708 2368 22764
rect 2424 22708 2472 22764
rect 2528 22708 2576 22764
rect 2632 22708 2642 22764
rect 38046 22708 38056 22764
rect 38112 22708 38160 22764
rect 38216 22708 38264 22764
rect 38320 22708 38368 22764
rect 38424 22708 38472 22764
rect 38528 22708 38576 22764
rect 38632 22708 38642 22764
rect 12898 22204 12908 22260
rect 12964 22204 38108 22260
rect 38164 22204 38668 22260
rect 38724 22204 38734 22260
rect 16370 22092 16380 22148
rect 16436 22092 28028 22148
rect 28084 22092 28094 22148
rect 34962 22092 34972 22148
rect 35028 22092 46284 22148
rect 46340 22092 46844 22148
rect 46900 22092 46910 22148
rect 49520 22036 50960 22120
rect 392 22008 1820 22036
rect -960 21980 1820 22008
rect 1876 21980 1886 22036
rect 47730 21980 47740 22036
rect 47796 21980 50960 22036
rect -960 21784 480 21980
rect 5766 21924 5776 21980
rect 5832 21924 5880 21980
rect 5936 21924 5984 21980
rect 6040 21924 6088 21980
rect 6144 21924 6192 21980
rect 6248 21924 6296 21980
rect 6352 21924 6362 21980
rect 41766 21924 41776 21980
rect 41832 21924 41880 21980
rect 41936 21924 41984 21980
rect 42040 21924 42088 21980
rect 42144 21924 42192 21980
rect 42248 21924 42296 21980
rect 42352 21924 42362 21980
rect 28018 21868 28028 21924
rect 28084 21868 37324 21924
rect 37380 21868 37390 21924
rect 49520 21896 50960 21980
rect 33394 21756 33404 21812
rect 33460 21756 37436 21812
rect 37492 21756 37502 21812
rect 38658 21532 38668 21588
rect 38724 21532 40348 21588
rect 40404 21532 40414 21588
rect 20514 21420 20524 21476
rect 20580 21420 36428 21476
rect 36484 21420 36764 21476
rect 36820 21420 38444 21476
rect 38500 21420 38510 21476
rect 22418 21308 22428 21364
rect 22484 21308 36876 21364
rect 36932 21308 37884 21364
rect 37940 21308 37950 21364
rect 38210 21308 38220 21364
rect 38276 21308 39900 21364
rect 39956 21308 39966 21364
rect 2046 21140 2056 21196
rect 2112 21140 2160 21196
rect 2216 21140 2264 21196
rect 2320 21140 2368 21196
rect 2424 21140 2472 21196
rect 2528 21140 2576 21196
rect 2632 21140 2642 21196
rect 38046 21140 38056 21196
rect 38112 21140 38160 21196
rect 38216 21140 38264 21196
rect 38320 21140 38368 21196
rect 38424 21140 38472 21196
rect 38528 21140 38576 21196
rect 38632 21140 38642 21196
rect 28354 20972 28364 21028
rect 28420 20972 29820 21028
rect 29876 20972 29886 21028
rect 36754 20972 36764 21028
rect 36820 20972 37996 21028
rect 38052 20972 38062 21028
rect 38322 20972 38332 21028
rect 38388 20972 38668 21028
rect 38724 20972 46060 21028
rect 46116 20972 46126 21028
rect 37996 20916 38052 20972
rect 37996 20860 47068 20916
rect 47124 20860 47134 20916
rect 34290 20636 34300 20692
rect 34356 20636 39452 20692
rect 39508 20636 39518 20692
rect 40002 20636 40012 20692
rect 40068 20636 40796 20692
rect 40852 20636 41580 20692
rect 41636 20636 41646 20692
rect 49520 20580 50960 20664
rect 17378 20524 17388 20580
rect 17444 20524 28812 20580
rect 28868 20524 30156 20580
rect 30212 20524 30222 20580
rect 32162 20524 32172 20580
rect 32228 20524 37660 20580
rect 37716 20524 37726 20580
rect 39106 20524 39116 20580
rect 39172 20524 39676 20580
rect 39732 20524 39742 20580
rect 47730 20524 47740 20580
rect 47796 20524 50960 20580
rect 49520 20440 50960 20524
rect 5766 20356 5776 20412
rect 5832 20356 5880 20412
rect 5936 20356 5984 20412
rect 6040 20356 6088 20412
rect 6144 20356 6192 20412
rect 6248 20356 6296 20412
rect 6352 20356 6362 20412
rect 41766 20356 41776 20412
rect 41832 20356 41880 20412
rect 41936 20356 41984 20412
rect 42040 20356 42088 20412
rect 42144 20356 42192 20412
rect 42248 20356 42296 20412
rect 42352 20356 42362 20412
rect 22642 20188 22652 20244
rect 22708 20188 33628 20244
rect 33684 20188 33694 20244
rect 36418 20188 36428 20244
rect 36484 20188 37436 20244
rect 37492 20188 38332 20244
rect 38388 20188 38398 20244
rect 29362 20076 29372 20132
rect 29428 20076 30828 20132
rect 30884 20076 30894 20132
rect 37986 20076 37996 20132
rect 38052 20076 44492 20132
rect 44548 20076 44558 20132
rect 29372 19908 29428 20076
rect 38210 19964 38220 20020
rect 38276 19964 38780 20020
rect 38836 19964 38846 20020
rect 25666 19852 25676 19908
rect 25732 19852 29428 19908
rect 23650 19740 23660 19796
rect 23716 19740 35980 19796
rect 36036 19740 36764 19796
rect 36820 19740 36830 19796
rect 2046 19572 2056 19628
rect 2112 19572 2160 19628
rect 2216 19572 2264 19628
rect 2320 19572 2368 19628
rect 2424 19572 2472 19628
rect 2528 19572 2576 19628
rect 2632 19572 2642 19628
rect 38046 19572 38056 19628
rect 38112 19572 38160 19628
rect 38216 19572 38264 19628
rect 38320 19572 38368 19628
rect 38424 19572 38472 19628
rect 38528 19572 38576 19628
rect 38632 19572 38642 19628
rect 36754 19404 36764 19460
rect 36820 19404 37996 19460
rect 38052 19404 38062 19460
rect 19730 19292 19740 19348
rect 19796 19292 36428 19348
rect 36484 19292 36494 19348
rect 49520 19124 50960 19208
rect 31266 19068 31276 19124
rect 31332 19068 37660 19124
rect 37716 19068 37726 19124
rect 38770 19068 38780 19124
rect 38836 19068 45836 19124
rect 45892 19068 45902 19124
rect 47730 19068 47740 19124
rect 47796 19068 50960 19124
rect 14466 18956 14476 19012
rect 14532 18956 34188 19012
rect 34244 18956 34860 19012
rect 34916 18956 34926 19012
rect 36194 18956 36204 19012
rect 36260 18956 37324 19012
rect 37380 18956 41244 19012
rect 41300 18956 41310 19012
rect 49520 18984 50960 19068
rect 33730 18844 33740 18900
rect 33796 18844 34300 18900
rect 34356 18844 34366 18900
rect 5766 18788 5776 18844
rect 5832 18788 5880 18844
rect 5936 18788 5984 18844
rect 6040 18788 6088 18844
rect 6144 18788 6192 18844
rect 6248 18788 6296 18844
rect 6352 18788 6362 18844
rect 41766 18788 41776 18844
rect 41832 18788 41880 18844
rect 41936 18788 41984 18844
rect 42040 18788 42088 18844
rect 42144 18788 42192 18844
rect 42248 18788 42296 18844
rect 42352 18788 42362 18844
rect 35746 18732 35756 18788
rect 35812 18732 36764 18788
rect 36820 18732 38108 18788
rect 38164 18732 38780 18788
rect 38836 18732 38846 18788
rect 33506 18620 33516 18676
rect 33572 18620 37212 18676
rect 37268 18620 37278 18676
rect 31266 18508 31276 18564
rect 31332 18508 37100 18564
rect 37156 18508 37166 18564
rect 37314 18508 37324 18564
rect 37380 18508 37660 18564
rect 37716 18508 37726 18564
rect 26852 18396 34860 18452
rect 34916 18396 34926 18452
rect 35074 18396 35084 18452
rect 35140 18396 35644 18452
rect 35700 18396 35710 18452
rect 36642 18396 36652 18452
rect 36708 18396 37548 18452
rect 37604 18396 38556 18452
rect 38612 18396 38780 18452
rect 38836 18396 40348 18452
rect 40404 18396 40414 18452
rect 26852 18340 26908 18396
rect 20850 18284 20860 18340
rect 20916 18284 26908 18340
rect 32610 18284 32620 18340
rect 32676 18284 36428 18340
rect 36484 18284 36494 18340
rect 35410 18060 35420 18116
rect 35476 18060 36204 18116
rect 36260 18060 36270 18116
rect 2046 18004 2056 18060
rect 2112 18004 2160 18060
rect 2216 18004 2264 18060
rect 2320 18004 2368 18060
rect 2424 18004 2472 18060
rect 2528 18004 2576 18060
rect 2632 18004 2642 18060
rect 38046 18004 38056 18060
rect 38112 18004 38160 18060
rect 38216 18004 38264 18060
rect 38320 18004 38368 18060
rect 38424 18004 38472 18060
rect 38528 18004 38576 18060
rect 38632 18004 38642 18060
rect 33954 17948 33964 18004
rect 34020 17948 35532 18004
rect 35588 17948 35598 18004
rect 34738 17836 34748 17892
rect 34804 17836 35420 17892
rect 35476 17836 35486 17892
rect 31602 17724 31612 17780
rect 31668 17724 32060 17780
rect 32116 17724 37436 17780
rect 37492 17724 37502 17780
rect 49520 17668 50960 17752
rect 29698 17612 29708 17668
rect 29764 17612 30380 17668
rect 30436 17612 30446 17668
rect 34850 17612 34860 17668
rect 34916 17612 35868 17668
rect 35924 17612 35934 17668
rect 36418 17612 36428 17668
rect 36484 17612 42812 17668
rect 42868 17612 42878 17668
rect 47842 17612 47852 17668
rect 47908 17612 50960 17668
rect 35298 17500 35308 17556
rect 35364 17500 37884 17556
rect 37940 17500 37950 17556
rect 49520 17528 50960 17612
rect 35634 17388 35644 17444
rect 35700 17388 46060 17444
rect 46116 17388 46126 17444
rect 5766 17220 5776 17276
rect 5832 17220 5880 17276
rect 5936 17220 5984 17276
rect 6040 17220 6088 17276
rect 6144 17220 6192 17276
rect 6248 17220 6296 17276
rect 6352 17220 6362 17276
rect 41766 17220 41776 17276
rect 41832 17220 41880 17276
rect 41936 17220 41984 17276
rect 42040 17220 42088 17276
rect 42144 17220 42192 17276
rect 42248 17220 42296 17276
rect 42352 17220 42362 17276
rect 35858 17164 35868 17220
rect 35924 17164 37436 17220
rect 37492 17164 38220 17220
rect 38276 17164 38668 17220
rect 38612 17108 38668 17164
rect 31490 17052 31500 17108
rect 31556 17052 32060 17108
rect 32116 17052 37772 17108
rect 37828 17052 37838 17108
rect 38612 17052 45724 17108
rect 45780 17052 45790 17108
rect 34290 16940 34300 16996
rect 34356 16940 36316 16996
rect 36372 16940 46956 16996
rect 47012 16940 47022 16996
rect 15474 16828 15484 16884
rect 15540 16828 17388 16884
rect 17444 16828 17454 16884
rect 33954 16828 33964 16884
rect 34020 16828 34860 16884
rect 34916 16828 35756 16884
rect 35812 16828 36428 16884
rect 36484 16828 36494 16884
rect 39442 16828 39452 16884
rect 39508 16828 46396 16884
rect 46452 16828 46844 16884
rect 46900 16828 46910 16884
rect 47730 16828 47740 16884
rect 47796 16828 49588 16884
rect 2046 16436 2056 16492
rect 2112 16436 2160 16492
rect 2216 16436 2264 16492
rect 2320 16436 2368 16492
rect 2424 16436 2472 16492
rect 2528 16436 2576 16492
rect 2632 16436 2642 16492
rect 38046 16436 38056 16492
rect 38112 16436 38160 16492
rect 38216 16436 38264 16492
rect 38320 16436 38368 16492
rect 38424 16436 38472 16492
rect 38528 16436 38576 16492
rect 38632 16436 38642 16492
rect 49532 16436 49588 16828
rect 30930 16380 30940 16436
rect 30996 16380 31052 16436
rect 31108 16380 31118 16436
rect 49308 16380 49588 16436
rect 29922 16268 29932 16324
rect 29988 16268 30380 16324
rect 30436 16268 30446 16324
rect 49308 16212 49364 16380
rect 49520 16212 50960 16296
rect 49308 16156 50960 16212
rect 28466 16044 28476 16100
rect 28532 16044 32844 16100
rect 32900 16044 33516 16100
rect 33572 16044 34188 16100
rect 34244 16044 34972 16100
rect 35028 16044 45948 16100
rect 46004 16044 46014 16100
rect 49520 16072 50960 16156
rect 31378 15932 31388 15988
rect 31444 15932 31836 15988
rect 31892 15932 31902 15988
rect 37874 15932 37884 15988
rect 37940 15932 40012 15988
rect 40068 15932 40078 15988
rect -960 15652 480 15848
rect 23762 15820 23772 15876
rect 23828 15820 27132 15876
rect 27188 15820 27198 15876
rect 28242 15820 28252 15876
rect 28308 15820 31052 15876
rect 31108 15820 31118 15876
rect 28914 15708 28924 15764
rect 28980 15708 33292 15764
rect 33348 15708 34300 15764
rect 34356 15708 34748 15764
rect 34804 15708 34814 15764
rect 5766 15652 5776 15708
rect 5832 15652 5880 15708
rect 5936 15652 5984 15708
rect 6040 15652 6088 15708
rect 6144 15652 6192 15708
rect 6248 15652 6296 15708
rect 6352 15652 6362 15708
rect 41766 15652 41776 15708
rect 41832 15652 41880 15708
rect 41936 15652 41984 15708
rect 42040 15652 42088 15708
rect 42144 15652 42192 15708
rect 42248 15652 42296 15708
rect 42352 15652 42362 15708
rect -960 15624 1820 15652
rect 392 15596 1820 15624
rect 1876 15596 1886 15652
rect 24994 15596 25004 15652
rect 25060 15596 37436 15652
rect 37492 15596 37660 15652
rect 37716 15596 37726 15652
rect 31014 15484 31052 15540
rect 31108 15484 31118 15540
rect 34290 15484 34300 15540
rect 34356 15484 34860 15540
rect 34916 15484 34926 15540
rect 39106 15484 39116 15540
rect 39172 15484 40796 15540
rect 40852 15484 40862 15540
rect 29138 15372 29148 15428
rect 29204 15372 30044 15428
rect 30100 15372 30110 15428
rect 38882 15372 38892 15428
rect 38948 15372 39340 15428
rect 39396 15372 39406 15428
rect 34402 15260 34412 15316
rect 34468 15260 34748 15316
rect 34804 15260 35644 15316
rect 35700 15260 36876 15316
rect 36932 15260 40012 15316
rect 40068 15260 40078 15316
rect 41458 15260 41468 15316
rect 41524 15260 46284 15316
rect 46340 15260 46844 15316
rect 46900 15260 46910 15316
rect 41468 15204 41524 15260
rect 38210 15148 38220 15204
rect 38276 15148 39340 15204
rect 39396 15148 41524 15204
rect 35522 15036 35532 15092
rect 35588 15036 35756 15092
rect 35812 15036 36428 15092
rect 36484 15036 36494 15092
rect 37650 15036 37660 15092
rect 37716 15036 37996 15092
rect 38052 15036 38062 15092
rect 38770 15036 38780 15092
rect 38836 15036 39452 15092
rect 39508 15036 39518 15092
rect 36194 14924 36204 14980
rect 36260 14924 36988 14980
rect 37044 14924 37054 14980
rect 2046 14868 2056 14924
rect 2112 14868 2160 14924
rect 2216 14868 2264 14924
rect 2320 14868 2368 14924
rect 2424 14868 2472 14924
rect 2528 14868 2576 14924
rect 2632 14868 2642 14924
rect 38046 14868 38056 14924
rect 38112 14868 38160 14924
rect 38216 14868 38264 14924
rect 38320 14868 38368 14924
rect 38424 14868 38472 14924
rect 38528 14868 38576 14924
rect 38632 14868 38642 14924
rect 38780 14756 38836 15036
rect 49520 14756 50960 14840
rect 31892 14700 33292 14756
rect 33348 14700 33740 14756
rect 33796 14700 34300 14756
rect 34356 14700 34860 14756
rect 34916 14700 34926 14756
rect 36082 14700 36092 14756
rect 36148 14700 36764 14756
rect 36820 14700 37324 14756
rect 37380 14700 38836 14756
rect 47842 14700 47852 14756
rect 47908 14700 50960 14756
rect 31892 14644 31948 14700
rect 30034 14588 30044 14644
rect 30100 14588 31948 14644
rect 36978 14588 36988 14644
rect 37044 14588 38444 14644
rect 38500 14588 46172 14644
rect 46228 14588 46238 14644
rect 49520 14616 50960 14700
rect 37650 14364 37660 14420
rect 37716 14364 38108 14420
rect 38164 14364 40012 14420
rect 40068 14364 40572 14420
rect 40628 14364 40638 14420
rect 35970 14252 35980 14308
rect 36036 14252 39676 14308
rect 39732 14252 39742 14308
rect 41580 14252 46508 14308
rect 46564 14252 46574 14308
rect 41580 14196 41636 14252
rect 37874 14140 37884 14196
rect 37940 14140 41636 14196
rect 5766 14084 5776 14140
rect 5832 14084 5880 14140
rect 5936 14084 5984 14140
rect 6040 14084 6088 14140
rect 6144 14084 6192 14140
rect 6248 14084 6296 14140
rect 6352 14084 6362 14140
rect 41766 14084 41776 14140
rect 41832 14084 41880 14140
rect 41936 14084 41984 14140
rect 42040 14084 42088 14140
rect 42144 14084 42192 14140
rect 42248 14084 42296 14140
rect 42352 14084 42362 14140
rect 38994 13916 39004 13972
rect 39060 13916 39900 13972
rect 39956 13916 39966 13972
rect 28802 13692 28812 13748
rect 28868 13692 34132 13748
rect 40114 13692 40124 13748
rect 40180 13692 40684 13748
rect 40740 13692 42476 13748
rect 42532 13692 46284 13748
rect 46340 13692 46844 13748
rect 46900 13692 46910 13748
rect 34076 13636 34132 13692
rect 34066 13580 34076 13636
rect 34132 13580 35532 13636
rect 35588 13580 35598 13636
rect 29474 13468 29484 13524
rect 29540 13468 30492 13524
rect 30548 13468 30558 13524
rect 32610 13468 32620 13524
rect 32676 13468 36204 13524
rect 36260 13468 36428 13524
rect 36484 13468 36494 13524
rect 47842 13468 47852 13524
rect 47908 13468 47918 13524
rect 2046 13300 2056 13356
rect 2112 13300 2160 13356
rect 2216 13300 2264 13356
rect 2320 13300 2368 13356
rect 2424 13300 2472 13356
rect 2528 13300 2576 13356
rect 2632 13300 2642 13356
rect 38046 13300 38056 13356
rect 38112 13300 38160 13356
rect 38216 13300 38264 13356
rect 38320 13300 38368 13356
rect 38424 13300 38472 13356
rect 38528 13300 38576 13356
rect 38632 13300 38642 13356
rect 47852 13300 47908 13468
rect 49520 13300 50960 13384
rect 47852 13244 50960 13300
rect 38546 13132 38556 13188
rect 38612 13132 39340 13188
rect 39396 13132 39406 13188
rect 49520 13160 50960 13244
rect 19058 13020 19068 13076
rect 19124 13020 23660 13076
rect 23716 13020 23726 13076
rect 16930 12796 16940 12852
rect 16996 12796 19628 12852
rect 19684 12796 20188 12852
rect 41906 12796 41916 12852
rect 41972 12796 42700 12852
rect 42756 12796 42766 12852
rect 20132 12740 20188 12796
rect 20132 12684 30940 12740
rect 30996 12684 31006 12740
rect 36082 12684 36092 12740
rect 36148 12684 36652 12740
rect 36708 12684 37436 12740
rect 37492 12684 37502 12740
rect 5766 12516 5776 12572
rect 5832 12516 5880 12572
rect 5936 12516 5984 12572
rect 6040 12516 6088 12572
rect 6144 12516 6192 12572
rect 6248 12516 6296 12572
rect 6352 12516 6362 12572
rect 41766 12516 41776 12572
rect 41832 12516 41880 12572
rect 41936 12516 41984 12572
rect 42040 12516 42088 12572
rect 42144 12516 42192 12572
rect 42248 12516 42296 12572
rect 42352 12516 42362 12572
rect 18386 12348 18396 12404
rect 18452 12348 20748 12404
rect 20804 12348 31836 12404
rect 31892 12348 31902 12404
rect 40786 12348 40796 12404
rect 40852 12348 40862 12404
rect 31826 12124 31836 12180
rect 31892 12124 32732 12180
rect 32788 12124 32798 12180
rect 40796 12068 40852 12348
rect 42578 12236 42588 12292
rect 42644 12236 43372 12292
rect 43428 12236 46284 12292
rect 46340 12236 46844 12292
rect 46900 12236 46910 12292
rect 40796 12012 41692 12068
rect 41748 12012 41758 12068
rect 49520 11844 50960 11928
rect 38780 11788 40348 11844
rect 40404 11788 40414 11844
rect 41122 11788 41132 11844
rect 41188 11788 42028 11844
rect 42084 11788 42094 11844
rect 47842 11788 47852 11844
rect 47908 11788 50960 11844
rect 2046 11732 2056 11788
rect 2112 11732 2160 11788
rect 2216 11732 2264 11788
rect 2320 11732 2368 11788
rect 2424 11732 2472 11788
rect 2528 11732 2576 11788
rect 2632 11732 2642 11788
rect 38046 11732 38056 11788
rect 38112 11732 38160 11788
rect 38216 11732 38264 11788
rect 38320 11732 38368 11788
rect 38424 11732 38472 11788
rect 38528 11732 38576 11788
rect 38632 11732 38642 11788
rect 32498 11676 32508 11732
rect 32564 11676 33404 11732
rect 33460 11676 33470 11732
rect 38780 11620 38836 11788
rect 41132 11732 41188 11788
rect 40450 11676 40460 11732
rect 40516 11676 41188 11732
rect 49520 11704 50960 11788
rect 38322 11564 38332 11620
rect 38388 11564 38836 11620
rect 21634 11452 21644 11508
rect 21700 11452 25676 11508
rect 25732 11452 25742 11508
rect 25890 11452 25900 11508
rect 25956 11452 28588 11508
rect 28644 11452 31164 11508
rect 31220 11452 31230 11508
rect 33842 11452 33852 11508
rect 33908 11452 36540 11508
rect 36596 11452 39564 11508
rect 39620 11452 39630 11508
rect 24546 11340 24556 11396
rect 24612 11340 24780 11396
rect 24836 11340 25116 11396
rect 25172 11340 27468 11396
rect 27524 11340 27916 11396
rect 27972 11340 28364 11396
rect 28420 11340 29596 11396
rect 29652 11340 29662 11396
rect 34066 11340 34076 11396
rect 34132 11340 35308 11396
rect 35364 11340 37212 11396
rect 37268 11340 37278 11396
rect 37650 11340 37660 11396
rect 37716 11340 40684 11396
rect 40740 11340 40750 11396
rect 34076 11284 34132 11340
rect 33170 11228 33180 11284
rect 33236 11228 34132 11284
rect 36530 11228 36540 11284
rect 36596 11228 40572 11284
rect 40628 11228 40638 11284
rect 41458 11228 41468 11284
rect 41524 11228 42364 11284
rect 42420 11228 42430 11284
rect 16930 11004 16940 11060
rect 16996 11004 35420 11060
rect 35476 11004 35486 11060
rect 5766 10948 5776 11004
rect 5832 10948 5880 11004
rect 5936 10948 5984 11004
rect 6040 10948 6088 11004
rect 6144 10948 6192 11004
rect 6248 10948 6296 11004
rect 6352 10948 6362 11004
rect 41766 10948 41776 11004
rect 41832 10948 41880 11004
rect 41936 10948 41984 11004
rect 42040 10948 42088 11004
rect 42144 10948 42192 11004
rect 42248 10948 42296 11004
rect 42352 10948 42362 11004
rect 20290 10780 20300 10836
rect 20356 10780 22876 10836
rect 22932 10780 31276 10836
rect 31332 10780 31342 10836
rect 2818 10668 2828 10724
rect 2884 10668 4172 10724
rect 4228 10668 4238 10724
rect 14802 10668 14812 10724
rect 14868 10668 17612 10724
rect 17668 10668 32284 10724
rect 32340 10668 32350 10724
rect 34626 10668 34636 10724
rect 34692 10668 37660 10724
rect 37716 10668 37726 10724
rect 30370 10556 30380 10612
rect 30436 10556 36876 10612
rect 36932 10556 36942 10612
rect 38770 10444 38780 10500
rect 38836 10444 40796 10500
rect 40852 10444 42028 10500
rect 42084 10444 42476 10500
rect 42532 10444 42542 10500
rect 49520 10388 50960 10472
rect 47842 10332 47852 10388
rect 47908 10332 50960 10388
rect 49520 10248 50960 10332
rect 2046 10164 2056 10220
rect 2112 10164 2160 10220
rect 2216 10164 2264 10220
rect 2320 10164 2368 10220
rect 2424 10164 2472 10220
rect 2528 10164 2576 10220
rect 2632 10164 2642 10220
rect 38046 10164 38056 10220
rect 38112 10164 38160 10220
rect 38216 10164 38264 10220
rect 38320 10164 38368 10220
rect 38424 10164 38472 10220
rect 38528 10164 38576 10220
rect 38632 10164 38642 10220
rect 21634 9996 21644 10052
rect 21700 9996 22652 10052
rect 22708 9996 22718 10052
rect 42578 9996 42588 10052
rect 42644 9996 46284 10052
rect 46340 9996 46844 10052
rect 46900 9996 46910 10052
rect 13458 9884 13468 9940
rect 13524 9884 15596 9940
rect 15652 9884 16044 9940
rect 16100 9884 16604 9940
rect 16660 9884 17052 9940
rect 17108 9884 18956 9940
rect 19012 9884 19022 9940
rect 31892 9884 32956 9940
rect 33012 9884 33516 9940
rect 33572 9884 33582 9940
rect 29922 9772 29932 9828
rect 29988 9772 30828 9828
rect 30884 9772 31836 9828
rect 31892 9772 31948 9884
rect -960 9492 480 9688
rect 17378 9660 17388 9716
rect 17444 9660 20076 9716
rect 20132 9660 31052 9716
rect 31108 9660 31118 9716
rect 2146 9548 2156 9604
rect 2212 9548 3612 9604
rect 3668 9548 5628 9604
rect 5684 9548 6860 9604
rect 6916 9548 6926 9604
rect 37538 9548 37548 9604
rect 37604 9548 42140 9604
rect 42196 9548 42206 9604
rect -960 9464 1820 9492
rect 392 9436 1820 9464
rect 1876 9436 1886 9492
rect 5766 9380 5776 9436
rect 5832 9380 5880 9436
rect 5936 9380 5984 9436
rect 6040 9380 6088 9436
rect 6144 9380 6192 9436
rect 6248 9380 6296 9436
rect 6352 9380 6362 9436
rect 41766 9380 41776 9436
rect 41832 9380 41880 9436
rect 41936 9380 41984 9436
rect 42040 9380 42088 9436
rect 42144 9380 42192 9436
rect 42248 9380 42296 9436
rect 42352 9380 42362 9436
rect 33506 9324 33516 9380
rect 33572 9324 39788 9380
rect 39844 9324 39854 9380
rect 19954 9212 19964 9268
rect 20020 9212 25004 9268
rect 25060 9212 25070 9268
rect 33954 9212 33964 9268
rect 34020 9212 35196 9268
rect 35252 9212 35756 9268
rect 35812 9212 35822 9268
rect 2930 9100 2940 9156
rect 2996 9100 4284 9156
rect 4340 9100 4350 9156
rect 3042 8988 3052 9044
rect 3108 8988 19180 9044
rect 19236 8988 19628 9044
rect 19684 8988 19694 9044
rect 49520 8932 50960 9016
rect 6850 8876 6860 8932
rect 6916 8876 11788 8932
rect 11844 8876 12572 8932
rect 12628 8876 13468 8932
rect 13524 8876 13534 8932
rect 16706 8876 16716 8932
rect 16772 8876 17724 8932
rect 17780 8876 23436 8932
rect 23492 8876 23502 8932
rect 30706 8876 30716 8932
rect 30772 8876 33516 8932
rect 33572 8876 33582 8932
rect 47842 8876 47852 8932
rect 47908 8876 50960 8932
rect 49520 8792 50960 8876
rect 2046 8596 2056 8652
rect 2112 8596 2160 8652
rect 2216 8596 2264 8652
rect 2320 8596 2368 8652
rect 2424 8596 2472 8652
rect 2528 8596 2576 8652
rect 2632 8596 2642 8652
rect 38046 8596 38056 8652
rect 38112 8596 38160 8652
rect 38216 8596 38264 8652
rect 38320 8596 38368 8652
rect 38424 8596 38472 8652
rect 38528 8596 38576 8652
rect 38632 8596 38642 8652
rect 38546 8428 38556 8484
rect 38612 8428 41132 8484
rect 41188 8428 42588 8484
rect 42644 8428 42654 8484
rect 8642 8316 8652 8372
rect 8708 8316 13020 8372
rect 13076 8316 13086 8372
rect 4946 8204 4956 8260
rect 5012 8204 5628 8260
rect 5684 8204 5694 8260
rect 8978 8204 8988 8260
rect 9044 8204 9660 8260
rect 9716 8204 9996 8260
rect 10052 8204 10062 8260
rect 41570 8204 41580 8260
rect 41636 8204 42028 8260
rect 42084 8204 42700 8260
rect 42756 8204 42766 8260
rect 2034 8092 2044 8148
rect 2100 8092 9548 8148
rect 9604 8092 10780 8148
rect 10836 8092 38892 8148
rect 38948 8092 38958 8148
rect 40674 8092 40684 8148
rect 40740 8092 41916 8148
rect 41972 8092 42588 8148
rect 42644 8092 46396 8148
rect 46452 8092 46462 8148
rect 13570 7980 13580 8036
rect 13636 7980 16492 8036
rect 16548 7980 17052 8036
rect 17108 7980 17388 8036
rect 17444 7980 17454 8036
rect 17826 7980 17836 8036
rect 17892 7980 20524 8036
rect 20580 7980 33180 8036
rect 33236 7980 33246 8036
rect 5766 7812 5776 7868
rect 5832 7812 5880 7868
rect 5936 7812 5984 7868
rect 6040 7812 6088 7868
rect 6144 7812 6192 7868
rect 6248 7812 6296 7868
rect 6352 7812 6362 7868
rect 41766 7812 41776 7868
rect 41832 7812 41880 7868
rect 41936 7812 41984 7868
rect 42040 7812 42088 7868
rect 42144 7812 42192 7868
rect 42248 7812 42296 7868
rect 42352 7812 42362 7868
rect 36418 7644 36428 7700
rect 36484 7644 39004 7700
rect 39060 7644 42812 7700
rect 42868 7644 42878 7700
rect 6402 7532 6412 7588
rect 6468 7532 6860 7588
rect 6916 7532 6926 7588
rect 49520 7476 50960 7560
rect 23426 7420 23436 7476
rect 23492 7420 24444 7476
rect 24500 7420 26236 7476
rect 26292 7420 28252 7476
rect 28308 7420 29148 7476
rect 29204 7420 29214 7476
rect 47730 7420 47740 7476
rect 47796 7420 50960 7476
rect 5170 7308 5180 7364
rect 5236 7308 5628 7364
rect 5684 7308 6188 7364
rect 6244 7308 9660 7364
rect 9716 7308 11788 7364
rect 11844 7308 13580 7364
rect 13636 7308 13646 7364
rect 49520 7336 50960 7420
rect 22866 7196 22876 7252
rect 22932 7196 42812 7252
rect 42868 7196 43932 7252
rect 43988 7196 43998 7252
rect 2046 7028 2056 7084
rect 2112 7028 2160 7084
rect 2216 7028 2264 7084
rect 2320 7028 2368 7084
rect 2424 7028 2472 7084
rect 2528 7028 2576 7084
rect 2632 7028 2642 7084
rect 38046 7028 38056 7084
rect 38112 7028 38160 7084
rect 38216 7028 38264 7084
rect 38320 7028 38368 7084
rect 38424 7028 38472 7084
rect 38528 7028 38576 7084
rect 38632 7028 38642 7084
rect 42242 6972 42252 7028
rect 42308 6972 42588 7028
rect 42644 6972 42654 7028
rect 20290 6860 20300 6916
rect 20356 6860 43260 6916
rect 43316 6860 43326 6916
rect 17378 6748 17388 6804
rect 17444 6748 17948 6804
rect 18004 6748 18014 6804
rect 38322 6748 38332 6804
rect 38388 6748 40796 6804
rect 40852 6748 40862 6804
rect 13010 6636 13020 6692
rect 13076 6636 14476 6692
rect 14532 6636 14542 6692
rect 16594 6636 16604 6692
rect 16660 6636 33628 6692
rect 33684 6636 33694 6692
rect 40674 6636 40684 6692
rect 40740 6636 43484 6692
rect 43540 6636 43550 6692
rect 46274 6636 46284 6692
rect 46340 6636 46844 6692
rect 46900 6636 46910 6692
rect 18722 6524 18732 6580
rect 18788 6524 21644 6580
rect 21700 6524 21710 6580
rect 26674 6524 26684 6580
rect 26740 6524 29596 6580
rect 29652 6524 36204 6580
rect 36260 6524 36270 6580
rect 36754 6524 36764 6580
rect 36820 6524 38108 6580
rect 38164 6524 38556 6580
rect 38612 6524 39788 6580
rect 39844 6524 39854 6580
rect 40114 6524 40124 6580
rect 40180 6524 41356 6580
rect 41412 6524 41422 6580
rect 41682 6524 41692 6580
rect 41748 6524 41916 6580
rect 41972 6524 46396 6580
rect 46452 6524 46462 6580
rect 40124 6468 40180 6524
rect 42476 6468 42532 6524
rect 39666 6412 39676 6468
rect 39732 6412 40180 6468
rect 42466 6412 42476 6468
rect 42532 6412 42542 6468
rect 37650 6300 37660 6356
rect 37716 6300 38892 6356
rect 38948 6300 38958 6356
rect 5766 6244 5776 6300
rect 5832 6244 5880 6300
rect 5936 6244 5984 6300
rect 6040 6244 6088 6300
rect 6144 6244 6192 6300
rect 6248 6244 6296 6300
rect 6352 6244 6362 6300
rect 41766 6244 41776 6300
rect 41832 6244 41880 6300
rect 41936 6244 41984 6300
rect 42040 6244 42088 6300
rect 42144 6244 42192 6300
rect 42248 6244 42296 6300
rect 42352 6244 42362 6300
rect 12674 6076 12684 6132
rect 12740 6076 13804 6132
rect 13860 6076 15932 6132
rect 15988 6076 15998 6132
rect 36194 6076 36204 6132
rect 36260 6076 37548 6132
rect 37604 6076 37614 6132
rect 38882 6076 38892 6132
rect 38948 6076 40348 6132
rect 40404 6076 41244 6132
rect 41300 6076 41916 6132
rect 41972 6076 46284 6132
rect 46340 6076 46350 6132
rect 49520 6020 50960 6104
rect 13346 5964 13356 6020
rect 13412 5964 16380 6020
rect 16436 5964 16446 6020
rect 33058 5964 33068 6020
rect 33124 5964 43484 6020
rect 43540 5964 43550 6020
rect 47730 5964 47740 6020
rect 47796 5964 50960 6020
rect 26450 5852 26460 5908
rect 26516 5852 29036 5908
rect 29092 5852 36652 5908
rect 36708 5852 36718 5908
rect 41346 5852 41356 5908
rect 41412 5852 41692 5908
rect 41748 5852 41758 5908
rect 42802 5852 42812 5908
rect 42868 5852 44604 5908
rect 44660 5852 44670 5908
rect 49520 5880 50960 5964
rect 39890 5628 39900 5684
rect 39956 5628 46396 5684
rect 46452 5628 46462 5684
rect 2046 5460 2056 5516
rect 2112 5460 2160 5516
rect 2216 5460 2264 5516
rect 2320 5460 2368 5516
rect 2424 5460 2472 5516
rect 2528 5460 2576 5516
rect 2632 5460 2642 5516
rect 38046 5460 38056 5516
rect 38112 5460 38160 5516
rect 38216 5460 38264 5516
rect 38320 5460 38368 5516
rect 38424 5460 38472 5516
rect 38528 5460 38576 5516
rect 38632 5460 38642 5516
rect 40674 5404 40684 5460
rect 40740 5404 41692 5460
rect 41748 5404 42700 5460
rect 42756 5404 43596 5460
rect 43652 5404 43662 5460
rect 40450 5292 40460 5348
rect 40516 5292 41468 5348
rect 41524 5292 41534 5348
rect 42242 5292 42252 5348
rect 42308 5292 43708 5348
rect 43764 5292 43774 5348
rect 8978 5180 8988 5236
rect 9044 5180 16940 5236
rect 16996 5180 18172 5236
rect 18228 5180 22876 5236
rect 22932 5180 22942 5236
rect 38322 5180 38332 5236
rect 38388 5180 44380 5236
rect 44436 5180 44446 5236
rect 30370 5068 30380 5124
rect 30436 5068 33068 5124
rect 33124 5068 33134 5124
rect 41346 5068 41356 5124
rect 41412 5068 44268 5124
rect 44324 5068 44334 5124
rect 26002 4956 26012 5012
rect 26068 4956 28028 5012
rect 28084 4956 29260 5012
rect 29316 4956 29484 5012
rect 29540 4956 29708 5012
rect 29764 4956 29932 5012
rect 29988 4956 33516 5012
rect 33572 4956 33852 5012
rect 33908 4956 33918 5012
rect 34850 4956 34860 5012
rect 34916 4956 37324 5012
rect 37380 4956 37548 5012
rect 37604 4956 38108 5012
rect 38164 4956 38892 5012
rect 38948 4956 38958 5012
rect 40226 4956 40236 5012
rect 40292 4956 43260 5012
rect 43316 4956 43326 5012
rect 34626 4844 34636 4900
rect 34692 4844 42924 4900
rect 42980 4844 42990 4900
rect 32498 4732 32508 4788
rect 32564 4732 39340 4788
rect 39396 4732 39406 4788
rect 42466 4732 42476 4788
rect 42532 4732 46396 4788
rect 46452 4732 46462 4788
rect 5766 4676 5776 4732
rect 5832 4676 5880 4732
rect 5936 4676 5984 4732
rect 6040 4676 6088 4732
rect 6144 4676 6192 4732
rect 6248 4676 6296 4732
rect 6352 4676 6362 4732
rect 41766 4676 41776 4732
rect 41832 4676 41880 4732
rect 41936 4676 41984 4732
rect 42040 4676 42088 4732
rect 42144 4676 42192 4732
rect 42248 4676 42296 4732
rect 42352 4676 42362 4732
rect 22530 4620 22540 4676
rect 22596 4620 24220 4676
rect 24276 4620 34412 4676
rect 34468 4620 34478 4676
rect 47842 4620 47852 4676
rect 47908 4620 48692 4676
rect 48636 4564 48692 4620
rect 49520 4564 50960 4648
rect 26450 4508 26460 4564
rect 26516 4508 29708 4564
rect 29764 4508 34188 4564
rect 34244 4508 34254 4564
rect 38434 4508 38444 4564
rect 38500 4508 47180 4564
rect 47236 4508 47740 4564
rect 47796 4508 47806 4564
rect 48636 4508 50960 4564
rect 20402 4396 20412 4452
rect 20468 4396 35756 4452
rect 35812 4396 35822 4452
rect 39330 4396 39340 4452
rect 39396 4396 40124 4452
rect 40180 4396 40796 4452
rect 40852 4396 42476 4452
rect 42532 4396 42542 4452
rect 49520 4424 50960 4508
rect 23314 4284 23324 4340
rect 23380 4284 23772 4340
rect 23828 4284 25676 4340
rect 25732 4284 25742 4340
rect 34066 4284 34076 4340
rect 34132 4284 34636 4340
rect 34692 4284 34702 4340
rect 2046 3892 2056 3948
rect 2112 3892 2160 3948
rect 2216 3892 2264 3948
rect 2320 3892 2368 3948
rect 2424 3892 2472 3948
rect 2528 3892 2576 3948
rect 2632 3892 2642 3948
rect 38046 3892 38056 3948
rect 38112 3892 38160 3948
rect 38216 3892 38264 3948
rect 38320 3892 38368 3948
rect 38424 3892 38472 3948
rect 38528 3892 38576 3948
rect 38632 3892 38642 3948
rect 29250 3612 29260 3668
rect 29316 3612 30156 3668
rect 30212 3612 30222 3668
rect 35410 3612 35420 3668
rect 35476 3612 37884 3668
rect 37940 3612 43148 3668
rect 43204 3612 43214 3668
rect 392 3528 1820 3556
rect -960 3500 1820 3528
rect 1876 3500 1886 3556
rect -960 3304 480 3500
rect 26338 3388 26348 3444
rect 26404 3388 29708 3444
rect 29764 3388 37100 3444
rect 37156 3388 37166 3444
rect 5766 3108 5776 3164
rect 5832 3108 5880 3164
rect 5936 3108 5984 3164
rect 6040 3108 6088 3164
rect 6144 3108 6192 3164
rect 6248 3108 6296 3164
rect 6352 3108 6362 3164
rect 41766 3108 41776 3164
rect 41832 3108 41880 3164
rect 41936 3108 41984 3164
rect 42040 3108 42088 3164
rect 42144 3108 42192 3164
rect 42248 3108 42296 3164
rect 42352 3108 42362 3164
rect 49520 3108 50960 3192
rect 47730 3052 47740 3108
rect 47796 3052 50960 3108
rect 49520 2968 50960 3052
rect 49520 1652 50960 1736
rect 48066 1596 48076 1652
rect 48132 1596 50960 1652
rect 49520 1512 50960 1596
<< via3 >>
rect 2056 46228 2112 46284
rect 2160 46228 2216 46284
rect 2264 46228 2320 46284
rect 2368 46228 2424 46284
rect 2472 46228 2528 46284
rect 2576 46228 2632 46284
rect 38056 46228 38112 46284
rect 38160 46228 38216 46284
rect 38264 46228 38320 46284
rect 38368 46228 38424 46284
rect 38472 46228 38528 46284
rect 38576 46228 38632 46284
rect 5776 45444 5832 45500
rect 5880 45444 5936 45500
rect 5984 45444 6040 45500
rect 6088 45444 6144 45500
rect 6192 45444 6248 45500
rect 6296 45444 6352 45500
rect 41776 45444 41832 45500
rect 41880 45444 41936 45500
rect 41984 45444 42040 45500
rect 42088 45444 42144 45500
rect 42192 45444 42248 45500
rect 42296 45444 42352 45500
rect 2056 44660 2112 44716
rect 2160 44660 2216 44716
rect 2264 44660 2320 44716
rect 2368 44660 2424 44716
rect 2472 44660 2528 44716
rect 2576 44660 2632 44716
rect 38056 44660 38112 44716
rect 38160 44660 38216 44716
rect 38264 44660 38320 44716
rect 38368 44660 38424 44716
rect 38472 44660 38528 44716
rect 38576 44660 38632 44716
rect 5776 43876 5832 43932
rect 5880 43876 5936 43932
rect 5984 43876 6040 43932
rect 6088 43876 6144 43932
rect 6192 43876 6248 43932
rect 6296 43876 6352 43932
rect 41776 43876 41832 43932
rect 41880 43876 41936 43932
rect 41984 43876 42040 43932
rect 42088 43876 42144 43932
rect 42192 43876 42248 43932
rect 42296 43876 42352 43932
rect 2056 43092 2112 43148
rect 2160 43092 2216 43148
rect 2264 43092 2320 43148
rect 2368 43092 2424 43148
rect 2472 43092 2528 43148
rect 2576 43092 2632 43148
rect 38056 43092 38112 43148
rect 38160 43092 38216 43148
rect 38264 43092 38320 43148
rect 38368 43092 38424 43148
rect 38472 43092 38528 43148
rect 38576 43092 38632 43148
rect 5776 42308 5832 42364
rect 5880 42308 5936 42364
rect 5984 42308 6040 42364
rect 6088 42308 6144 42364
rect 6192 42308 6248 42364
rect 6296 42308 6352 42364
rect 41776 42308 41832 42364
rect 41880 42308 41936 42364
rect 41984 42308 42040 42364
rect 42088 42308 42144 42364
rect 42192 42308 42248 42364
rect 42296 42308 42352 42364
rect 2056 41524 2112 41580
rect 2160 41524 2216 41580
rect 2264 41524 2320 41580
rect 2368 41524 2424 41580
rect 2472 41524 2528 41580
rect 2576 41524 2632 41580
rect 38056 41524 38112 41580
rect 38160 41524 38216 41580
rect 38264 41524 38320 41580
rect 38368 41524 38424 41580
rect 38472 41524 38528 41580
rect 38576 41524 38632 41580
rect 5776 40740 5832 40796
rect 5880 40740 5936 40796
rect 5984 40740 6040 40796
rect 6088 40740 6144 40796
rect 6192 40740 6248 40796
rect 6296 40740 6352 40796
rect 41776 40740 41832 40796
rect 41880 40740 41936 40796
rect 41984 40740 42040 40796
rect 42088 40740 42144 40796
rect 42192 40740 42248 40796
rect 42296 40740 42352 40796
rect 2056 39956 2112 40012
rect 2160 39956 2216 40012
rect 2264 39956 2320 40012
rect 2368 39956 2424 40012
rect 2472 39956 2528 40012
rect 2576 39956 2632 40012
rect 38056 39956 38112 40012
rect 38160 39956 38216 40012
rect 38264 39956 38320 40012
rect 38368 39956 38424 40012
rect 38472 39956 38528 40012
rect 38576 39956 38632 40012
rect 5776 39172 5832 39228
rect 5880 39172 5936 39228
rect 5984 39172 6040 39228
rect 6088 39172 6144 39228
rect 6192 39172 6248 39228
rect 6296 39172 6352 39228
rect 41776 39172 41832 39228
rect 41880 39172 41936 39228
rect 41984 39172 42040 39228
rect 42088 39172 42144 39228
rect 42192 39172 42248 39228
rect 42296 39172 42352 39228
rect 2056 38388 2112 38444
rect 2160 38388 2216 38444
rect 2264 38388 2320 38444
rect 2368 38388 2424 38444
rect 2472 38388 2528 38444
rect 2576 38388 2632 38444
rect 38056 38388 38112 38444
rect 38160 38388 38216 38444
rect 38264 38388 38320 38444
rect 38368 38388 38424 38444
rect 38472 38388 38528 38444
rect 38576 38388 38632 38444
rect 5776 37604 5832 37660
rect 5880 37604 5936 37660
rect 5984 37604 6040 37660
rect 6088 37604 6144 37660
rect 6192 37604 6248 37660
rect 6296 37604 6352 37660
rect 41776 37604 41832 37660
rect 41880 37604 41936 37660
rect 41984 37604 42040 37660
rect 42088 37604 42144 37660
rect 42192 37604 42248 37660
rect 42296 37604 42352 37660
rect 2056 36820 2112 36876
rect 2160 36820 2216 36876
rect 2264 36820 2320 36876
rect 2368 36820 2424 36876
rect 2472 36820 2528 36876
rect 2576 36820 2632 36876
rect 38056 36820 38112 36876
rect 38160 36820 38216 36876
rect 38264 36820 38320 36876
rect 38368 36820 38424 36876
rect 38472 36820 38528 36876
rect 38576 36820 38632 36876
rect 5776 36036 5832 36092
rect 5880 36036 5936 36092
rect 5984 36036 6040 36092
rect 6088 36036 6144 36092
rect 6192 36036 6248 36092
rect 6296 36036 6352 36092
rect 41776 36036 41832 36092
rect 41880 36036 41936 36092
rect 41984 36036 42040 36092
rect 42088 36036 42144 36092
rect 42192 36036 42248 36092
rect 42296 36036 42352 36092
rect 2056 35252 2112 35308
rect 2160 35252 2216 35308
rect 2264 35252 2320 35308
rect 2368 35252 2424 35308
rect 2472 35252 2528 35308
rect 2576 35252 2632 35308
rect 38056 35252 38112 35308
rect 38160 35252 38216 35308
rect 38264 35252 38320 35308
rect 38368 35252 38424 35308
rect 38472 35252 38528 35308
rect 38576 35252 38632 35308
rect 5776 34468 5832 34524
rect 5880 34468 5936 34524
rect 5984 34468 6040 34524
rect 6088 34468 6144 34524
rect 6192 34468 6248 34524
rect 6296 34468 6352 34524
rect 41776 34468 41832 34524
rect 41880 34468 41936 34524
rect 41984 34468 42040 34524
rect 42088 34468 42144 34524
rect 42192 34468 42248 34524
rect 42296 34468 42352 34524
rect 2056 33684 2112 33740
rect 2160 33684 2216 33740
rect 2264 33684 2320 33740
rect 2368 33684 2424 33740
rect 2472 33684 2528 33740
rect 2576 33684 2632 33740
rect 38056 33684 38112 33740
rect 38160 33684 38216 33740
rect 38264 33684 38320 33740
rect 38368 33684 38424 33740
rect 38472 33684 38528 33740
rect 38576 33684 38632 33740
rect 5776 32900 5832 32956
rect 5880 32900 5936 32956
rect 5984 32900 6040 32956
rect 6088 32900 6144 32956
rect 6192 32900 6248 32956
rect 6296 32900 6352 32956
rect 41776 32900 41832 32956
rect 41880 32900 41936 32956
rect 41984 32900 42040 32956
rect 42088 32900 42144 32956
rect 42192 32900 42248 32956
rect 42296 32900 42352 32956
rect 2056 32116 2112 32172
rect 2160 32116 2216 32172
rect 2264 32116 2320 32172
rect 2368 32116 2424 32172
rect 2472 32116 2528 32172
rect 2576 32116 2632 32172
rect 38056 32116 38112 32172
rect 38160 32116 38216 32172
rect 38264 32116 38320 32172
rect 38368 32116 38424 32172
rect 38472 32116 38528 32172
rect 38576 32116 38632 32172
rect 5776 31332 5832 31388
rect 5880 31332 5936 31388
rect 5984 31332 6040 31388
rect 6088 31332 6144 31388
rect 6192 31332 6248 31388
rect 6296 31332 6352 31388
rect 41776 31332 41832 31388
rect 41880 31332 41936 31388
rect 41984 31332 42040 31388
rect 42088 31332 42144 31388
rect 42192 31332 42248 31388
rect 42296 31332 42352 31388
rect 2056 30548 2112 30604
rect 2160 30548 2216 30604
rect 2264 30548 2320 30604
rect 2368 30548 2424 30604
rect 2472 30548 2528 30604
rect 2576 30548 2632 30604
rect 38056 30548 38112 30604
rect 38160 30548 38216 30604
rect 38264 30548 38320 30604
rect 38368 30548 38424 30604
rect 38472 30548 38528 30604
rect 38576 30548 38632 30604
rect 5776 29764 5832 29820
rect 5880 29764 5936 29820
rect 5984 29764 6040 29820
rect 6088 29764 6144 29820
rect 6192 29764 6248 29820
rect 6296 29764 6352 29820
rect 41776 29764 41832 29820
rect 41880 29764 41936 29820
rect 41984 29764 42040 29820
rect 42088 29764 42144 29820
rect 42192 29764 42248 29820
rect 42296 29764 42352 29820
rect 2056 28980 2112 29036
rect 2160 28980 2216 29036
rect 2264 28980 2320 29036
rect 2368 28980 2424 29036
rect 2472 28980 2528 29036
rect 2576 28980 2632 29036
rect 38056 28980 38112 29036
rect 38160 28980 38216 29036
rect 38264 28980 38320 29036
rect 38368 28980 38424 29036
rect 38472 28980 38528 29036
rect 38576 28980 38632 29036
rect 5776 28196 5832 28252
rect 5880 28196 5936 28252
rect 5984 28196 6040 28252
rect 6088 28196 6144 28252
rect 6192 28196 6248 28252
rect 6296 28196 6352 28252
rect 41776 28196 41832 28252
rect 41880 28196 41936 28252
rect 41984 28196 42040 28252
rect 42088 28196 42144 28252
rect 42192 28196 42248 28252
rect 42296 28196 42352 28252
rect 2056 27412 2112 27468
rect 2160 27412 2216 27468
rect 2264 27412 2320 27468
rect 2368 27412 2424 27468
rect 2472 27412 2528 27468
rect 2576 27412 2632 27468
rect 38056 27412 38112 27468
rect 38160 27412 38216 27468
rect 38264 27412 38320 27468
rect 38368 27412 38424 27468
rect 38472 27412 38528 27468
rect 38576 27412 38632 27468
rect 5776 26628 5832 26684
rect 5880 26628 5936 26684
rect 5984 26628 6040 26684
rect 6088 26628 6144 26684
rect 6192 26628 6248 26684
rect 6296 26628 6352 26684
rect 41776 26628 41832 26684
rect 41880 26628 41936 26684
rect 41984 26628 42040 26684
rect 42088 26628 42144 26684
rect 42192 26628 42248 26684
rect 42296 26628 42352 26684
rect 2056 25844 2112 25900
rect 2160 25844 2216 25900
rect 2264 25844 2320 25900
rect 2368 25844 2424 25900
rect 2472 25844 2528 25900
rect 2576 25844 2632 25900
rect 38056 25844 38112 25900
rect 38160 25844 38216 25900
rect 38264 25844 38320 25900
rect 38368 25844 38424 25900
rect 38472 25844 38528 25900
rect 38576 25844 38632 25900
rect 5776 25060 5832 25116
rect 5880 25060 5936 25116
rect 5984 25060 6040 25116
rect 6088 25060 6144 25116
rect 6192 25060 6248 25116
rect 6296 25060 6352 25116
rect 41776 25060 41832 25116
rect 41880 25060 41936 25116
rect 41984 25060 42040 25116
rect 42088 25060 42144 25116
rect 42192 25060 42248 25116
rect 42296 25060 42352 25116
rect 2056 24276 2112 24332
rect 2160 24276 2216 24332
rect 2264 24276 2320 24332
rect 2368 24276 2424 24332
rect 2472 24276 2528 24332
rect 2576 24276 2632 24332
rect 38056 24276 38112 24332
rect 38160 24276 38216 24332
rect 38264 24276 38320 24332
rect 38368 24276 38424 24332
rect 38472 24276 38528 24332
rect 38576 24276 38632 24332
rect 5776 23492 5832 23548
rect 5880 23492 5936 23548
rect 5984 23492 6040 23548
rect 6088 23492 6144 23548
rect 6192 23492 6248 23548
rect 6296 23492 6352 23548
rect 41776 23492 41832 23548
rect 41880 23492 41936 23548
rect 41984 23492 42040 23548
rect 42088 23492 42144 23548
rect 42192 23492 42248 23548
rect 42296 23492 42352 23548
rect 2056 22708 2112 22764
rect 2160 22708 2216 22764
rect 2264 22708 2320 22764
rect 2368 22708 2424 22764
rect 2472 22708 2528 22764
rect 2576 22708 2632 22764
rect 38056 22708 38112 22764
rect 38160 22708 38216 22764
rect 38264 22708 38320 22764
rect 38368 22708 38424 22764
rect 38472 22708 38528 22764
rect 38576 22708 38632 22764
rect 5776 21924 5832 21980
rect 5880 21924 5936 21980
rect 5984 21924 6040 21980
rect 6088 21924 6144 21980
rect 6192 21924 6248 21980
rect 6296 21924 6352 21980
rect 41776 21924 41832 21980
rect 41880 21924 41936 21980
rect 41984 21924 42040 21980
rect 42088 21924 42144 21980
rect 42192 21924 42248 21980
rect 42296 21924 42352 21980
rect 2056 21140 2112 21196
rect 2160 21140 2216 21196
rect 2264 21140 2320 21196
rect 2368 21140 2424 21196
rect 2472 21140 2528 21196
rect 2576 21140 2632 21196
rect 38056 21140 38112 21196
rect 38160 21140 38216 21196
rect 38264 21140 38320 21196
rect 38368 21140 38424 21196
rect 38472 21140 38528 21196
rect 38576 21140 38632 21196
rect 5776 20356 5832 20412
rect 5880 20356 5936 20412
rect 5984 20356 6040 20412
rect 6088 20356 6144 20412
rect 6192 20356 6248 20412
rect 6296 20356 6352 20412
rect 41776 20356 41832 20412
rect 41880 20356 41936 20412
rect 41984 20356 42040 20412
rect 42088 20356 42144 20412
rect 42192 20356 42248 20412
rect 42296 20356 42352 20412
rect 2056 19572 2112 19628
rect 2160 19572 2216 19628
rect 2264 19572 2320 19628
rect 2368 19572 2424 19628
rect 2472 19572 2528 19628
rect 2576 19572 2632 19628
rect 38056 19572 38112 19628
rect 38160 19572 38216 19628
rect 38264 19572 38320 19628
rect 38368 19572 38424 19628
rect 38472 19572 38528 19628
rect 38576 19572 38632 19628
rect 5776 18788 5832 18844
rect 5880 18788 5936 18844
rect 5984 18788 6040 18844
rect 6088 18788 6144 18844
rect 6192 18788 6248 18844
rect 6296 18788 6352 18844
rect 41776 18788 41832 18844
rect 41880 18788 41936 18844
rect 41984 18788 42040 18844
rect 42088 18788 42144 18844
rect 42192 18788 42248 18844
rect 42296 18788 42352 18844
rect 2056 18004 2112 18060
rect 2160 18004 2216 18060
rect 2264 18004 2320 18060
rect 2368 18004 2424 18060
rect 2472 18004 2528 18060
rect 2576 18004 2632 18060
rect 38056 18004 38112 18060
rect 38160 18004 38216 18060
rect 38264 18004 38320 18060
rect 38368 18004 38424 18060
rect 38472 18004 38528 18060
rect 38576 18004 38632 18060
rect 5776 17220 5832 17276
rect 5880 17220 5936 17276
rect 5984 17220 6040 17276
rect 6088 17220 6144 17276
rect 6192 17220 6248 17276
rect 6296 17220 6352 17276
rect 41776 17220 41832 17276
rect 41880 17220 41936 17276
rect 41984 17220 42040 17276
rect 42088 17220 42144 17276
rect 42192 17220 42248 17276
rect 42296 17220 42352 17276
rect 2056 16436 2112 16492
rect 2160 16436 2216 16492
rect 2264 16436 2320 16492
rect 2368 16436 2424 16492
rect 2472 16436 2528 16492
rect 2576 16436 2632 16492
rect 38056 16436 38112 16492
rect 38160 16436 38216 16492
rect 38264 16436 38320 16492
rect 38368 16436 38424 16492
rect 38472 16436 38528 16492
rect 38576 16436 38632 16492
rect 31052 16380 31108 16436
rect 5776 15652 5832 15708
rect 5880 15652 5936 15708
rect 5984 15652 6040 15708
rect 6088 15652 6144 15708
rect 6192 15652 6248 15708
rect 6296 15652 6352 15708
rect 41776 15652 41832 15708
rect 41880 15652 41936 15708
rect 41984 15652 42040 15708
rect 42088 15652 42144 15708
rect 42192 15652 42248 15708
rect 42296 15652 42352 15708
rect 31052 15484 31108 15540
rect 2056 14868 2112 14924
rect 2160 14868 2216 14924
rect 2264 14868 2320 14924
rect 2368 14868 2424 14924
rect 2472 14868 2528 14924
rect 2576 14868 2632 14924
rect 38056 14868 38112 14924
rect 38160 14868 38216 14924
rect 38264 14868 38320 14924
rect 38368 14868 38424 14924
rect 38472 14868 38528 14924
rect 38576 14868 38632 14924
rect 5776 14084 5832 14140
rect 5880 14084 5936 14140
rect 5984 14084 6040 14140
rect 6088 14084 6144 14140
rect 6192 14084 6248 14140
rect 6296 14084 6352 14140
rect 41776 14084 41832 14140
rect 41880 14084 41936 14140
rect 41984 14084 42040 14140
rect 42088 14084 42144 14140
rect 42192 14084 42248 14140
rect 42296 14084 42352 14140
rect 2056 13300 2112 13356
rect 2160 13300 2216 13356
rect 2264 13300 2320 13356
rect 2368 13300 2424 13356
rect 2472 13300 2528 13356
rect 2576 13300 2632 13356
rect 38056 13300 38112 13356
rect 38160 13300 38216 13356
rect 38264 13300 38320 13356
rect 38368 13300 38424 13356
rect 38472 13300 38528 13356
rect 38576 13300 38632 13356
rect 5776 12516 5832 12572
rect 5880 12516 5936 12572
rect 5984 12516 6040 12572
rect 6088 12516 6144 12572
rect 6192 12516 6248 12572
rect 6296 12516 6352 12572
rect 41776 12516 41832 12572
rect 41880 12516 41936 12572
rect 41984 12516 42040 12572
rect 42088 12516 42144 12572
rect 42192 12516 42248 12572
rect 42296 12516 42352 12572
rect 2056 11732 2112 11788
rect 2160 11732 2216 11788
rect 2264 11732 2320 11788
rect 2368 11732 2424 11788
rect 2472 11732 2528 11788
rect 2576 11732 2632 11788
rect 38056 11732 38112 11788
rect 38160 11732 38216 11788
rect 38264 11732 38320 11788
rect 38368 11732 38424 11788
rect 38472 11732 38528 11788
rect 38576 11732 38632 11788
rect 5776 10948 5832 11004
rect 5880 10948 5936 11004
rect 5984 10948 6040 11004
rect 6088 10948 6144 11004
rect 6192 10948 6248 11004
rect 6296 10948 6352 11004
rect 41776 10948 41832 11004
rect 41880 10948 41936 11004
rect 41984 10948 42040 11004
rect 42088 10948 42144 11004
rect 42192 10948 42248 11004
rect 42296 10948 42352 11004
rect 2056 10164 2112 10220
rect 2160 10164 2216 10220
rect 2264 10164 2320 10220
rect 2368 10164 2424 10220
rect 2472 10164 2528 10220
rect 2576 10164 2632 10220
rect 38056 10164 38112 10220
rect 38160 10164 38216 10220
rect 38264 10164 38320 10220
rect 38368 10164 38424 10220
rect 38472 10164 38528 10220
rect 38576 10164 38632 10220
rect 5776 9380 5832 9436
rect 5880 9380 5936 9436
rect 5984 9380 6040 9436
rect 6088 9380 6144 9436
rect 6192 9380 6248 9436
rect 6296 9380 6352 9436
rect 41776 9380 41832 9436
rect 41880 9380 41936 9436
rect 41984 9380 42040 9436
rect 42088 9380 42144 9436
rect 42192 9380 42248 9436
rect 42296 9380 42352 9436
rect 2056 8596 2112 8652
rect 2160 8596 2216 8652
rect 2264 8596 2320 8652
rect 2368 8596 2424 8652
rect 2472 8596 2528 8652
rect 2576 8596 2632 8652
rect 38056 8596 38112 8652
rect 38160 8596 38216 8652
rect 38264 8596 38320 8652
rect 38368 8596 38424 8652
rect 38472 8596 38528 8652
rect 38576 8596 38632 8652
rect 5776 7812 5832 7868
rect 5880 7812 5936 7868
rect 5984 7812 6040 7868
rect 6088 7812 6144 7868
rect 6192 7812 6248 7868
rect 6296 7812 6352 7868
rect 41776 7812 41832 7868
rect 41880 7812 41936 7868
rect 41984 7812 42040 7868
rect 42088 7812 42144 7868
rect 42192 7812 42248 7868
rect 42296 7812 42352 7868
rect 2056 7028 2112 7084
rect 2160 7028 2216 7084
rect 2264 7028 2320 7084
rect 2368 7028 2424 7084
rect 2472 7028 2528 7084
rect 2576 7028 2632 7084
rect 38056 7028 38112 7084
rect 38160 7028 38216 7084
rect 38264 7028 38320 7084
rect 38368 7028 38424 7084
rect 38472 7028 38528 7084
rect 38576 7028 38632 7084
rect 5776 6244 5832 6300
rect 5880 6244 5936 6300
rect 5984 6244 6040 6300
rect 6088 6244 6144 6300
rect 6192 6244 6248 6300
rect 6296 6244 6352 6300
rect 41776 6244 41832 6300
rect 41880 6244 41936 6300
rect 41984 6244 42040 6300
rect 42088 6244 42144 6300
rect 42192 6244 42248 6300
rect 42296 6244 42352 6300
rect 2056 5460 2112 5516
rect 2160 5460 2216 5516
rect 2264 5460 2320 5516
rect 2368 5460 2424 5516
rect 2472 5460 2528 5516
rect 2576 5460 2632 5516
rect 38056 5460 38112 5516
rect 38160 5460 38216 5516
rect 38264 5460 38320 5516
rect 38368 5460 38424 5516
rect 38472 5460 38528 5516
rect 38576 5460 38632 5516
rect 5776 4676 5832 4732
rect 5880 4676 5936 4732
rect 5984 4676 6040 4732
rect 6088 4676 6144 4732
rect 6192 4676 6248 4732
rect 6296 4676 6352 4732
rect 41776 4676 41832 4732
rect 41880 4676 41936 4732
rect 41984 4676 42040 4732
rect 42088 4676 42144 4732
rect 42192 4676 42248 4732
rect 42296 4676 42352 4732
rect 2056 3892 2112 3948
rect 2160 3892 2216 3948
rect 2264 3892 2320 3948
rect 2368 3892 2424 3948
rect 2472 3892 2528 3948
rect 2576 3892 2632 3948
rect 38056 3892 38112 3948
rect 38160 3892 38216 3948
rect 38264 3892 38320 3948
rect 38368 3892 38424 3948
rect 38472 3892 38528 3948
rect 38576 3892 38632 3948
rect 5776 3108 5832 3164
rect 5880 3108 5936 3164
rect 5984 3108 6040 3164
rect 6088 3108 6144 3164
rect 6192 3108 6248 3164
rect 6296 3108 6352 3164
rect 41776 3108 41832 3164
rect 41880 3108 41936 3164
rect 41984 3108 42040 3164
rect 42088 3108 42144 3164
rect 42192 3108 42248 3164
rect 42296 3108 42352 3164
<< metal4 >>
rect 2034 46284 2654 46316
rect 2034 46228 2056 46284
rect 2112 46228 2160 46284
rect 2216 46228 2264 46284
rect 2320 46228 2368 46284
rect 2424 46228 2472 46284
rect 2528 46228 2576 46284
rect 2632 46228 2654 46284
rect 2034 44716 2654 46228
rect 2034 44660 2056 44716
rect 2112 44660 2160 44716
rect 2216 44660 2264 44716
rect 2320 44660 2368 44716
rect 2424 44660 2472 44716
rect 2528 44660 2576 44716
rect 2632 44660 2654 44716
rect 2034 43148 2654 44660
rect 2034 43092 2056 43148
rect 2112 43092 2160 43148
rect 2216 43092 2264 43148
rect 2320 43092 2368 43148
rect 2424 43092 2472 43148
rect 2528 43092 2576 43148
rect 2632 43092 2654 43148
rect 2034 41580 2654 43092
rect 2034 41524 2056 41580
rect 2112 41524 2160 41580
rect 2216 41524 2264 41580
rect 2320 41524 2368 41580
rect 2424 41524 2472 41580
rect 2528 41524 2576 41580
rect 2632 41524 2654 41580
rect 2034 40012 2654 41524
rect 2034 39956 2056 40012
rect 2112 39956 2160 40012
rect 2216 39956 2264 40012
rect 2320 39956 2368 40012
rect 2424 39956 2472 40012
rect 2528 39956 2576 40012
rect 2632 39956 2654 40012
rect 2034 38444 2654 39956
rect 2034 38388 2056 38444
rect 2112 38388 2160 38444
rect 2216 38388 2264 38444
rect 2320 38388 2368 38444
rect 2424 38388 2472 38444
rect 2528 38388 2576 38444
rect 2632 38388 2654 38444
rect 2034 36876 2654 38388
rect 2034 36820 2056 36876
rect 2112 36820 2160 36876
rect 2216 36820 2264 36876
rect 2320 36820 2368 36876
rect 2424 36820 2472 36876
rect 2528 36820 2576 36876
rect 2632 36820 2654 36876
rect 2034 35308 2654 36820
rect 2034 35252 2056 35308
rect 2112 35252 2160 35308
rect 2216 35252 2264 35308
rect 2320 35252 2368 35308
rect 2424 35252 2472 35308
rect 2528 35252 2576 35308
rect 2632 35252 2654 35308
rect 2034 33740 2654 35252
rect 2034 33684 2056 33740
rect 2112 33684 2160 33740
rect 2216 33684 2264 33740
rect 2320 33684 2368 33740
rect 2424 33684 2472 33740
rect 2528 33684 2576 33740
rect 2632 33684 2654 33740
rect 2034 32172 2654 33684
rect 2034 32116 2056 32172
rect 2112 32116 2160 32172
rect 2216 32116 2264 32172
rect 2320 32116 2368 32172
rect 2424 32116 2472 32172
rect 2528 32116 2576 32172
rect 2632 32116 2654 32172
rect 2034 30604 2654 32116
rect 2034 30548 2056 30604
rect 2112 30548 2160 30604
rect 2216 30548 2264 30604
rect 2320 30548 2368 30604
rect 2424 30548 2472 30604
rect 2528 30548 2576 30604
rect 2632 30548 2654 30604
rect 2034 29036 2654 30548
rect 2034 28980 2056 29036
rect 2112 28980 2160 29036
rect 2216 28980 2264 29036
rect 2320 28980 2368 29036
rect 2424 28980 2472 29036
rect 2528 28980 2576 29036
rect 2632 28980 2654 29036
rect 2034 27468 2654 28980
rect 2034 27412 2056 27468
rect 2112 27412 2160 27468
rect 2216 27412 2264 27468
rect 2320 27412 2368 27468
rect 2424 27412 2472 27468
rect 2528 27412 2576 27468
rect 2632 27412 2654 27468
rect 2034 25900 2654 27412
rect 2034 25844 2056 25900
rect 2112 25844 2160 25900
rect 2216 25844 2264 25900
rect 2320 25844 2368 25900
rect 2424 25844 2472 25900
rect 2528 25844 2576 25900
rect 2632 25844 2654 25900
rect 2034 24332 2654 25844
rect 2034 24276 2056 24332
rect 2112 24276 2160 24332
rect 2216 24276 2264 24332
rect 2320 24276 2368 24332
rect 2424 24276 2472 24332
rect 2528 24276 2576 24332
rect 2632 24276 2654 24332
rect 2034 22764 2654 24276
rect 2034 22708 2056 22764
rect 2112 22708 2160 22764
rect 2216 22708 2264 22764
rect 2320 22708 2368 22764
rect 2424 22708 2472 22764
rect 2528 22708 2576 22764
rect 2632 22708 2654 22764
rect 2034 21196 2654 22708
rect 2034 21140 2056 21196
rect 2112 21140 2160 21196
rect 2216 21140 2264 21196
rect 2320 21140 2368 21196
rect 2424 21140 2472 21196
rect 2528 21140 2576 21196
rect 2632 21140 2654 21196
rect 2034 19628 2654 21140
rect 2034 19572 2056 19628
rect 2112 19572 2160 19628
rect 2216 19572 2264 19628
rect 2320 19572 2368 19628
rect 2424 19572 2472 19628
rect 2528 19572 2576 19628
rect 2632 19572 2654 19628
rect 2034 18060 2654 19572
rect 2034 18004 2056 18060
rect 2112 18004 2160 18060
rect 2216 18004 2264 18060
rect 2320 18004 2368 18060
rect 2424 18004 2472 18060
rect 2528 18004 2576 18060
rect 2632 18004 2654 18060
rect 2034 16492 2654 18004
rect 2034 16436 2056 16492
rect 2112 16436 2160 16492
rect 2216 16436 2264 16492
rect 2320 16436 2368 16492
rect 2424 16436 2472 16492
rect 2528 16436 2576 16492
rect 2632 16436 2654 16492
rect 2034 14924 2654 16436
rect 2034 14868 2056 14924
rect 2112 14868 2160 14924
rect 2216 14868 2264 14924
rect 2320 14868 2368 14924
rect 2424 14868 2472 14924
rect 2528 14868 2576 14924
rect 2632 14868 2654 14924
rect 2034 13356 2654 14868
rect 2034 13300 2056 13356
rect 2112 13300 2160 13356
rect 2216 13300 2264 13356
rect 2320 13300 2368 13356
rect 2424 13300 2472 13356
rect 2528 13300 2576 13356
rect 2632 13300 2654 13356
rect 2034 11788 2654 13300
rect 2034 11732 2056 11788
rect 2112 11732 2160 11788
rect 2216 11732 2264 11788
rect 2320 11732 2368 11788
rect 2424 11732 2472 11788
rect 2528 11732 2576 11788
rect 2632 11732 2654 11788
rect 2034 10220 2654 11732
rect 2034 10164 2056 10220
rect 2112 10164 2160 10220
rect 2216 10164 2264 10220
rect 2320 10164 2368 10220
rect 2424 10164 2472 10220
rect 2528 10164 2576 10220
rect 2632 10164 2654 10220
rect 2034 8652 2654 10164
rect 2034 8596 2056 8652
rect 2112 8596 2160 8652
rect 2216 8596 2264 8652
rect 2320 8596 2368 8652
rect 2424 8596 2472 8652
rect 2528 8596 2576 8652
rect 2632 8596 2654 8652
rect 2034 7084 2654 8596
rect 2034 7028 2056 7084
rect 2112 7028 2160 7084
rect 2216 7028 2264 7084
rect 2320 7028 2368 7084
rect 2424 7028 2472 7084
rect 2528 7028 2576 7084
rect 2632 7028 2654 7084
rect 2034 5516 2654 7028
rect 2034 5460 2056 5516
rect 2112 5460 2160 5516
rect 2216 5460 2264 5516
rect 2320 5460 2368 5516
rect 2424 5460 2472 5516
rect 2528 5460 2576 5516
rect 2632 5460 2654 5516
rect 2034 3948 2654 5460
rect 2034 3892 2056 3948
rect 2112 3892 2160 3948
rect 2216 3892 2264 3948
rect 2320 3892 2368 3948
rect 2424 3892 2472 3948
rect 2528 3892 2576 3948
rect 2632 3892 2654 3948
rect 2034 3076 2654 3892
rect 5754 45500 6374 46316
rect 5754 45444 5776 45500
rect 5832 45444 5880 45500
rect 5936 45444 5984 45500
rect 6040 45444 6088 45500
rect 6144 45444 6192 45500
rect 6248 45444 6296 45500
rect 6352 45444 6374 45500
rect 5754 43932 6374 45444
rect 5754 43876 5776 43932
rect 5832 43876 5880 43932
rect 5936 43876 5984 43932
rect 6040 43876 6088 43932
rect 6144 43876 6192 43932
rect 6248 43876 6296 43932
rect 6352 43876 6374 43932
rect 5754 42364 6374 43876
rect 5754 42308 5776 42364
rect 5832 42308 5880 42364
rect 5936 42308 5984 42364
rect 6040 42308 6088 42364
rect 6144 42308 6192 42364
rect 6248 42308 6296 42364
rect 6352 42308 6374 42364
rect 5754 40796 6374 42308
rect 5754 40740 5776 40796
rect 5832 40740 5880 40796
rect 5936 40740 5984 40796
rect 6040 40740 6088 40796
rect 6144 40740 6192 40796
rect 6248 40740 6296 40796
rect 6352 40740 6374 40796
rect 5754 39228 6374 40740
rect 5754 39172 5776 39228
rect 5832 39172 5880 39228
rect 5936 39172 5984 39228
rect 6040 39172 6088 39228
rect 6144 39172 6192 39228
rect 6248 39172 6296 39228
rect 6352 39172 6374 39228
rect 5754 37660 6374 39172
rect 5754 37604 5776 37660
rect 5832 37604 5880 37660
rect 5936 37604 5984 37660
rect 6040 37604 6088 37660
rect 6144 37604 6192 37660
rect 6248 37604 6296 37660
rect 6352 37604 6374 37660
rect 5754 36092 6374 37604
rect 5754 36036 5776 36092
rect 5832 36036 5880 36092
rect 5936 36036 5984 36092
rect 6040 36036 6088 36092
rect 6144 36036 6192 36092
rect 6248 36036 6296 36092
rect 6352 36036 6374 36092
rect 5754 34524 6374 36036
rect 5754 34468 5776 34524
rect 5832 34468 5880 34524
rect 5936 34468 5984 34524
rect 6040 34468 6088 34524
rect 6144 34468 6192 34524
rect 6248 34468 6296 34524
rect 6352 34468 6374 34524
rect 5754 32956 6374 34468
rect 5754 32900 5776 32956
rect 5832 32900 5880 32956
rect 5936 32900 5984 32956
rect 6040 32900 6088 32956
rect 6144 32900 6192 32956
rect 6248 32900 6296 32956
rect 6352 32900 6374 32956
rect 5754 31388 6374 32900
rect 5754 31332 5776 31388
rect 5832 31332 5880 31388
rect 5936 31332 5984 31388
rect 6040 31332 6088 31388
rect 6144 31332 6192 31388
rect 6248 31332 6296 31388
rect 6352 31332 6374 31388
rect 5754 29820 6374 31332
rect 5754 29764 5776 29820
rect 5832 29764 5880 29820
rect 5936 29764 5984 29820
rect 6040 29764 6088 29820
rect 6144 29764 6192 29820
rect 6248 29764 6296 29820
rect 6352 29764 6374 29820
rect 5754 28252 6374 29764
rect 5754 28196 5776 28252
rect 5832 28196 5880 28252
rect 5936 28196 5984 28252
rect 6040 28196 6088 28252
rect 6144 28196 6192 28252
rect 6248 28196 6296 28252
rect 6352 28196 6374 28252
rect 5754 26684 6374 28196
rect 5754 26628 5776 26684
rect 5832 26628 5880 26684
rect 5936 26628 5984 26684
rect 6040 26628 6088 26684
rect 6144 26628 6192 26684
rect 6248 26628 6296 26684
rect 6352 26628 6374 26684
rect 5754 25116 6374 26628
rect 5754 25060 5776 25116
rect 5832 25060 5880 25116
rect 5936 25060 5984 25116
rect 6040 25060 6088 25116
rect 6144 25060 6192 25116
rect 6248 25060 6296 25116
rect 6352 25060 6374 25116
rect 5754 23548 6374 25060
rect 5754 23492 5776 23548
rect 5832 23492 5880 23548
rect 5936 23492 5984 23548
rect 6040 23492 6088 23548
rect 6144 23492 6192 23548
rect 6248 23492 6296 23548
rect 6352 23492 6374 23548
rect 5754 21980 6374 23492
rect 5754 21924 5776 21980
rect 5832 21924 5880 21980
rect 5936 21924 5984 21980
rect 6040 21924 6088 21980
rect 6144 21924 6192 21980
rect 6248 21924 6296 21980
rect 6352 21924 6374 21980
rect 5754 20412 6374 21924
rect 5754 20356 5776 20412
rect 5832 20356 5880 20412
rect 5936 20356 5984 20412
rect 6040 20356 6088 20412
rect 6144 20356 6192 20412
rect 6248 20356 6296 20412
rect 6352 20356 6374 20412
rect 5754 18844 6374 20356
rect 5754 18788 5776 18844
rect 5832 18788 5880 18844
rect 5936 18788 5984 18844
rect 6040 18788 6088 18844
rect 6144 18788 6192 18844
rect 6248 18788 6296 18844
rect 6352 18788 6374 18844
rect 5754 17276 6374 18788
rect 5754 17220 5776 17276
rect 5832 17220 5880 17276
rect 5936 17220 5984 17276
rect 6040 17220 6088 17276
rect 6144 17220 6192 17276
rect 6248 17220 6296 17276
rect 6352 17220 6374 17276
rect 5754 15708 6374 17220
rect 38034 46284 38654 46316
rect 38034 46228 38056 46284
rect 38112 46228 38160 46284
rect 38216 46228 38264 46284
rect 38320 46228 38368 46284
rect 38424 46228 38472 46284
rect 38528 46228 38576 46284
rect 38632 46228 38654 46284
rect 38034 44716 38654 46228
rect 38034 44660 38056 44716
rect 38112 44660 38160 44716
rect 38216 44660 38264 44716
rect 38320 44660 38368 44716
rect 38424 44660 38472 44716
rect 38528 44660 38576 44716
rect 38632 44660 38654 44716
rect 38034 43148 38654 44660
rect 38034 43092 38056 43148
rect 38112 43092 38160 43148
rect 38216 43092 38264 43148
rect 38320 43092 38368 43148
rect 38424 43092 38472 43148
rect 38528 43092 38576 43148
rect 38632 43092 38654 43148
rect 38034 41580 38654 43092
rect 38034 41524 38056 41580
rect 38112 41524 38160 41580
rect 38216 41524 38264 41580
rect 38320 41524 38368 41580
rect 38424 41524 38472 41580
rect 38528 41524 38576 41580
rect 38632 41524 38654 41580
rect 38034 40012 38654 41524
rect 38034 39956 38056 40012
rect 38112 39956 38160 40012
rect 38216 39956 38264 40012
rect 38320 39956 38368 40012
rect 38424 39956 38472 40012
rect 38528 39956 38576 40012
rect 38632 39956 38654 40012
rect 38034 38444 38654 39956
rect 38034 38388 38056 38444
rect 38112 38388 38160 38444
rect 38216 38388 38264 38444
rect 38320 38388 38368 38444
rect 38424 38388 38472 38444
rect 38528 38388 38576 38444
rect 38632 38388 38654 38444
rect 38034 36876 38654 38388
rect 38034 36820 38056 36876
rect 38112 36820 38160 36876
rect 38216 36820 38264 36876
rect 38320 36820 38368 36876
rect 38424 36820 38472 36876
rect 38528 36820 38576 36876
rect 38632 36820 38654 36876
rect 38034 35308 38654 36820
rect 38034 35252 38056 35308
rect 38112 35252 38160 35308
rect 38216 35252 38264 35308
rect 38320 35252 38368 35308
rect 38424 35252 38472 35308
rect 38528 35252 38576 35308
rect 38632 35252 38654 35308
rect 38034 33740 38654 35252
rect 38034 33684 38056 33740
rect 38112 33684 38160 33740
rect 38216 33684 38264 33740
rect 38320 33684 38368 33740
rect 38424 33684 38472 33740
rect 38528 33684 38576 33740
rect 38632 33684 38654 33740
rect 38034 32172 38654 33684
rect 38034 32116 38056 32172
rect 38112 32116 38160 32172
rect 38216 32116 38264 32172
rect 38320 32116 38368 32172
rect 38424 32116 38472 32172
rect 38528 32116 38576 32172
rect 38632 32116 38654 32172
rect 38034 30604 38654 32116
rect 38034 30548 38056 30604
rect 38112 30548 38160 30604
rect 38216 30548 38264 30604
rect 38320 30548 38368 30604
rect 38424 30548 38472 30604
rect 38528 30548 38576 30604
rect 38632 30548 38654 30604
rect 38034 29036 38654 30548
rect 38034 28980 38056 29036
rect 38112 28980 38160 29036
rect 38216 28980 38264 29036
rect 38320 28980 38368 29036
rect 38424 28980 38472 29036
rect 38528 28980 38576 29036
rect 38632 28980 38654 29036
rect 38034 27468 38654 28980
rect 38034 27412 38056 27468
rect 38112 27412 38160 27468
rect 38216 27412 38264 27468
rect 38320 27412 38368 27468
rect 38424 27412 38472 27468
rect 38528 27412 38576 27468
rect 38632 27412 38654 27468
rect 38034 25900 38654 27412
rect 38034 25844 38056 25900
rect 38112 25844 38160 25900
rect 38216 25844 38264 25900
rect 38320 25844 38368 25900
rect 38424 25844 38472 25900
rect 38528 25844 38576 25900
rect 38632 25844 38654 25900
rect 38034 24332 38654 25844
rect 38034 24276 38056 24332
rect 38112 24276 38160 24332
rect 38216 24276 38264 24332
rect 38320 24276 38368 24332
rect 38424 24276 38472 24332
rect 38528 24276 38576 24332
rect 38632 24276 38654 24332
rect 38034 22764 38654 24276
rect 38034 22708 38056 22764
rect 38112 22708 38160 22764
rect 38216 22708 38264 22764
rect 38320 22708 38368 22764
rect 38424 22708 38472 22764
rect 38528 22708 38576 22764
rect 38632 22708 38654 22764
rect 38034 21196 38654 22708
rect 38034 21140 38056 21196
rect 38112 21140 38160 21196
rect 38216 21140 38264 21196
rect 38320 21140 38368 21196
rect 38424 21140 38472 21196
rect 38528 21140 38576 21196
rect 38632 21140 38654 21196
rect 38034 19628 38654 21140
rect 38034 19572 38056 19628
rect 38112 19572 38160 19628
rect 38216 19572 38264 19628
rect 38320 19572 38368 19628
rect 38424 19572 38472 19628
rect 38528 19572 38576 19628
rect 38632 19572 38654 19628
rect 38034 18060 38654 19572
rect 38034 18004 38056 18060
rect 38112 18004 38160 18060
rect 38216 18004 38264 18060
rect 38320 18004 38368 18060
rect 38424 18004 38472 18060
rect 38528 18004 38576 18060
rect 38632 18004 38654 18060
rect 38034 16492 38654 18004
rect 5754 15652 5776 15708
rect 5832 15652 5880 15708
rect 5936 15652 5984 15708
rect 6040 15652 6088 15708
rect 6144 15652 6192 15708
rect 6248 15652 6296 15708
rect 6352 15652 6374 15708
rect 5754 14140 6374 15652
rect 31052 16436 31108 16446
rect 31052 15540 31108 16380
rect 31052 15474 31108 15484
rect 38034 16436 38056 16492
rect 38112 16436 38160 16492
rect 38216 16436 38264 16492
rect 38320 16436 38368 16492
rect 38424 16436 38472 16492
rect 38528 16436 38576 16492
rect 38632 16436 38654 16492
rect 5754 14084 5776 14140
rect 5832 14084 5880 14140
rect 5936 14084 5984 14140
rect 6040 14084 6088 14140
rect 6144 14084 6192 14140
rect 6248 14084 6296 14140
rect 6352 14084 6374 14140
rect 5754 12572 6374 14084
rect 5754 12516 5776 12572
rect 5832 12516 5880 12572
rect 5936 12516 5984 12572
rect 6040 12516 6088 12572
rect 6144 12516 6192 12572
rect 6248 12516 6296 12572
rect 6352 12516 6374 12572
rect 5754 11004 6374 12516
rect 5754 10948 5776 11004
rect 5832 10948 5880 11004
rect 5936 10948 5984 11004
rect 6040 10948 6088 11004
rect 6144 10948 6192 11004
rect 6248 10948 6296 11004
rect 6352 10948 6374 11004
rect 5754 9436 6374 10948
rect 5754 9380 5776 9436
rect 5832 9380 5880 9436
rect 5936 9380 5984 9436
rect 6040 9380 6088 9436
rect 6144 9380 6192 9436
rect 6248 9380 6296 9436
rect 6352 9380 6374 9436
rect 5754 7868 6374 9380
rect 5754 7812 5776 7868
rect 5832 7812 5880 7868
rect 5936 7812 5984 7868
rect 6040 7812 6088 7868
rect 6144 7812 6192 7868
rect 6248 7812 6296 7868
rect 6352 7812 6374 7868
rect 5754 6300 6374 7812
rect 5754 6244 5776 6300
rect 5832 6244 5880 6300
rect 5936 6244 5984 6300
rect 6040 6244 6088 6300
rect 6144 6244 6192 6300
rect 6248 6244 6296 6300
rect 6352 6244 6374 6300
rect 5754 4732 6374 6244
rect 5754 4676 5776 4732
rect 5832 4676 5880 4732
rect 5936 4676 5984 4732
rect 6040 4676 6088 4732
rect 6144 4676 6192 4732
rect 6248 4676 6296 4732
rect 6352 4676 6374 4732
rect 5754 3164 6374 4676
rect 5754 3108 5776 3164
rect 5832 3108 5880 3164
rect 5936 3108 5984 3164
rect 6040 3108 6088 3164
rect 6144 3108 6192 3164
rect 6248 3108 6296 3164
rect 6352 3108 6374 3164
rect 5754 3076 6374 3108
rect 38034 14924 38654 16436
rect 38034 14868 38056 14924
rect 38112 14868 38160 14924
rect 38216 14868 38264 14924
rect 38320 14868 38368 14924
rect 38424 14868 38472 14924
rect 38528 14868 38576 14924
rect 38632 14868 38654 14924
rect 38034 13356 38654 14868
rect 38034 13300 38056 13356
rect 38112 13300 38160 13356
rect 38216 13300 38264 13356
rect 38320 13300 38368 13356
rect 38424 13300 38472 13356
rect 38528 13300 38576 13356
rect 38632 13300 38654 13356
rect 38034 11788 38654 13300
rect 38034 11732 38056 11788
rect 38112 11732 38160 11788
rect 38216 11732 38264 11788
rect 38320 11732 38368 11788
rect 38424 11732 38472 11788
rect 38528 11732 38576 11788
rect 38632 11732 38654 11788
rect 38034 10220 38654 11732
rect 38034 10164 38056 10220
rect 38112 10164 38160 10220
rect 38216 10164 38264 10220
rect 38320 10164 38368 10220
rect 38424 10164 38472 10220
rect 38528 10164 38576 10220
rect 38632 10164 38654 10220
rect 38034 8652 38654 10164
rect 38034 8596 38056 8652
rect 38112 8596 38160 8652
rect 38216 8596 38264 8652
rect 38320 8596 38368 8652
rect 38424 8596 38472 8652
rect 38528 8596 38576 8652
rect 38632 8596 38654 8652
rect 38034 7084 38654 8596
rect 38034 7028 38056 7084
rect 38112 7028 38160 7084
rect 38216 7028 38264 7084
rect 38320 7028 38368 7084
rect 38424 7028 38472 7084
rect 38528 7028 38576 7084
rect 38632 7028 38654 7084
rect 38034 5516 38654 7028
rect 38034 5460 38056 5516
rect 38112 5460 38160 5516
rect 38216 5460 38264 5516
rect 38320 5460 38368 5516
rect 38424 5460 38472 5516
rect 38528 5460 38576 5516
rect 38632 5460 38654 5516
rect 38034 3948 38654 5460
rect 38034 3892 38056 3948
rect 38112 3892 38160 3948
rect 38216 3892 38264 3948
rect 38320 3892 38368 3948
rect 38424 3892 38472 3948
rect 38528 3892 38576 3948
rect 38632 3892 38654 3948
rect 38034 3076 38654 3892
rect 41754 45500 42374 46316
rect 41754 45444 41776 45500
rect 41832 45444 41880 45500
rect 41936 45444 41984 45500
rect 42040 45444 42088 45500
rect 42144 45444 42192 45500
rect 42248 45444 42296 45500
rect 42352 45444 42374 45500
rect 41754 43932 42374 45444
rect 41754 43876 41776 43932
rect 41832 43876 41880 43932
rect 41936 43876 41984 43932
rect 42040 43876 42088 43932
rect 42144 43876 42192 43932
rect 42248 43876 42296 43932
rect 42352 43876 42374 43932
rect 41754 42364 42374 43876
rect 41754 42308 41776 42364
rect 41832 42308 41880 42364
rect 41936 42308 41984 42364
rect 42040 42308 42088 42364
rect 42144 42308 42192 42364
rect 42248 42308 42296 42364
rect 42352 42308 42374 42364
rect 41754 40796 42374 42308
rect 41754 40740 41776 40796
rect 41832 40740 41880 40796
rect 41936 40740 41984 40796
rect 42040 40740 42088 40796
rect 42144 40740 42192 40796
rect 42248 40740 42296 40796
rect 42352 40740 42374 40796
rect 41754 39228 42374 40740
rect 41754 39172 41776 39228
rect 41832 39172 41880 39228
rect 41936 39172 41984 39228
rect 42040 39172 42088 39228
rect 42144 39172 42192 39228
rect 42248 39172 42296 39228
rect 42352 39172 42374 39228
rect 41754 37660 42374 39172
rect 41754 37604 41776 37660
rect 41832 37604 41880 37660
rect 41936 37604 41984 37660
rect 42040 37604 42088 37660
rect 42144 37604 42192 37660
rect 42248 37604 42296 37660
rect 42352 37604 42374 37660
rect 41754 36092 42374 37604
rect 41754 36036 41776 36092
rect 41832 36036 41880 36092
rect 41936 36036 41984 36092
rect 42040 36036 42088 36092
rect 42144 36036 42192 36092
rect 42248 36036 42296 36092
rect 42352 36036 42374 36092
rect 41754 34524 42374 36036
rect 41754 34468 41776 34524
rect 41832 34468 41880 34524
rect 41936 34468 41984 34524
rect 42040 34468 42088 34524
rect 42144 34468 42192 34524
rect 42248 34468 42296 34524
rect 42352 34468 42374 34524
rect 41754 32956 42374 34468
rect 41754 32900 41776 32956
rect 41832 32900 41880 32956
rect 41936 32900 41984 32956
rect 42040 32900 42088 32956
rect 42144 32900 42192 32956
rect 42248 32900 42296 32956
rect 42352 32900 42374 32956
rect 41754 31388 42374 32900
rect 41754 31332 41776 31388
rect 41832 31332 41880 31388
rect 41936 31332 41984 31388
rect 42040 31332 42088 31388
rect 42144 31332 42192 31388
rect 42248 31332 42296 31388
rect 42352 31332 42374 31388
rect 41754 29820 42374 31332
rect 41754 29764 41776 29820
rect 41832 29764 41880 29820
rect 41936 29764 41984 29820
rect 42040 29764 42088 29820
rect 42144 29764 42192 29820
rect 42248 29764 42296 29820
rect 42352 29764 42374 29820
rect 41754 28252 42374 29764
rect 41754 28196 41776 28252
rect 41832 28196 41880 28252
rect 41936 28196 41984 28252
rect 42040 28196 42088 28252
rect 42144 28196 42192 28252
rect 42248 28196 42296 28252
rect 42352 28196 42374 28252
rect 41754 26684 42374 28196
rect 41754 26628 41776 26684
rect 41832 26628 41880 26684
rect 41936 26628 41984 26684
rect 42040 26628 42088 26684
rect 42144 26628 42192 26684
rect 42248 26628 42296 26684
rect 42352 26628 42374 26684
rect 41754 25116 42374 26628
rect 41754 25060 41776 25116
rect 41832 25060 41880 25116
rect 41936 25060 41984 25116
rect 42040 25060 42088 25116
rect 42144 25060 42192 25116
rect 42248 25060 42296 25116
rect 42352 25060 42374 25116
rect 41754 23548 42374 25060
rect 41754 23492 41776 23548
rect 41832 23492 41880 23548
rect 41936 23492 41984 23548
rect 42040 23492 42088 23548
rect 42144 23492 42192 23548
rect 42248 23492 42296 23548
rect 42352 23492 42374 23548
rect 41754 21980 42374 23492
rect 41754 21924 41776 21980
rect 41832 21924 41880 21980
rect 41936 21924 41984 21980
rect 42040 21924 42088 21980
rect 42144 21924 42192 21980
rect 42248 21924 42296 21980
rect 42352 21924 42374 21980
rect 41754 20412 42374 21924
rect 41754 20356 41776 20412
rect 41832 20356 41880 20412
rect 41936 20356 41984 20412
rect 42040 20356 42088 20412
rect 42144 20356 42192 20412
rect 42248 20356 42296 20412
rect 42352 20356 42374 20412
rect 41754 18844 42374 20356
rect 41754 18788 41776 18844
rect 41832 18788 41880 18844
rect 41936 18788 41984 18844
rect 42040 18788 42088 18844
rect 42144 18788 42192 18844
rect 42248 18788 42296 18844
rect 42352 18788 42374 18844
rect 41754 17276 42374 18788
rect 41754 17220 41776 17276
rect 41832 17220 41880 17276
rect 41936 17220 41984 17276
rect 42040 17220 42088 17276
rect 42144 17220 42192 17276
rect 42248 17220 42296 17276
rect 42352 17220 42374 17276
rect 41754 15708 42374 17220
rect 41754 15652 41776 15708
rect 41832 15652 41880 15708
rect 41936 15652 41984 15708
rect 42040 15652 42088 15708
rect 42144 15652 42192 15708
rect 42248 15652 42296 15708
rect 42352 15652 42374 15708
rect 41754 14140 42374 15652
rect 41754 14084 41776 14140
rect 41832 14084 41880 14140
rect 41936 14084 41984 14140
rect 42040 14084 42088 14140
rect 42144 14084 42192 14140
rect 42248 14084 42296 14140
rect 42352 14084 42374 14140
rect 41754 12572 42374 14084
rect 41754 12516 41776 12572
rect 41832 12516 41880 12572
rect 41936 12516 41984 12572
rect 42040 12516 42088 12572
rect 42144 12516 42192 12572
rect 42248 12516 42296 12572
rect 42352 12516 42374 12572
rect 41754 11004 42374 12516
rect 41754 10948 41776 11004
rect 41832 10948 41880 11004
rect 41936 10948 41984 11004
rect 42040 10948 42088 11004
rect 42144 10948 42192 11004
rect 42248 10948 42296 11004
rect 42352 10948 42374 11004
rect 41754 9436 42374 10948
rect 41754 9380 41776 9436
rect 41832 9380 41880 9436
rect 41936 9380 41984 9436
rect 42040 9380 42088 9436
rect 42144 9380 42192 9436
rect 42248 9380 42296 9436
rect 42352 9380 42374 9436
rect 41754 7868 42374 9380
rect 41754 7812 41776 7868
rect 41832 7812 41880 7868
rect 41936 7812 41984 7868
rect 42040 7812 42088 7868
rect 42144 7812 42192 7868
rect 42248 7812 42296 7868
rect 42352 7812 42374 7868
rect 41754 6300 42374 7812
rect 41754 6244 41776 6300
rect 41832 6244 41880 6300
rect 41936 6244 41984 6300
rect 42040 6244 42088 6300
rect 42144 6244 42192 6300
rect 42248 6244 42296 6300
rect 42352 6244 42374 6300
rect 41754 4732 42374 6244
rect 41754 4676 41776 4732
rect 41832 4676 41880 4732
rect 41936 4676 41984 4732
rect 42040 4676 42088 4732
rect 42144 4676 42192 4732
rect 42248 4676 42296 4732
rect 42352 4676 42374 4732
rect 41754 3164 42374 4676
rect 41754 3108 41776 3164
rect 41832 3108 41880 3164
rect 41936 3108 41984 3164
rect 42040 3108 42088 3164
rect 42144 3108 42192 3164
rect 42248 3108 42296 3164
rect 42352 3108 42374 3164
rect 41754 3076 42374 3108
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__078__A1 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 43344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__078__A2
timestamp 1666464484
transform -1 0 42896 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__079__I
timestamp 1666464484
transform 1 0 38640 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__080__A1
timestamp 1666464484
transform -1 0 33824 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__080__A2
timestamp 1666464484
transform 1 0 34832 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__081__A2
timestamp 1666464484
transform 1 0 39088 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__084__I1
timestamp 1666464484
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__084__S
timestamp 1666464484
transform -1 0 42784 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__086__I0
timestamp 1666464484
transform 1 0 40768 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__086__I1
timestamp 1666464484
transform -1 0 38192 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__086__S
timestamp 1666464484
transform -1 0 40768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__088__I0
timestamp 1666464484
transform -1 0 38640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__088__I1
timestamp 1666464484
transform 1 0 38864 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__088__S
timestamp 1666464484
transform 1 0 41440 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__090__I0
timestamp 1666464484
transform 1 0 41888 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__090__I1
timestamp 1666464484
transform -1 0 41664 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__090__S
timestamp 1666464484
transform 1 0 43680 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__093__I0
timestamp 1666464484
transform 1 0 41888 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__093__I1
timestamp 1666464484
transform 1 0 40768 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__095__I0
timestamp 1666464484
transform 1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__095__I1
timestamp 1666464484
transform 1 0 41104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__097__I0
timestamp 1666464484
transform 1 0 41216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__097__I1
timestamp 1666464484
transform 1 0 40768 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__099__I0
timestamp 1666464484
transform 1 0 43344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__099__I1
timestamp 1666464484
transform -1 0 41216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__102__I0
timestamp 1666464484
transform 1 0 40656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__102__I1
timestamp 1666464484
transform 1 0 38528 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__104__I0
timestamp 1666464484
transform 1 0 41440 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__104__I1
timestamp 1666464484
transform 1 0 36736 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__106__I0
timestamp 1666464484
transform -1 0 36176 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__106__I1
timestamp 1666464484
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__108__I0
timestamp 1666464484
transform 1 0 37408 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__108__I1
timestamp 1666464484
transform 1 0 36400 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__111__I0
timestamp 1666464484
transform 1 0 36176 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__111__I1
timestamp 1666464484
transform 1 0 35616 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__113__I0
timestamp 1666464484
transform 1 0 34048 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__113__I1
timestamp 1666464484
transform 1 0 33264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__115__I0
timestamp 1666464484
transform 1 0 33712 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__115__I1
timestamp 1666464484
transform 1 0 33488 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__117__I0
timestamp 1666464484
transform 1 0 32816 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__117__I1
timestamp 1666464484
transform 1 0 33264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__121__I0
timestamp 1666464484
transform 1 0 34272 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__121__I1
timestamp 1666464484
transform 1 0 34720 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__121__S
timestamp 1666464484
transform -1 0 38080 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__123__I0
timestamp 1666464484
transform 1 0 33936 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__123__I1
timestamp 1666464484
transform 1 0 34832 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__123__S
timestamp 1666464484
transform 1 0 38304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__125__I0
timestamp 1666464484
transform 1 0 38304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__125__I1
timestamp 1666464484
transform 1 0 37408 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__125__S
timestamp 1666464484
transform -1 0 38976 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__127__I0
timestamp 1666464484
transform 1 0 36176 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__127__I1
timestamp 1666464484
transform 1 0 35728 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__127__S
timestamp 1666464484
transform 1 0 38528 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__130__I0
timestamp 1666464484
transform 1 0 38080 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__130__I1
timestamp 1666464484
transform 1 0 36736 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__132__I0
timestamp 1666464484
transform 1 0 35952 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__132__I1
timestamp 1666464484
transform 1 0 36400 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__134__I0
timestamp 1666464484
transform 1 0 36288 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__134__I1
timestamp 1666464484
transform 1 0 36736 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__136__I0
timestamp 1666464484
transform 1 0 36400 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__136__I1
timestamp 1666464484
transform 1 0 36848 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__137__I
timestamp 1666464484
transform 1 0 32032 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__139__I0
timestamp 1666464484
transform 1 0 36848 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__139__I1
timestamp 1666464484
transform 1 0 37296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__140__I
timestamp 1666464484
transform -1 0 32144 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__141__I0
timestamp 1666464484
transform 1 0 39648 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__141__I1
timestamp 1666464484
transform 1 0 36736 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__142__I
timestamp 1666464484
transform 1 0 31808 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__143__I0
timestamp 1666464484
transform 1 0 36960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__143__I1
timestamp 1666464484
transform 1 0 37408 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__144__I
timestamp 1666464484
transform -1 0 30912 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__145__I0
timestamp 1666464484
transform 1 0 37072 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__145__I1
timestamp 1666464484
transform 1 0 37520 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__146__I
timestamp 1666464484
transform -1 0 30128 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__148__I0
timestamp 1666464484
transform 1 0 39648 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__148__I1
timestamp 1666464484
transform 1 0 36736 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__148__S
timestamp 1666464484
transform 1 0 40096 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__149__I
timestamp 1666464484
transform 1 0 30352 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__150__I0
timestamp 1666464484
transform 1 0 36848 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__150__I1
timestamp 1666464484
transform 1 0 37296 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__150__S
timestamp 1666464484
transform 1 0 39648 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__151__I
timestamp 1666464484
transform -1 0 30128 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__152__I0
timestamp 1666464484
transform 1 0 36176 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__152__I1
timestamp 1666464484
transform 1 0 36624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__152__S
timestamp 1666464484
transform 1 0 38752 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__153__I
timestamp 1666464484
transform 1 0 27888 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__154__I0
timestamp 1666464484
transform 1 0 29344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__154__I1
timestamp 1666464484
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__154__S
timestamp 1666464484
transform 1 0 31472 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__156__CLK
timestamp 1666464484
transform 1 0 6832 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__156__D
timestamp 1666464484
transform 1 0 2912 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__157__CLK
timestamp 1666464484
transform 1 0 9632 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__158__CLK
timestamp 1666464484
transform -1 0 16576 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__158__D
timestamp 1666464484
transform -1 0 17024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__159__CLK
timestamp 1666464484
transform 1 0 6720 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__159__D
timestamp 1666464484
transform 1 0 2800 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__160__CLK
timestamp 1666464484
transform -1 0 9072 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__161__CLK
timestamp 1666464484
transform 1 0 12432 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__161__D
timestamp 1666464484
transform -1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__162__CLK
timestamp 1666464484
transform 1 0 5600 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__163__CLK
timestamp 1666464484
transform 1 0 5152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__164__CLK
timestamp 1666464484
transform 1 0 13552 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__164__D
timestamp 1666464484
transform -1 0 9632 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__165__CLK
timestamp 1666464484
transform 1 0 29232 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__165__D
timestamp 1666464484
transform -1 0 33152 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__166__CLK
timestamp 1666464484
transform 1 0 33488 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__167__CLK
timestamp 1666464484
transform 1 0 34048 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__167__D
timestamp 1666464484
transform -1 0 37968 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__168__CLK
timestamp 1666464484
transform -1 0 37408 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__169__CLK
timestamp 1666464484
transform 1 0 34832 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__169__D
timestamp 1666464484
transform 1 0 37520 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__170__CLK
timestamp 1666464484
transform -1 0 35280 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__170__D
timestamp 1666464484
transform 1 0 38976 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__171__CLK
timestamp 1666464484
transform 1 0 35168 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__172__CLK
timestamp 1666464484
transform 1 0 37184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__173__CLK
timestamp 1666464484
transform 1 0 34608 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__174__CLK
timestamp 1666464484
transform 1 0 33488 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__174__D
timestamp 1666464484
transform 1 0 37632 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__175__CLK
timestamp 1666464484
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__175__D
timestamp 1666464484
transform -1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__176__CLK
timestamp 1666464484
transform 1 0 33936 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__176__D
timestamp 1666464484
transform 1 0 33488 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__177__CLK
timestamp 1666464484
transform 1 0 29904 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__177__D
timestamp 1666464484
transform -1 0 29680 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__178__CLK
timestamp 1666464484
transform -1 0 29344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__178__D
timestamp 1666464484
transform 1 0 29680 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__179__CLK
timestamp 1666464484
transform -1 0 30240 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__179__D
timestamp 1666464484
transform -1 0 29792 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__180__CLK
timestamp 1666464484
transform 1 0 29456 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__180__D
timestamp 1666464484
transform 1 0 29008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__181__CLK
timestamp 1666464484
transform 1 0 23744 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__181__D
timestamp 1666464484
transform 1 0 24192 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__182__CLK
timestamp 1666464484
transform 1 0 17360 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__182__D
timestamp 1666464484
transform -1 0 21728 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__183__CLK
timestamp 1666464484
transform 1 0 16464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__183__D
timestamp 1666464484
transform -1 0 20608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__184__CLK
timestamp 1666464484
transform 1 0 13440 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__184__D
timestamp 1666464484
transform 1 0 17584 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__185__CLK
timestamp 1666464484
transform 1 0 15568 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__185__D
timestamp 1666464484
transform -1 0 19712 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__186__CLK
timestamp 1666464484
transform 1 0 16016 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__186__D
timestamp 1666464484
transform -1 0 20160 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__187__CLK
timestamp 1666464484
transform 1 0 17024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__187__D
timestamp 1666464484
transform 1 0 20720 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__188__CLK
timestamp 1666464484
transform 1 0 18928 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__188__D
timestamp 1666464484
transform 1 0 22848 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__189__CLK
timestamp 1666464484
transform 1 0 27888 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__189__D
timestamp 1666464484
transform -1 0 28672 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__190__CLK
timestamp 1666464484
transform 1 0 30800 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__191__CLK
timestamp 1666464484
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__192__CLK
timestamp 1666464484
transform 1 0 32928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__193__CLK
timestamp 1666464484
transform 1 0 32928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__194__CLK
timestamp 1666464484
transform 1 0 31808 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__195__CLK
timestamp 1666464484
transform 1 0 24752 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__196__CLK
timestamp 1666464484
transform 1 0 15904 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__196__D
timestamp 1666464484
transform 1 0 16352 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__205__I
timestamp 1666464484
transform 1 0 38864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__I
timestamp 1666464484
transform 1 0 17360 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clock_I
timestamp 1666464484
transform -1 0 19264 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_0__f_clock_I
timestamp 1666464484
transform 1 0 17584 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_1__f_clock_I
timestamp 1666464484
transform -1 0 17808 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_2__f_clock_I
timestamp 1666464484
transform 1 0 28672 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_3__f_clock_I
timestamp 1666464484
transform 1 0 26208 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1666464484
transform -1 0 1904 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1666464484
transform -1 0 1904 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1666464484
transform -1 0 1904 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output4_I
timestamp 1666464484
transform 1 0 47152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output5_I
timestamp 1666464484
transform -1 0 46480 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output6_I
timestamp 1666464484
transform -1 0 46480 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output7_I
timestamp 1666464484
transform 1 0 46256 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output8_I
timestamp 1666464484
transform 1 0 46256 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output9_I
timestamp 1666464484
transform 1 0 46256 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output10_I
timestamp 1666464484
transform 1 0 46256 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output11_I
timestamp 1666464484
transform 1 0 46256 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output12_I
timestamp 1666464484
transform 1 0 46256 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output13_I
timestamp 1666464484
transform 1 0 46256 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output14_I
timestamp 1666464484
transform -1 0 46480 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output15_I
timestamp 1666464484
transform -1 0 46480 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output16_I
timestamp 1666464484
transform -1 0 46480 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output17_I
timestamp 1666464484
transform -1 0 46480 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output18_I
timestamp 1666464484
transform -1 0 46480 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output19_I
timestamp 1666464484
transform -1 0 46480 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output20_I
timestamp 1666464484
transform -1 0 46480 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output21_I
timestamp 1666464484
transform -1 0 46480 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output22_I
timestamp 1666464484
transform 1 0 46256 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output23_I
timestamp 1666464484
transform 1 0 46256 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output24_I
timestamp 1666464484
transform 1 0 46256 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output25_I
timestamp 1666464484
transform 1 0 46256 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output26_I
timestamp 1666464484
transform 1 0 45808 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output27_I
timestamp 1666464484
transform 1 0 46256 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output28_I
timestamp 1666464484
transform -1 0 46480 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output29_I
timestamp 1666464484
transform 1 0 44128 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output30_I
timestamp 1666464484
transform 1 0 46256 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output31_I
timestamp 1666464484
transform -1 0 46480 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output32_I
timestamp 1666464484
transform 1 0 46256 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output33_I
timestamp 1666464484
transform 1 0 46256 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output34_I
timestamp 1666464484
transform 1 0 46256 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output35_I
timestamp 1666464484
transform 1 0 46256 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output36_I
timestamp 1666464484
transform -1 0 46480 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output37_I
timestamp 1666464484
transform 1 0 3472 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 1568 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 2352 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 4144 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 5040 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37
timestamp 1666464484
transform 1 0 5488 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53
timestamp 1666464484
transform 1 0 7280 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61
timestamp 1666464484
transform 1 0 8176 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63
timestamp 1666464484
transform 1 0 8400 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68
timestamp 1666464484
transform 1 0 8960 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_72 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 9408 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1666464484
transform 1 0 12992 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_107 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 13328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_111
timestamp 1666464484
transform 1 0 13776 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_117
timestamp 1666464484
transform 1 0 14448 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_133
timestamp 1666464484
transform 1 0 16240 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_137
timestamp 1666464484
transform 1 0 16688 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_139
timestamp 1666464484
transform 1 0 16912 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_142
timestamp 1666464484
transform 1 0 17248 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_158
timestamp 1666464484
transform 1 0 19040 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_166
timestamp 1666464484
transform 1 0 19936 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_174
timestamp 1666464484
transform 1 0 20832 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_177
timestamp 1666464484
transform 1 0 21168 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_193
timestamp 1666464484
transform 1 0 22960 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_201
timestamp 1666464484
transform 1 0 23856 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_209
timestamp 1666464484
transform 1 0 24752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_212
timestamp 1666464484
transform 1 0 25088 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_214
timestamp 1666464484
transform 1 0 25312 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_244
timestamp 1666464484
transform 1 0 28672 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_247
timestamp 1666464484
transform 1 0 29008 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_250
timestamp 1666464484
transform 1 0 29344 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_254
timestamp 1666464484
transform 1 0 29792 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_258
timestamp 1666464484
transform 1 0 30240 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_274
timestamp 1666464484
transform 1 0 32032 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_278
timestamp 1666464484
transform 1 0 32480 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_282
timestamp 1666464484
transform 1 0 32928 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_314
timestamp 1666464484
transform 1 0 36512 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_317
timestamp 1666464484
transform 1 0 36848 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_319
timestamp 1666464484
transform 1 0 37072 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_322
timestamp 1666464484
transform 1 0 37408 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_324
timestamp 1666464484
transform 1 0 37632 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_327
timestamp 1666464484
transform 1 0 37968 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_343
timestamp 1666464484
transform 1 0 39760 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_347
timestamp 1666464484
transform 1 0 40208 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_349
timestamp 1666464484
transform 1 0 40432 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_352
timestamp 1666464484
transform 1 0 40768 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_384
timestamp 1666464484
transform 1 0 44352 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_387
timestamp 1666464484
transform 1 0 44688 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_395
timestamp 1666464484
transform 1 0 45584 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_399
timestamp 1666464484
transform 1 0 46032 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_403
timestamp 1666464484
transform 1 0 46480 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_419
timestamp 1666464484
transform 1 0 48272 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_2
timestamp 1666464484
transform 1 0 1568 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_5 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 1904 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_69
timestamp 1666464484
transform 1 0 9072 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_73
timestamp 1666464484
transform 1 0 9520 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_137
timestamp 1666464484
transform 1 0 16688 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_141
timestamp 1666464484
transform 1 0 17136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_144
timestamp 1666464484
transform 1 0 17472 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_160
timestamp 1666464484
transform 1 0 19264 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_168
timestamp 1666464484
transform 1 0 20160 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_198
timestamp 1666464484
transform 1 0 23520 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_202
timestamp 1666464484
transform 1 0 23968 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_206
timestamp 1666464484
transform 1 0 24416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_210
timestamp 1666464484
transform 1 0 24864 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_212
timestamp 1666464484
transform 1 0 25088 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_215
timestamp 1666464484
transform 1 0 25424 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_245
timestamp 1666464484
transform 1 0 28784 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_251
timestamp 1666464484
transform 1 0 29456 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_255
timestamp 1666464484
transform 1 0 29904 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_271
timestamp 1666464484
transform 1 0 31696 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_279
timestamp 1666464484
transform 1 0 32592 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_283
timestamp 1666464484
transform 1 0 33040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_286
timestamp 1666464484
transform 1 0 33376 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_289
timestamp 1666464484
transform 1 0 33712 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_291
timestamp 1666464484
transform 1 0 33936 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_294
timestamp 1666464484
transform 1 0 34272 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_325
timestamp 1666464484
transform 1 0 37744 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_333
timestamp 1666464484
transform 1 0 38640 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_337
timestamp 1666464484
transform 1 0 39088 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_345
timestamp 1666464484
transform 1 0 39984 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_348
timestamp 1666464484
transform 1 0 40320 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_352
timestamp 1666464484
transform 1 0 40768 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_354
timestamp 1666464484
transform 1 0 40992 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_357
timestamp 1666464484
transform 1 0 41328 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_360
timestamp 1666464484
transform 1 0 41664 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_364
timestamp 1666464484
transform 1 0 42112 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_370
timestamp 1666464484
transform 1 0 42784 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_402
timestamp 1666464484
transform 1 0 46368 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_406
timestamp 1666464484
transform 1 0 46816 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_408
timestamp 1666464484
transform 1 0 47040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_411
timestamp 1666464484
transform 1 0 47376 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_419
timestamp 1666464484
transform 1 0 48272 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_2
timestamp 1666464484
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1666464484
transform 1 0 5152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_37
timestamp 1666464484
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_101
timestamp 1666464484
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1666464484
transform 1 0 13104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_108
timestamp 1666464484
transform 1 0 13440 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_124
timestamp 1666464484
transform 1 0 15232 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_132
timestamp 1666464484
transform 1 0 16128 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_136
timestamp 1666464484
transform 1 0 16576 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_140
timestamp 1666464484
transform 1 0 17024 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_171
timestamp 1666464484
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_175
timestamp 1666464484
transform 1 0 20944 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_179
timestamp 1666464484
transform 1 0 21392 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_187
timestamp 1666464484
transform 1 0 22288 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_191
timestamp 1666464484
transform 1 0 22736 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_242
timestamp 1666464484
transform 1 0 28448 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_246
timestamp 1666464484
transform 1 0 28896 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_250
timestamp 1666464484
transform 1 0 29344 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_280
timestamp 1666464484
transform 1 0 32704 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_284
timestamp 1666464484
transform 1 0 33152 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_288
timestamp 1666464484
transform 1 0 33600 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_318
timestamp 1666464484
transform 1 0 36960 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_321
timestamp 1666464484
transform 1 0 37296 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_351
timestamp 1666464484
transform 1 0 40656 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_368
timestamp 1666464484
transform 1 0 42560 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_376
timestamp 1666464484
transform 1 0 43456 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_380
timestamp 1666464484
transform 1 0 43904 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_388
timestamp 1666464484
transform 1 0 44800 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_392
timestamp 1666464484
transform 1 0 45248 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_400
timestamp 1666464484
transform 1 0 46144 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_403
timestamp 1666464484
transform 1 0 46480 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_419
timestamp 1666464484
transform 1 0 48272 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_2
timestamp 1666464484
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_66
timestamp 1666464484
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1666464484
transform 1 0 9184 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_73
timestamp 1666464484
transform 1 0 9520 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_89
timestamp 1666464484
transform 1 0 11312 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_97
timestamp 1666464484
transform 1 0 12208 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_128
timestamp 1666464484
transform 1 0 15680 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_132
timestamp 1666464484
transform 1 0 16128 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_136
timestamp 1666464484
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_140
timestamp 1666464484
transform 1 0 17024 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_144
timestamp 1666464484
transform 1 0 17472 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_208
timestamp 1666464484
transform 1 0 24640 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_212
timestamp 1666464484
transform 1 0 25088 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_215
timestamp 1666464484
transform 1 0 25424 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_245
timestamp 1666464484
transform 1 0 28784 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_249
timestamp 1666464484
transform 1 0 29232 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_253
timestamp 1666464484
transform 1 0 29680 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_269
timestamp 1666464484
transform 1 0 31472 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_277
timestamp 1666464484
transform 1 0 32368 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_281
timestamp 1666464484
transform 1 0 32816 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_283
timestamp 1666464484
transform 1 0 33040 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_286
timestamp 1666464484
transform 1 0 33376 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_294
timestamp 1666464484
transform 1 0 34272 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_298
timestamp 1666464484
transform 1 0 34720 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_301
timestamp 1666464484
transform 1 0 35056 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_332
timestamp 1666464484
transform 1 0 38528 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_334
timestamp 1666464484
transform 1 0 38752 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_350
timestamp 1666464484
transform 1 0 40544 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_354
timestamp 1666464484
transform 1 0 40992 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_357
timestamp 1666464484
transform 1 0 41328 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_373
timestamp 1666464484
transform 1 0 43120 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_381
timestamp 1666464484
transform 1 0 44016 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_389
timestamp 1666464484
transform 1 0 44912 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_405
timestamp 1666464484
transform 1 0 46704 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_413
timestamp 1666464484
transform 1 0 47600 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_417
timestamp 1666464484
transform 1 0 48048 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_419
timestamp 1666464484
transform 1 0 48272 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_2
timestamp 1666464484
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1666464484
transform 1 0 5152 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_37
timestamp 1666464484
transform 1 0 5488 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_69
timestamp 1666464484
transform 1 0 9072 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_85
timestamp 1666464484
transform 1 0 10864 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_93
timestamp 1666464484
transform 1 0 11760 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_97
timestamp 1666464484
transform 1 0 12208 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_101
timestamp 1666464484
transform 1 0 12656 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1666464484
transform 1 0 13104 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_108
timestamp 1666464484
transform 1 0 13440 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_138
timestamp 1666464484
transform 1 0 16800 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_142
timestamp 1666464484
transform 1 0 17248 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_145
timestamp 1666464484
transform 1 0 17584 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_176
timestamp 1666464484
transform 1 0 21056 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_179
timestamp 1666464484
transform 1 0 21392 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_182
timestamp 1666464484
transform 1 0 21728 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_214
timestamp 1666464484
transform 1 0 25312 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_247
timestamp 1666464484
transform 1 0 29008 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_250
timestamp 1666464484
transform 1 0 29344 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_253
timestamp 1666464484
transform 1 0 29680 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_257
timestamp 1666464484
transform 1 0 30128 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_289
timestamp 1666464484
transform 1 0 33712 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_305
timestamp 1666464484
transform 1 0 35504 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_313
timestamp 1666464484
transform 1 0 36400 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_317
timestamp 1666464484
transform 1 0 36848 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_321
timestamp 1666464484
transform 1 0 37296 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_325
timestamp 1666464484
transform 1 0 37744 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_329
timestamp 1666464484
transform 1 0 38192 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_333
timestamp 1666464484
transform 1 0 38640 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_337
timestamp 1666464484
transform 1 0 39088 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_354
timestamp 1666464484
transform 1 0 40992 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_371
timestamp 1666464484
transform 1 0 42896 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_379
timestamp 1666464484
transform 1 0 43792 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_387
timestamp 1666464484
transform 1 0 44688 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_389
timestamp 1666464484
transform 1 0 44912 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_392
timestamp 1666464484
transform 1 0 45248 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_400
timestamp 1666464484
transform 1 0 46144 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_403
timestamp 1666464484
transform 1 0 46480 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_419
timestamp 1666464484
transform 1 0 48272 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_2
timestamp 1666464484
transform 1 0 1568 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_36
timestamp 1666464484
transform 1 0 5376 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_40
timestamp 1666464484
transform 1 0 5824 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1666464484
transform 1 0 9184 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_73
timestamp 1666464484
transform 1 0 9520 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_76
timestamp 1666464484
transform 1 0 9856 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_84
timestamp 1666464484
transform 1 0 10752 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_88
timestamp 1666464484
transform 1 0 11200 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_140
timestamp 1666464484
transform 1 0 17024 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_144
timestamp 1666464484
transform 1 0 17472 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_147
timestamp 1666464484
transform 1 0 17808 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_211
timestamp 1666464484
transform 1 0 24976 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_215
timestamp 1666464484
transform 1 0 25424 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_219
timestamp 1666464484
transform 1 0 25872 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_221
timestamp 1666464484
transform 1 0 26096 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_224
timestamp 1666464484
transform 1 0 26432 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_276
timestamp 1666464484
transform 1 0 32256 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_286
timestamp 1666464484
transform 1 0 33376 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_294
timestamp 1666464484
transform 1 0 34272 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_298
timestamp 1666464484
transform 1 0 34720 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_300
timestamp 1666464484
transform 1 0 34944 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_303
timestamp 1666464484
transform 1 0 35280 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_334
timestamp 1666464484
transform 1 0 38752 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_338
timestamp 1666464484
transform 1 0 39200 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_346
timestamp 1666464484
transform 1 0 40096 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_350
timestamp 1666464484
transform 1 0 40544 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_354
timestamp 1666464484
transform 1 0 40992 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_357
timestamp 1666464484
transform 1 0 41328 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_360
timestamp 1666464484
transform 1 0 41664 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_364
timestamp 1666464484
transform 1 0 42112 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_368
timestamp 1666464484
transform 1 0 42560 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_371
timestamp 1666464484
transform 1 0 42896 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_375
timestamp 1666464484
transform 1 0 43344 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_385
timestamp 1666464484
transform 1 0 44464 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_417
timestamp 1666464484
transform 1 0 48048 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_419
timestamp 1666464484
transform 1 0 48272 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_2
timestamp 1666464484
transform 1 0 1568 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_4
timestamp 1666464484
transform 1 0 1792 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1666464484
transform 1 0 5152 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_37
timestamp 1666464484
transform 1 0 5488 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_67
timestamp 1666464484
transform 1 0 8848 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_71
timestamp 1666464484
transform 1 0 9296 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_74
timestamp 1666464484
transform 1 0 9632 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_105
timestamp 1666464484
transform 1 0 13104 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_108
timestamp 1666464484
transform 1 0 13440 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_111
timestamp 1666464484
transform 1 0 13776 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_127
timestamp 1666464484
transform 1 0 15568 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_137
timestamp 1666464484
transform 1 0 16688 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_168
timestamp 1666464484
transform 1 0 20160 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_172
timestamp 1666464484
transform 1 0 20608 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_176
timestamp 1666464484
transform 1 0 21056 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_179
timestamp 1666464484
transform 1 0 21392 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_243
timestamp 1666464484
transform 1 0 28560 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_247
timestamp 1666464484
transform 1 0 29008 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_250
timestamp 1666464484
transform 1 0 29344 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_314
timestamp 1666464484
transform 1 0 36512 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_318
timestamp 1666464484
transform 1 0 36960 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_321
timestamp 1666464484
transform 1 0 37296 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_337
timestamp 1666464484
transform 1 0 39088 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_345
timestamp 1666464484
transform 1 0 39984 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_349
timestamp 1666464484
transform 1 0 40432 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_353
timestamp 1666464484
transform 1 0 40880 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_357
timestamp 1666464484
transform 1 0 41328 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_374
timestamp 1666464484
transform 1 0 43232 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_392
timestamp 1666464484
transform 1 0 45248 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_400
timestamp 1666464484
transform 1 0 46144 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_403
timestamp 1666464484
transform 1 0 46480 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_419
timestamp 1666464484
transform 1 0 48272 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_2
timestamp 1666464484
transform 1 0 1568 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_7
timestamp 1666464484
transform 1 0 2128 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_11
timestamp 1666464484
transform 1 0 2576 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_13
timestamp 1666464484
transform 1 0 2800 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_16
timestamp 1666464484
transform 1 0 3136 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_47
timestamp 1666464484
transform 1 0 6608 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_51
timestamp 1666464484
transform 1 0 7056 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_69
timestamp 1666464484
transform 1 0 9072 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_73
timestamp 1666464484
transform 1 0 9520 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_89
timestamp 1666464484
transform 1 0 11312 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_140
timestamp 1666464484
transform 1 0 17024 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_144
timestamp 1666464484
transform 1 0 17472 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_147
timestamp 1666464484
transform 1 0 17808 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_155
timestamp 1666464484
transform 1 0 18704 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_157
timestamp 1666464484
transform 1 0 18928 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_160
timestamp 1666464484
transform 1 0 19264 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_212
timestamp 1666464484
transform 1 0 25088 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_215
timestamp 1666464484
transform 1 0 25424 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_247
timestamp 1666464484
transform 1 0 29008 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_251
timestamp 1666464484
transform 1 0 29456 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_253
timestamp 1666464484
transform 1 0 29680 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_283
timestamp 1666464484
transform 1 0 33040 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_286
timestamp 1666464484
transform 1 0 33376 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_289
timestamp 1666464484
transform 1 0 33712 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_293
timestamp 1666464484
transform 1 0 34160 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_301
timestamp 1666464484
transform 1 0 35056 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_304
timestamp 1666464484
transform 1 0 35392 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_335
timestamp 1666464484
transform 1 0 38864 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_351
timestamp 1666464484
transform 1 0 40656 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_357
timestamp 1666464484
transform 1 0 41328 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_389
timestamp 1666464484
transform 1 0 44912 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_397
timestamp 1666464484
transform 1 0 45808 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_403
timestamp 1666464484
transform 1 0 46480 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_419
timestamp 1666464484
transform 1 0 48272 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_2
timestamp 1666464484
transform 1 0 1568 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_4
timestamp 1666464484
transform 1 0 1792 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1666464484
transform 1 0 5152 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_37
timestamp 1666464484
transform 1 0 5488 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_40
timestamp 1666464484
transform 1 0 5824 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_104
timestamp 1666464484
transform 1 0 12992 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_108
timestamp 1666464484
transform 1 0 13440 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_124
timestamp 1666464484
transform 1 0 15232 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_128
timestamp 1666464484
transform 1 0 15680 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_130
timestamp 1666464484
transform 1 0 15904 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_133
timestamp 1666464484
transform 1 0 16240 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_164
timestamp 1666464484
transform 1 0 19712 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_168
timestamp 1666464484
transform 1 0 20160 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_176
timestamp 1666464484
transform 1 0 21056 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_179
timestamp 1666464484
transform 1 0 21392 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_243
timestamp 1666464484
transform 1 0 28560 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_247
timestamp 1666464484
transform 1 0 29008 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_250
timestamp 1666464484
transform 1 0 29344 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_280
timestamp 1666464484
transform 1 0 32704 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_284
timestamp 1666464484
transform 1 0 33152 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_286
timestamp 1666464484
transform 1 0 33376 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_289
timestamp 1666464484
transform 1 0 33712 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_305
timestamp 1666464484
transform 1 0 35504 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_313
timestamp 1666464484
transform 1 0 36400 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_317
timestamp 1666464484
transform 1 0 36848 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_321
timestamp 1666464484
transform 1 0 37296 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_353
timestamp 1666464484
transform 1 0 40880 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_355
timestamp 1666464484
transform 1 0 41104 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_358
timestamp 1666464484
transform 1 0 41440 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_362
timestamp 1666464484
transform 1 0 41888 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_369
timestamp 1666464484
transform 1 0 42672 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_385
timestamp 1666464484
transform 1 0 44464 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_389
timestamp 1666464484
transform 1 0 44912 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_392
timestamp 1666464484
transform 1 0 45248 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_408
timestamp 1666464484
transform 1 0 47040 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_416
timestamp 1666464484
transform 1 0 47936 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_2
timestamp 1666464484
transform 1 0 1568 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_10
timestamp 1666464484
transform 1 0 2464 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_12
timestamp 1666464484
transform 1 0 2688 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_15
timestamp 1666464484
transform 1 0 3024 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_46
timestamp 1666464484
transform 1 0 6496 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_50
timestamp 1666464484
transform 1 0 6944 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_66
timestamp 1666464484
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_70
timestamp 1666464484
transform 1 0 9184 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_73
timestamp 1666464484
transform 1 0 9520 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_105
timestamp 1666464484
transform 1 0 13104 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_107
timestamp 1666464484
transform 1 0 13328 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_110
timestamp 1666464484
transform 1 0 13664 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_141
timestamp 1666464484
transform 1 0 17136 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_144
timestamp 1666464484
transform 1 0 17472 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_147
timestamp 1666464484
transform 1 0 17808 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_155
timestamp 1666464484
transform 1 0 18704 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_159
timestamp 1666464484
transform 1 0 19152 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_190
timestamp 1666464484
transform 1 0 22624 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_194
timestamp 1666464484
transform 1 0 23072 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_202
timestamp 1666464484
transform 1 0 23968 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_206
timestamp 1666464484
transform 1 0 24416 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_208
timestamp 1666464484
transform 1 0 24640 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_211
timestamp 1666464484
transform 1 0 24976 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_215
timestamp 1666464484
transform 1 0 25424 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_231
timestamp 1666464484
transform 1 0 27216 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_261
timestamp 1666464484
transform 1 0 30576 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_265
timestamp 1666464484
transform 1 0 31024 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_273
timestamp 1666464484
transform 1 0 31920 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_277
timestamp 1666464484
transform 1 0 32368 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_279
timestamp 1666464484
transform 1 0 32592 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_282
timestamp 1666464484
transform 1 0 32928 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_286
timestamp 1666464484
transform 1 0 33376 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_288
timestamp 1666464484
transform 1 0 33600 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_318
timestamp 1666464484
transform 1 0 36960 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_322
timestamp 1666464484
transform 1 0 37408 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_326
timestamp 1666464484
transform 1 0 37856 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_342
timestamp 1666464484
transform 1 0 39648 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_350
timestamp 1666464484
transform 1 0 40544 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_354
timestamp 1666464484
transform 1 0 40992 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_357
timestamp 1666464484
transform 1 0 41328 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_373
timestamp 1666464484
transform 1 0 43120 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_389
timestamp 1666464484
transform 1 0 44912 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_397
timestamp 1666464484
transform 1 0 45808 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_403
timestamp 1666464484
transform 1 0 46480 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_419
timestamp 1666464484
transform 1 0 48272 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_2
timestamp 1666464484
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1666464484
transform 1 0 5152 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_37
timestamp 1666464484
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_101
timestamp 1666464484
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1666464484
transform 1 0 13104 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_108
timestamp 1666464484
transform 1 0 13440 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_142
timestamp 1666464484
transform 1 0 17248 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_173
timestamp 1666464484
transform 1 0 20720 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_179
timestamp 1666464484
transform 1 0 21392 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_209
timestamp 1666464484
transform 1 0 24752 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_240
timestamp 1666464484
transform 1 0 28224 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_244
timestamp 1666464484
transform 1 0 28672 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_250
timestamp 1666464484
transform 1 0 29344 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_280
timestamp 1666464484
transform 1 0 32704 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_311
timestamp 1666464484
transform 1 0 36176 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_315
timestamp 1666464484
transform 1 0 36624 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_321
timestamp 1666464484
transform 1 0 37296 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_351
timestamp 1666464484
transform 1 0 40656 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_353
timestamp 1666464484
transform 1 0 40880 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_356
timestamp 1666464484
transform 1 0 41216 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_368
timestamp 1666464484
transform 1 0 42560 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_376
timestamp 1666464484
transform 1 0 43456 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_384
timestamp 1666464484
transform 1 0 44352 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_388
timestamp 1666464484
transform 1 0 44800 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_392
timestamp 1666464484
transform 1 0 45248 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_408
timestamp 1666464484
transform 1 0 47040 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_416
timestamp 1666464484
transform 1 0 47936 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_2
timestamp 1666464484
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_66
timestamp 1666464484
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_70
timestamp 1666464484
transform 1 0 9184 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_73
timestamp 1666464484
transform 1 0 9520 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_137
timestamp 1666464484
transform 1 0 16688 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_141
timestamp 1666464484
transform 1 0 17136 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_144
timestamp 1666464484
transform 1 0 17472 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_160
timestamp 1666464484
transform 1 0 19264 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_168
timestamp 1666464484
transform 1 0 20160 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_172
timestamp 1666464484
transform 1 0 20608 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_175
timestamp 1666464484
transform 1 0 20944 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_207
timestamp 1666464484
transform 1 0 24528 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_211
timestamp 1666464484
transform 1 0 24976 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_215
timestamp 1666464484
transform 1 0 25424 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_231
timestamp 1666464484
transform 1 0 27216 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_235
timestamp 1666464484
transform 1 0 27664 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_239
timestamp 1666464484
transform 1 0 28112 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_270
timestamp 1666464484
transform 1 0 31584 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_274
timestamp 1666464484
transform 1 0 32032 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_278
timestamp 1666464484
transform 1 0 32480 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_282
timestamp 1666464484
transform 1 0 32928 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_286
timestamp 1666464484
transform 1 0 33376 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_294
timestamp 1666464484
transform 1 0 34272 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_296
timestamp 1666464484
transform 1 0 34496 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_299
timestamp 1666464484
transform 1 0 34832 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_330
timestamp 1666464484
transform 1 0 38304 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_346
timestamp 1666464484
transform 1 0 40096 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_354
timestamp 1666464484
transform 1 0 40992 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_357
timestamp 1666464484
transform 1 0 41328 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_373
timestamp 1666464484
transform 1 0 43120 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_377
timestamp 1666464484
transform 1 0 43568 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_393
timestamp 1666464484
transform 1 0 45360 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_403
timestamp 1666464484
transform 1 0 46480 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_419
timestamp 1666464484
transform 1 0 48272 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_2
timestamp 1666464484
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1666464484
transform 1 0 5152 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_37
timestamp 1666464484
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_101
timestamp 1666464484
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_105
timestamp 1666464484
transform 1 0 13104 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_108
timestamp 1666464484
transform 1 0 13440 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_124
timestamp 1666464484
transform 1 0 15232 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_126
timestamp 1666464484
transform 1 0 15456 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_129
timestamp 1666464484
transform 1 0 15792 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_160
timestamp 1666464484
transform 1 0 19264 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_164
timestamp 1666464484
transform 1 0 19712 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_172
timestamp 1666464484
transform 1 0 20608 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_176
timestamp 1666464484
transform 1 0 21056 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_179
timestamp 1666464484
transform 1 0 21392 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_243
timestamp 1666464484
transform 1 0 28560 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_247
timestamp 1666464484
transform 1 0 29008 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_250
timestamp 1666464484
transform 1 0 29344 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_280
timestamp 1666464484
transform 1 0 32704 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_284
timestamp 1666464484
transform 1 0 33152 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_300
timestamp 1666464484
transform 1 0 34944 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_308
timestamp 1666464484
transform 1 0 35840 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_312
timestamp 1666464484
transform 1 0 36288 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_314
timestamp 1666464484
transform 1 0 36512 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_317
timestamp 1666464484
transform 1 0 36848 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_321
timestamp 1666464484
transform 1 0 37296 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_324
timestamp 1666464484
transform 1 0 37632 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_334
timestamp 1666464484
transform 1 0 38752 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_342
timestamp 1666464484
transform 1 0 39648 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_346
timestamp 1666464484
transform 1 0 40096 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_354
timestamp 1666464484
transform 1 0 40992 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_364
timestamp 1666464484
transform 1 0 42112 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_380
timestamp 1666464484
transform 1 0 43904 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_388
timestamp 1666464484
transform 1 0 44800 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_392
timestamp 1666464484
transform 1 0 45248 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_408
timestamp 1666464484
transform 1 0 47040 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_416
timestamp 1666464484
transform 1 0 47936 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_2
timestamp 1666464484
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_66
timestamp 1666464484
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_70
timestamp 1666464484
transform 1 0 9184 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_73
timestamp 1666464484
transform 1 0 9520 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_137
timestamp 1666464484
transform 1 0 16688 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_141
timestamp 1666464484
transform 1 0 17136 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_144
timestamp 1666464484
transform 1 0 17472 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_208
timestamp 1666464484
transform 1 0 24640 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_212
timestamp 1666464484
transform 1 0 25088 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_215
timestamp 1666464484
transform 1 0 25424 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_279
timestamp 1666464484
transform 1 0 32592 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_283
timestamp 1666464484
transform 1 0 33040 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_286
timestamp 1666464484
transform 1 0 33376 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_290
timestamp 1666464484
transform 1 0 33824 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_294
timestamp 1666464484
transform 1 0 34272 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_302
timestamp 1666464484
transform 1 0 35168 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_306
timestamp 1666464484
transform 1 0 35616 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_308
timestamp 1666464484
transform 1 0 35840 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_311
timestamp 1666464484
transform 1 0 36176 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_315
timestamp 1666464484
transform 1 0 36624 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_332
timestamp 1666464484
transform 1 0 38528 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_349
timestamp 1666464484
transform 1 0 40432 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_353
timestamp 1666464484
transform 1 0 40880 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_357
timestamp 1666464484
transform 1 0 41328 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_389
timestamp 1666464484
transform 1 0 44912 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_397
timestamp 1666464484
transform 1 0 45808 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_403
timestamp 1666464484
transform 1 0 46480 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_419
timestamp 1666464484
transform 1 0 48272 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_2
timestamp 1666464484
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_34
timestamp 1666464484
transform 1 0 5152 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_37
timestamp 1666464484
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_101
timestamp 1666464484
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_105
timestamp 1666464484
transform 1 0 13104 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_108
timestamp 1666464484
transform 1 0 13440 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_172
timestamp 1666464484
transform 1 0 20608 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_176
timestamp 1666464484
transform 1 0 21056 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_179
timestamp 1666464484
transform 1 0 21392 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_243
timestamp 1666464484
transform 1 0 28560 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_247
timestamp 1666464484
transform 1 0 29008 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_250
timestamp 1666464484
transform 1 0 29344 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_282
timestamp 1666464484
transform 1 0 32928 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_284
timestamp 1666464484
transform 1 0 33152 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_287
timestamp 1666464484
transform 1 0 33488 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_291
timestamp 1666464484
transform 1 0 33936 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_293
timestamp 1666464484
transform 1 0 34160 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_309
timestamp 1666464484
transform 1 0 35952 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_313
timestamp 1666464484
transform 1 0 36400 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_315
timestamp 1666464484
transform 1 0 36624 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_318
timestamp 1666464484
transform 1 0 36960 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_321
timestamp 1666464484
transform 1 0 37296 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_337
timestamp 1666464484
transform 1 0 39088 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_347
timestamp 1666464484
transform 1 0 40208 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_357
timestamp 1666464484
transform 1 0 41328 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_389
timestamp 1666464484
transform 1 0 44912 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_392
timestamp 1666464484
transform 1 0 45248 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_408
timestamp 1666464484
transform 1 0 47040 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_416
timestamp 1666464484
transform 1 0 47936 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_2
timestamp 1666464484
transform 1 0 1568 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_5
timestamp 1666464484
transform 1 0 1904 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_69
timestamp 1666464484
transform 1 0 9072 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_73
timestamp 1666464484
transform 1 0 9520 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_137
timestamp 1666464484
transform 1 0 16688 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_141
timestamp 1666464484
transform 1 0 17136 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_144
timestamp 1666464484
transform 1 0 17472 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_208
timestamp 1666464484
transform 1 0 24640 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_212
timestamp 1666464484
transform 1 0 25088 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_215
timestamp 1666464484
transform 1 0 25424 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_253
timestamp 1666464484
transform 1 0 29680 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_257
timestamp 1666464484
transform 1 0 30128 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_261
timestamp 1666464484
transform 1 0 30576 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_264
timestamp 1666464484
transform 1 0 30912 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_280
timestamp 1666464484
transform 1 0 32704 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_286
timestamp 1666464484
transform 1 0 33376 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_289
timestamp 1666464484
transform 1 0 33712 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_306
timestamp 1666464484
transform 1 0 35616 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_323
timestamp 1666464484
transform 1 0 37520 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_340
timestamp 1666464484
transform 1 0 39424 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_352
timestamp 1666464484
transform 1 0 40768 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_354
timestamp 1666464484
transform 1 0 40992 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_357
timestamp 1666464484
transform 1 0 41328 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_360
timestamp 1666464484
transform 1 0 41664 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_392
timestamp 1666464484
transform 1 0 45248 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_400
timestamp 1666464484
transform 1 0 46144 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_403
timestamp 1666464484
transform 1 0 46480 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_419
timestamp 1666464484
transform 1 0 48272 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_2
timestamp 1666464484
transform 1 0 1568 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_9
timestamp 1666464484
transform 1 0 2352 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_25
timestamp 1666464484
transform 1 0 4144 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_33
timestamp 1666464484
transform 1 0 5040 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_37
timestamp 1666464484
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_101
timestamp 1666464484
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_105
timestamp 1666464484
transform 1 0 13104 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_108
timestamp 1666464484
transform 1 0 13440 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_172
timestamp 1666464484
transform 1 0 20608 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_176
timestamp 1666464484
transform 1 0 21056 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_179
timestamp 1666464484
transform 1 0 21392 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_211
timestamp 1666464484
transform 1 0 24976 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_227
timestamp 1666464484
transform 1 0 26768 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_235
timestamp 1666464484
transform 1 0 27664 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_239
timestamp 1666464484
transform 1 0 28112 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_247
timestamp 1666464484
transform 1 0 29008 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_250
timestamp 1666464484
transform 1 0 29344 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_254
timestamp 1666464484
transform 1 0 29792 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_262
timestamp 1666464484
transform 1 0 30688 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_270
timestamp 1666464484
transform 1 0 31584 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_274
timestamp 1666464484
transform 1 0 32032 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_278
timestamp 1666464484
transform 1 0 32480 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_280
timestamp 1666464484
transform 1 0 32704 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_283
timestamp 1666464484
transform 1 0 33040 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_287
timestamp 1666464484
transform 1 0 33488 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_304
timestamp 1666464484
transform 1 0 35392 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_308
timestamp 1666464484
transform 1 0 35840 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_316
timestamp 1666464484
transform 1 0 36736 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_318
timestamp 1666464484
transform 1 0 36960 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_321
timestamp 1666464484
transform 1 0 37296 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_324
timestamp 1666464484
transform 1 0 37632 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_328
timestamp 1666464484
transform 1 0 38080 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_332
timestamp 1666464484
transform 1 0 38528 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_336
timestamp 1666464484
transform 1 0 38976 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_340
timestamp 1666464484
transform 1 0 39424 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_347
timestamp 1666464484
transform 1 0 40208 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_355
timestamp 1666464484
transform 1 0 41104 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_387
timestamp 1666464484
transform 1 0 44688 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_389
timestamp 1666464484
transform 1 0 44912 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_392
timestamp 1666464484
transform 1 0 45248 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_408
timestamp 1666464484
transform 1 0 47040 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_416
timestamp 1666464484
transform 1 0 47936 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_2
timestamp 1666464484
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_66
timestamp 1666464484
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_70
timestamp 1666464484
transform 1 0 9184 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_73
timestamp 1666464484
transform 1 0 9520 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_137
timestamp 1666464484
transform 1 0 16688 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_141
timestamp 1666464484
transform 1 0 17136 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_144
timestamp 1666464484
transform 1 0 17472 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_208
timestamp 1666464484
transform 1 0 24640 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_212
timestamp 1666464484
transform 1 0 25088 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_17_215
timestamp 1666464484
transform 1 0 25424 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_247
timestamp 1666464484
transform 1 0 29008 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_263
timestamp 1666464484
transform 1 0 30800 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_271
timestamp 1666464484
transform 1 0 31696 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_275
timestamp 1666464484
transform 1 0 32144 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_283
timestamp 1666464484
transform 1 0 33040 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_286
timestamp 1666464484
transform 1 0 33376 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_296
timestamp 1666464484
transform 1 0 34496 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_300
timestamp 1666464484
transform 1 0 34944 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_317
timestamp 1666464484
transform 1 0 36848 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_334
timestamp 1666464484
transform 1 0 38752 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_342
timestamp 1666464484
transform 1 0 39648 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_350
timestamp 1666464484
transform 1 0 40544 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_354
timestamp 1666464484
transform 1 0 40992 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_357
timestamp 1666464484
transform 1 0 41328 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_17_364
timestamp 1666464484
transform 1 0 42112 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_396
timestamp 1666464484
transform 1 0 45696 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_400
timestamp 1666464484
transform 1 0 46144 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_403
timestamp 1666464484
transform 1 0 46480 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_419
timestamp 1666464484
transform 1 0 48272 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_18_2
timestamp 1666464484
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_34
timestamp 1666464484
transform 1 0 5152 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_37
timestamp 1666464484
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_101
timestamp 1666464484
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_105
timestamp 1666464484
transform 1 0 13104 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_108
timestamp 1666464484
transform 1 0 13440 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_172
timestamp 1666464484
transform 1 0 20608 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_176
timestamp 1666464484
transform 1 0 21056 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_179
timestamp 1666464484
transform 1 0 21392 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_243
timestamp 1666464484
transform 1 0 28560 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_247
timestamp 1666464484
transform 1 0 29008 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_250
timestamp 1666464484
transform 1 0 29344 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_257
timestamp 1666464484
transform 1 0 30128 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_261
timestamp 1666464484
transform 1 0 30576 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_265
timestamp 1666464484
transform 1 0 31024 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_272
timestamp 1666464484
transform 1 0 31808 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_276
timestamp 1666464484
transform 1 0 32256 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_284
timestamp 1666464484
transform 1 0 33152 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_288
timestamp 1666464484
transform 1 0 33600 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_290
timestamp 1666464484
transform 1 0 33824 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_293
timestamp 1666464484
transform 1 0 34160 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_301
timestamp 1666464484
transform 1 0 35056 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_318
timestamp 1666464484
transform 1 0 36960 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_321
timestamp 1666464484
transform 1 0 37296 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_328
timestamp 1666464484
transform 1 0 38080 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_18_332
timestamp 1666464484
transform 1 0 38528 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_364
timestamp 1666464484
transform 1 0 42112 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_380
timestamp 1666464484
transform 1 0 43904 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_388
timestamp 1666464484
transform 1 0 44800 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_392
timestamp 1666464484
transform 1 0 45248 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_408
timestamp 1666464484
transform 1 0 47040 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_416
timestamp 1666464484
transform 1 0 47936 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_2
timestamp 1666464484
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_66
timestamp 1666464484
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_70
timestamp 1666464484
transform 1 0 9184 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_73
timestamp 1666464484
transform 1 0 9520 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_137
timestamp 1666464484
transform 1 0 16688 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_141
timestamp 1666464484
transform 1 0 17136 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_144
timestamp 1666464484
transform 1 0 17472 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_208
timestamp 1666464484
transform 1 0 24640 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_212
timestamp 1666464484
transform 1 0 25088 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_19_215
timestamp 1666464484
transform 1 0 25424 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_253
timestamp 1666464484
transform 1 0 29680 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_257
timestamp 1666464484
transform 1 0 30128 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_261
timestamp 1666464484
transform 1 0 30576 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_269
timestamp 1666464484
transform 1 0 31472 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_277
timestamp 1666464484
transform 1 0 32368 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_281
timestamp 1666464484
transform 1 0 32816 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_283
timestamp 1666464484
transform 1 0 33040 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_286
timestamp 1666464484
transform 1 0 33376 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_294
timestamp 1666464484
transform 1 0 34272 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_298
timestamp 1666464484
transform 1 0 34720 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_301
timestamp 1666464484
transform 1 0 35056 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_309
timestamp 1666464484
transform 1 0 35952 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_326
timestamp 1666464484
transform 1 0 37856 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_330
timestamp 1666464484
transform 1 0 38304 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_334
timestamp 1666464484
transform 1 0 38752 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_350
timestamp 1666464484
transform 1 0 40544 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_354
timestamp 1666464484
transform 1 0 40992 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_19_357
timestamp 1666464484
transform 1 0 41328 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_389
timestamp 1666464484
transform 1 0 44912 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_397
timestamp 1666464484
transform 1 0 45808 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_403
timestamp 1666464484
transform 1 0 46480 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_419
timestamp 1666464484
transform 1 0 48272 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_2
timestamp 1666464484
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_34
timestamp 1666464484
transform 1 0 5152 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_37
timestamp 1666464484
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_101
timestamp 1666464484
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_105
timestamp 1666464484
transform 1 0 13104 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_108
timestamp 1666464484
transform 1 0 13440 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_172
timestamp 1666464484
transform 1 0 20608 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_176
timestamp 1666464484
transform 1 0 21056 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_179
timestamp 1666464484
transform 1 0 21392 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_243
timestamp 1666464484
transform 1 0 28560 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_247
timestamp 1666464484
transform 1 0 29008 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_250
timestamp 1666464484
transform 1 0 29344 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_258
timestamp 1666464484
transform 1 0 30240 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_262
timestamp 1666464484
transform 1 0 30688 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_269
timestamp 1666464484
transform 1 0 31472 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_285
timestamp 1666464484
transform 1 0 33264 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_287
timestamp 1666464484
transform 1 0 33488 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_290
timestamp 1666464484
transform 1 0 33824 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_297
timestamp 1666464484
transform 1 0 34608 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_301
timestamp 1666464484
transform 1 0 35056 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_305
timestamp 1666464484
transform 1 0 35504 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_309
timestamp 1666464484
transform 1 0 35952 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_313
timestamp 1666464484
transform 1 0 36400 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_315
timestamp 1666464484
transform 1 0 36624 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_318
timestamp 1666464484
transform 1 0 36960 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_321
timestamp 1666464484
transform 1 0 37296 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_337
timestamp 1666464484
transform 1 0 39088 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_369
timestamp 1666464484
transform 1 0 42672 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_385
timestamp 1666464484
transform 1 0 44464 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_389
timestamp 1666464484
transform 1 0 44912 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_392
timestamp 1666464484
transform 1 0 45248 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_400
timestamp 1666464484
transform 1 0 46144 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_403
timestamp 1666464484
transform 1 0 46480 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_419
timestamp 1666464484
transform 1 0 48272 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_2
timestamp 1666464484
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_66
timestamp 1666464484
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_70
timestamp 1666464484
transform 1 0 9184 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_73
timestamp 1666464484
transform 1 0 9520 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_137
timestamp 1666464484
transform 1 0 16688 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_141
timestamp 1666464484
transform 1 0 17136 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_144
timestamp 1666464484
transform 1 0 17472 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_208
timestamp 1666464484
transform 1 0 24640 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_212
timestamp 1666464484
transform 1 0 25088 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_21_215
timestamp 1666464484
transform 1 0 25424 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_247
timestamp 1666464484
transform 1 0 29008 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_249
timestamp 1666464484
transform 1 0 29232 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_252
timestamp 1666464484
transform 1 0 29568 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_268
timestamp 1666464484
transform 1 0 31360 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_272
timestamp 1666464484
transform 1 0 31808 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_274
timestamp 1666464484
transform 1 0 32032 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_281
timestamp 1666464484
transform 1 0 32816 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_283
timestamp 1666464484
transform 1 0 33040 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_286
timestamp 1666464484
transform 1 0 33376 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_293
timestamp 1666464484
transform 1 0 34160 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_301
timestamp 1666464484
transform 1 0 35056 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_311
timestamp 1666464484
transform 1 0 36176 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_315
timestamp 1666464484
transform 1 0 36624 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_332
timestamp 1666464484
transform 1 0 38528 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_336
timestamp 1666464484
transform 1 0 38976 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_339
timestamp 1666464484
transform 1 0 39312 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_21_357
timestamp 1666464484
transform 1 0 41328 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_389
timestamp 1666464484
transform 1 0 44912 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_405
timestamp 1666464484
transform 1 0 46704 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_413
timestamp 1666464484
transform 1 0 47600 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_417
timestamp 1666464484
transform 1 0 48048 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_419
timestamp 1666464484
transform 1 0 48272 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_2
timestamp 1666464484
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_34
timestamp 1666464484
transform 1 0 5152 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_37
timestamp 1666464484
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_101
timestamp 1666464484
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_105
timestamp 1666464484
transform 1 0 13104 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_108
timestamp 1666464484
transform 1 0 13440 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_172
timestamp 1666464484
transform 1 0 20608 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_176
timestamp 1666464484
transform 1 0 21056 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_179
timestamp 1666464484
transform 1 0 21392 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_243
timestamp 1666464484
transform 1 0 28560 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_247
timestamp 1666464484
transform 1 0 29008 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_250
timestamp 1666464484
transform 1 0 29344 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_267
timestamp 1666464484
transform 1 0 31248 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_271
timestamp 1666464484
transform 1 0 31696 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_279
timestamp 1666464484
transform 1 0 32592 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_289
timestamp 1666464484
transform 1 0 33712 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_305
timestamp 1666464484
transform 1 0 35504 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_309
timestamp 1666464484
transform 1 0 35952 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_311
timestamp 1666464484
transform 1 0 36176 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_314
timestamp 1666464484
transform 1 0 36512 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_318
timestamp 1666464484
transform 1 0 36960 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_321
timestamp 1666464484
transform 1 0 37296 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_337
timestamp 1666464484
transform 1 0 39088 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_346
timestamp 1666464484
transform 1 0 40096 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_354
timestamp 1666464484
transform 1 0 40992 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_386
timestamp 1666464484
transform 1 0 44576 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_392
timestamp 1666464484
transform 1 0 45248 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_400
timestamp 1666464484
transform 1 0 46144 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_403
timestamp 1666464484
transform 1 0 46480 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_419
timestamp 1666464484
transform 1 0 48272 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_2
timestamp 1666464484
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_66
timestamp 1666464484
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_70
timestamp 1666464484
transform 1 0 9184 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_73
timestamp 1666464484
transform 1 0 9520 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_137
timestamp 1666464484
transform 1 0 16688 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_141
timestamp 1666464484
transform 1 0 17136 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_144
timestamp 1666464484
transform 1 0 17472 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_208
timestamp 1666464484
transform 1 0 24640 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_212
timestamp 1666464484
transform 1 0 25088 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_215
timestamp 1666464484
transform 1 0 25424 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_279
timestamp 1666464484
transform 1 0 32592 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_283
timestamp 1666464484
transform 1 0 33040 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_286
timestamp 1666464484
transform 1 0 33376 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_302
timestamp 1666464484
transform 1 0 35168 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_310
timestamp 1666464484
transform 1 0 36064 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_312
timestamp 1666464484
transform 1 0 36288 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_315
timestamp 1666464484
transform 1 0 36624 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_319
timestamp 1666464484
transform 1 0 37072 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_336
timestamp 1666464484
transform 1 0 38976 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_352
timestamp 1666464484
transform 1 0 40768 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_354
timestamp 1666464484
transform 1 0 40992 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_23_357
timestamp 1666464484
transform 1 0 41328 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_389
timestamp 1666464484
transform 1 0 44912 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_405
timestamp 1666464484
transform 1 0 46704 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_413
timestamp 1666464484
transform 1 0 47600 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_417
timestamp 1666464484
transform 1 0 48048 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_419
timestamp 1666464484
transform 1 0 48272 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_2
timestamp 1666464484
transform 1 0 1568 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_7
timestamp 1666464484
transform 1 0 2128 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_23
timestamp 1666464484
transform 1 0 3920 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_31
timestamp 1666464484
transform 1 0 4816 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_37
timestamp 1666464484
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_101
timestamp 1666464484
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_105
timestamp 1666464484
transform 1 0 13104 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_108
timestamp 1666464484
transform 1 0 13440 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_172
timestamp 1666464484
transform 1 0 20608 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_176
timestamp 1666464484
transform 1 0 21056 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_179
timestamp 1666464484
transform 1 0 21392 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_211
timestamp 1666464484
transform 1 0 24976 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_227
timestamp 1666464484
transform 1 0 26768 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_235
timestamp 1666464484
transform 1 0 27664 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_243
timestamp 1666464484
transform 1 0 28560 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_247
timestamp 1666464484
transform 1 0 29008 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_250
timestamp 1666464484
transform 1 0 29344 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_314
timestamp 1666464484
transform 1 0 36512 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_318
timestamp 1666464484
transform 1 0 36960 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_321
timestamp 1666464484
transform 1 0 37296 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_325
timestamp 1666464484
transform 1 0 37744 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_331
timestamp 1666464484
transform 1 0 38416 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_335
timestamp 1666464484
transform 1 0 38864 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_367
timestamp 1666464484
transform 1 0 42448 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_383
timestamp 1666464484
transform 1 0 44240 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_387
timestamp 1666464484
transform 1 0 44688 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_389
timestamp 1666464484
transform 1 0 44912 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_392
timestamp 1666464484
transform 1 0 45248 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_400
timestamp 1666464484
transform 1 0 46144 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_403
timestamp 1666464484
transform 1 0 46480 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_419
timestamp 1666464484
transform 1 0 48272 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_2
timestamp 1666464484
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_66
timestamp 1666464484
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_70
timestamp 1666464484
transform 1 0 9184 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_73
timestamp 1666464484
transform 1 0 9520 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_137
timestamp 1666464484
transform 1 0 16688 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_141
timestamp 1666464484
transform 1 0 17136 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_144
timestamp 1666464484
transform 1 0 17472 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_208
timestamp 1666464484
transform 1 0 24640 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_212
timestamp 1666464484
transform 1 0 25088 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_215
timestamp 1666464484
transform 1 0 25424 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_279
timestamp 1666464484
transform 1 0 32592 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_283
timestamp 1666464484
transform 1 0 33040 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_286
timestamp 1666464484
transform 1 0 33376 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_302
timestamp 1666464484
transform 1 0 35168 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_310
timestamp 1666464484
transform 1 0 36064 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_314
timestamp 1666464484
transform 1 0 36512 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_316
timestamp 1666464484
transform 1 0 36736 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_319
timestamp 1666464484
transform 1 0 37072 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_323
timestamp 1666464484
transform 1 0 37520 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_340
timestamp 1666464484
transform 1 0 39424 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_348
timestamp 1666464484
transform 1 0 40320 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_352
timestamp 1666464484
transform 1 0 40768 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_354
timestamp 1666464484
transform 1 0 40992 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_25_357
timestamp 1666464484
transform 1 0 41328 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_389
timestamp 1666464484
transform 1 0 44912 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_405
timestamp 1666464484
transform 1 0 46704 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_413
timestamp 1666464484
transform 1 0 47600 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_417
timestamp 1666464484
transform 1 0 48048 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_419
timestamp 1666464484
transform 1 0 48272 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_2
timestamp 1666464484
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_34
timestamp 1666464484
transform 1 0 5152 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_37
timestamp 1666464484
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_101
timestamp 1666464484
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_105
timestamp 1666464484
transform 1 0 13104 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_108
timestamp 1666464484
transform 1 0 13440 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_172
timestamp 1666464484
transform 1 0 20608 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_176
timestamp 1666464484
transform 1 0 21056 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_179
timestamp 1666464484
transform 1 0 21392 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_243
timestamp 1666464484
transform 1 0 28560 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_247
timestamp 1666464484
transform 1 0 29008 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_250
timestamp 1666464484
transform 1 0 29344 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_314
timestamp 1666464484
transform 1 0 36512 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_318
timestamp 1666464484
transform 1 0 36960 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_321
timestamp 1666464484
transform 1 0 37296 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_340
timestamp 1666464484
transform 1 0 39424 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_344
timestamp 1666464484
transform 1 0 39872 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_346
timestamp 1666464484
transform 1 0 40096 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_355
timestamp 1666464484
transform 1 0 41104 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_387
timestamp 1666464484
transform 1 0 44688 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_389
timestamp 1666464484
transform 1 0 44912 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_392
timestamp 1666464484
transform 1 0 45248 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_400
timestamp 1666464484
transform 1 0 46144 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_403
timestamp 1666464484
transform 1 0 46480 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_419
timestamp 1666464484
transform 1 0 48272 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_2
timestamp 1666464484
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_66
timestamp 1666464484
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_70
timestamp 1666464484
transform 1 0 9184 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_73
timestamp 1666464484
transform 1 0 9520 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_137
timestamp 1666464484
transform 1 0 16688 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_141
timestamp 1666464484
transform 1 0 17136 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_144
timestamp 1666464484
transform 1 0 17472 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_208
timestamp 1666464484
transform 1 0 24640 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_212
timestamp 1666464484
transform 1 0 25088 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_215
timestamp 1666464484
transform 1 0 25424 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_279
timestamp 1666464484
transform 1 0 32592 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_283
timestamp 1666464484
transform 1 0 33040 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_27_286
timestamp 1666464484
transform 1 0 33376 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_320
timestamp 1666464484
transform 1 0 37184 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_324
timestamp 1666464484
transform 1 0 37632 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_341
timestamp 1666464484
transform 1 0 39536 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_349
timestamp 1666464484
transform 1 0 40432 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_353
timestamp 1666464484
transform 1 0 40880 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_27_357
timestamp 1666464484
transform 1 0 41328 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_389
timestamp 1666464484
transform 1 0 44912 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_405
timestamp 1666464484
transform 1 0 46704 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_413
timestamp 1666464484
transform 1 0 47600 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_417
timestamp 1666464484
transform 1 0 48048 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_419
timestamp 1666464484
transform 1 0 48272 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_2
timestamp 1666464484
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_34
timestamp 1666464484
transform 1 0 5152 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_37
timestamp 1666464484
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_101
timestamp 1666464484
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_105
timestamp 1666464484
transform 1 0 13104 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_108
timestamp 1666464484
transform 1 0 13440 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_172
timestamp 1666464484
transform 1 0 20608 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_176
timestamp 1666464484
transform 1 0 21056 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_179
timestamp 1666464484
transform 1 0 21392 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_243
timestamp 1666464484
transform 1 0 28560 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_247
timestamp 1666464484
transform 1 0 29008 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_250
timestamp 1666464484
transform 1 0 29344 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_314
timestamp 1666464484
transform 1 0 36512 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_318
timestamp 1666464484
transform 1 0 36960 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_321
timestamp 1666464484
transform 1 0 37296 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_337
timestamp 1666464484
transform 1 0 39088 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_345
timestamp 1666464484
transform 1 0 39984 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_354
timestamp 1666464484
transform 1 0 40992 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_386
timestamp 1666464484
transform 1 0 44576 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_392
timestamp 1666464484
transform 1 0 45248 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_400
timestamp 1666464484
transform 1 0 46144 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_403
timestamp 1666464484
transform 1 0 46480 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_419
timestamp 1666464484
transform 1 0 48272 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_2
timestamp 1666464484
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_66
timestamp 1666464484
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_70
timestamp 1666464484
transform 1 0 9184 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_73
timestamp 1666464484
transform 1 0 9520 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_137
timestamp 1666464484
transform 1 0 16688 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_141
timestamp 1666464484
transform 1 0 17136 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_144
timestamp 1666464484
transform 1 0 17472 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_208
timestamp 1666464484
transform 1 0 24640 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_212
timestamp 1666464484
transform 1 0 25088 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_215
timestamp 1666464484
transform 1 0 25424 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_279
timestamp 1666464484
transform 1 0 32592 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_283
timestamp 1666464484
transform 1 0 33040 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_29_286
timestamp 1666464484
transform 1 0 33376 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_318
timestamp 1666464484
transform 1 0 36960 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_321
timestamp 1666464484
transform 1 0 37296 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_325
timestamp 1666464484
transform 1 0 37744 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_342
timestamp 1666464484
transform 1 0 39648 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_350
timestamp 1666464484
transform 1 0 40544 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_354
timestamp 1666464484
transform 1 0 40992 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_29_357
timestamp 1666464484
transform 1 0 41328 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_389
timestamp 1666464484
transform 1 0 44912 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_405
timestamp 1666464484
transform 1 0 46704 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_413
timestamp 1666464484
transform 1 0 47600 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_417
timestamp 1666464484
transform 1 0 48048 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_419
timestamp 1666464484
transform 1 0 48272 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_2
timestamp 1666464484
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_34
timestamp 1666464484
transform 1 0 5152 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_37
timestamp 1666464484
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_101
timestamp 1666464484
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_105
timestamp 1666464484
transform 1 0 13104 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_108
timestamp 1666464484
transform 1 0 13440 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_172
timestamp 1666464484
transform 1 0 20608 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_176
timestamp 1666464484
transform 1 0 21056 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_179
timestamp 1666464484
transform 1 0 21392 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_243
timestamp 1666464484
transform 1 0 28560 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_247
timestamp 1666464484
transform 1 0 29008 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_250
timestamp 1666464484
transform 1 0 29344 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_314
timestamp 1666464484
transform 1 0 36512 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_318
timestamp 1666464484
transform 1 0 36960 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_321
timestamp 1666464484
transform 1 0 37296 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_329
timestamp 1666464484
transform 1 0 38192 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_333
timestamp 1666464484
transform 1 0 38640 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_336
timestamp 1666464484
transform 1 0 38976 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_340
timestamp 1666464484
transform 1 0 39424 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_349
timestamp 1666464484
transform 1 0 40432 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_381
timestamp 1666464484
transform 1 0 44016 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_389
timestamp 1666464484
transform 1 0 44912 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_392
timestamp 1666464484
transform 1 0 45248 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_400
timestamp 1666464484
transform 1 0 46144 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_403
timestamp 1666464484
transform 1 0 46480 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_419
timestamp 1666464484
transform 1 0 48272 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_2
timestamp 1666464484
transform 1 0 1568 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_5
timestamp 1666464484
transform 1 0 1904 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_69
timestamp 1666464484
transform 1 0 9072 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_73
timestamp 1666464484
transform 1 0 9520 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_137
timestamp 1666464484
transform 1 0 16688 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_141
timestamp 1666464484
transform 1 0 17136 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_144
timestamp 1666464484
transform 1 0 17472 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_208
timestamp 1666464484
transform 1 0 24640 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_212
timestamp 1666464484
transform 1 0 25088 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_215
timestamp 1666464484
transform 1 0 25424 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_279
timestamp 1666464484
transform 1 0 32592 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_283
timestamp 1666464484
transform 1 0 33040 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_286
timestamp 1666464484
transform 1 0 33376 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_302
timestamp 1666464484
transform 1 0 35168 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_310
timestamp 1666464484
transform 1 0 36064 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_313
timestamp 1666464484
transform 1 0 36400 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_317
timestamp 1666464484
transform 1 0 36848 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_334
timestamp 1666464484
transform 1 0 38752 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_344
timestamp 1666464484
transform 1 0 39872 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_352
timestamp 1666464484
transform 1 0 40768 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_354
timestamp 1666464484
transform 1 0 40992 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_31_357
timestamp 1666464484
transform 1 0 41328 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_389
timestamp 1666464484
transform 1 0 44912 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_405
timestamp 1666464484
transform 1 0 46704 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_413
timestamp 1666464484
transform 1 0 47600 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_417
timestamp 1666464484
transform 1 0 48048 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_419
timestamp 1666464484
transform 1 0 48272 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_2
timestamp 1666464484
transform 1 0 1568 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_9
timestamp 1666464484
transform 1 0 2352 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_25
timestamp 1666464484
transform 1 0 4144 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_33
timestamp 1666464484
transform 1 0 5040 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_37
timestamp 1666464484
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_101
timestamp 1666464484
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_105
timestamp 1666464484
transform 1 0 13104 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_108
timestamp 1666464484
transform 1 0 13440 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_172
timestamp 1666464484
transform 1 0 20608 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_176
timestamp 1666464484
transform 1 0 21056 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_179
timestamp 1666464484
transform 1 0 21392 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_243
timestamp 1666464484
transform 1 0 28560 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_247
timestamp 1666464484
transform 1 0 29008 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_250
timestamp 1666464484
transform 1 0 29344 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_314
timestamp 1666464484
transform 1 0 36512 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_318
timestamp 1666464484
transform 1 0 36960 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_321
timestamp 1666464484
transform 1 0 37296 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_340
timestamp 1666464484
transform 1 0 39424 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_344
timestamp 1666464484
transform 1 0 39872 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_348
timestamp 1666464484
transform 1 0 40320 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_380
timestamp 1666464484
transform 1 0 43904 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_388
timestamp 1666464484
transform 1 0 44800 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_392
timestamp 1666464484
transform 1 0 45248 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_400
timestamp 1666464484
transform 1 0 46144 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_403
timestamp 1666464484
transform 1 0 46480 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_419
timestamp 1666464484
transform 1 0 48272 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_2
timestamp 1666464484
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_66
timestamp 1666464484
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_70
timestamp 1666464484
transform 1 0 9184 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_73
timestamp 1666464484
transform 1 0 9520 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_137
timestamp 1666464484
transform 1 0 16688 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_141
timestamp 1666464484
transform 1 0 17136 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_144
timestamp 1666464484
transform 1 0 17472 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_208
timestamp 1666464484
transform 1 0 24640 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_212
timestamp 1666464484
transform 1 0 25088 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_215
timestamp 1666464484
transform 1 0 25424 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_279
timestamp 1666464484
transform 1 0 32592 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_283
timestamp 1666464484
transform 1 0 33040 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_286
timestamp 1666464484
transform 1 0 33376 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_302
timestamp 1666464484
transform 1 0 35168 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_310
timestamp 1666464484
transform 1 0 36064 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_314
timestamp 1666464484
transform 1 0 36512 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_316
timestamp 1666464484
transform 1 0 36736 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_319
timestamp 1666464484
transform 1 0 37072 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_323
timestamp 1666464484
transform 1 0 37520 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_340
timestamp 1666464484
transform 1 0 39424 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_344
timestamp 1666464484
transform 1 0 39872 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_352
timestamp 1666464484
transform 1 0 40768 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_354
timestamp 1666464484
transform 1 0 40992 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_33_357
timestamp 1666464484
transform 1 0 41328 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_389
timestamp 1666464484
transform 1 0 44912 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_397
timestamp 1666464484
transform 1 0 45808 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_403
timestamp 1666464484
transform 1 0 46480 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_419
timestamp 1666464484
transform 1 0 48272 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_2
timestamp 1666464484
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_34
timestamp 1666464484
transform 1 0 5152 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_37
timestamp 1666464484
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_101
timestamp 1666464484
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_105
timestamp 1666464484
transform 1 0 13104 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_108
timestamp 1666464484
transform 1 0 13440 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_172
timestamp 1666464484
transform 1 0 20608 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_176
timestamp 1666464484
transform 1 0 21056 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_179
timestamp 1666464484
transform 1 0 21392 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_243
timestamp 1666464484
transform 1 0 28560 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_247
timestamp 1666464484
transform 1 0 29008 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_250
timestamp 1666464484
transform 1 0 29344 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_314
timestamp 1666464484
transform 1 0 36512 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_318
timestamp 1666464484
transform 1 0 36960 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_321
timestamp 1666464484
transform 1 0 37296 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_385
timestamp 1666464484
transform 1 0 44464 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_389
timestamp 1666464484
transform 1 0 44912 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_392
timestamp 1666464484
transform 1 0 45248 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_408
timestamp 1666464484
transform 1 0 47040 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_416
timestamp 1666464484
transform 1 0 47936 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_2
timestamp 1666464484
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_66
timestamp 1666464484
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_70
timestamp 1666464484
transform 1 0 9184 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_73
timestamp 1666464484
transform 1 0 9520 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_137
timestamp 1666464484
transform 1 0 16688 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_141
timestamp 1666464484
transform 1 0 17136 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_144
timestamp 1666464484
transform 1 0 17472 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_208
timestamp 1666464484
transform 1 0 24640 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_212
timestamp 1666464484
transform 1 0 25088 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_215
timestamp 1666464484
transform 1 0 25424 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_279
timestamp 1666464484
transform 1 0 32592 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_283
timestamp 1666464484
transform 1 0 33040 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_286
timestamp 1666464484
transform 1 0 33376 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_350
timestamp 1666464484
transform 1 0 40544 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_354
timestamp 1666464484
transform 1 0 40992 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_35_357
timestamp 1666464484
transform 1 0 41328 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_389
timestamp 1666464484
transform 1 0 44912 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_397
timestamp 1666464484
transform 1 0 45808 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_403
timestamp 1666464484
transform 1 0 46480 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_419
timestamp 1666464484
transform 1 0 48272 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_2
timestamp 1666464484
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_34
timestamp 1666464484
transform 1 0 5152 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_37
timestamp 1666464484
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_101
timestamp 1666464484
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_105
timestamp 1666464484
transform 1 0 13104 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_108
timestamp 1666464484
transform 1 0 13440 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_172
timestamp 1666464484
transform 1 0 20608 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_176
timestamp 1666464484
transform 1 0 21056 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_179
timestamp 1666464484
transform 1 0 21392 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_243
timestamp 1666464484
transform 1 0 28560 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_247
timestamp 1666464484
transform 1 0 29008 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_250
timestamp 1666464484
transform 1 0 29344 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_314
timestamp 1666464484
transform 1 0 36512 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_318
timestamp 1666464484
transform 1 0 36960 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_321
timestamp 1666464484
transform 1 0 37296 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_385
timestamp 1666464484
transform 1 0 44464 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_389
timestamp 1666464484
transform 1 0 44912 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_392
timestamp 1666464484
transform 1 0 45248 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_408
timestamp 1666464484
transform 1 0 47040 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_416
timestamp 1666464484
transform 1 0 47936 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_2
timestamp 1666464484
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_66
timestamp 1666464484
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_70
timestamp 1666464484
transform 1 0 9184 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_73
timestamp 1666464484
transform 1 0 9520 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_137
timestamp 1666464484
transform 1 0 16688 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_141
timestamp 1666464484
transform 1 0 17136 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_144
timestamp 1666464484
transform 1 0 17472 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_208
timestamp 1666464484
transform 1 0 24640 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_212
timestamp 1666464484
transform 1 0 25088 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_215
timestamp 1666464484
transform 1 0 25424 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_279
timestamp 1666464484
transform 1 0 32592 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_283
timestamp 1666464484
transform 1 0 33040 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_286
timestamp 1666464484
transform 1 0 33376 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_350
timestamp 1666464484
transform 1 0 40544 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_354
timestamp 1666464484
transform 1 0 40992 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_357
timestamp 1666464484
transform 1 0 41328 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_389
timestamp 1666464484
transform 1 0 44912 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_397
timestamp 1666464484
transform 1 0 45808 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_403
timestamp 1666464484
transform 1 0 46480 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_419
timestamp 1666464484
transform 1 0 48272 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_2
timestamp 1666464484
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_34
timestamp 1666464484
transform 1 0 5152 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_37
timestamp 1666464484
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_101
timestamp 1666464484
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_105
timestamp 1666464484
transform 1 0 13104 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_108
timestamp 1666464484
transform 1 0 13440 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_172
timestamp 1666464484
transform 1 0 20608 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_176
timestamp 1666464484
transform 1 0 21056 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_179
timestamp 1666464484
transform 1 0 21392 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_243
timestamp 1666464484
transform 1 0 28560 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_247
timestamp 1666464484
transform 1 0 29008 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_250
timestamp 1666464484
transform 1 0 29344 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_314
timestamp 1666464484
transform 1 0 36512 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_318
timestamp 1666464484
transform 1 0 36960 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_321
timestamp 1666464484
transform 1 0 37296 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_385
timestamp 1666464484
transform 1 0 44464 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_389
timestamp 1666464484
transform 1 0 44912 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_392
timestamp 1666464484
transform 1 0 45248 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_408
timestamp 1666464484
transform 1 0 47040 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_416
timestamp 1666464484
transform 1 0 47936 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_2
timestamp 1666464484
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_66
timestamp 1666464484
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_70
timestamp 1666464484
transform 1 0 9184 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_73
timestamp 1666464484
transform 1 0 9520 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_137
timestamp 1666464484
transform 1 0 16688 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_141
timestamp 1666464484
transform 1 0 17136 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_144
timestamp 1666464484
transform 1 0 17472 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_208
timestamp 1666464484
transform 1 0 24640 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_212
timestamp 1666464484
transform 1 0 25088 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_215
timestamp 1666464484
transform 1 0 25424 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_279
timestamp 1666464484
transform 1 0 32592 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_283
timestamp 1666464484
transform 1 0 33040 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_286
timestamp 1666464484
transform 1 0 33376 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_350
timestamp 1666464484
transform 1 0 40544 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_354
timestamp 1666464484
transform 1 0 40992 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_39_357
timestamp 1666464484
transform 1 0 41328 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_389
timestamp 1666464484
transform 1 0 44912 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_397
timestamp 1666464484
transform 1 0 45808 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_403
timestamp 1666464484
transform 1 0 46480 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_419
timestamp 1666464484
transform 1 0 48272 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_2
timestamp 1666464484
transform 1 0 1568 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_7
timestamp 1666464484
transform 1 0 2128 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_23
timestamp 1666464484
transform 1 0 3920 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_31
timestamp 1666464484
transform 1 0 4816 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_37
timestamp 1666464484
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_101
timestamp 1666464484
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_105
timestamp 1666464484
transform 1 0 13104 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_108
timestamp 1666464484
transform 1 0 13440 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_172
timestamp 1666464484
transform 1 0 20608 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_176
timestamp 1666464484
transform 1 0 21056 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_179
timestamp 1666464484
transform 1 0 21392 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_243
timestamp 1666464484
transform 1 0 28560 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_247
timestamp 1666464484
transform 1 0 29008 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_250
timestamp 1666464484
transform 1 0 29344 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_314
timestamp 1666464484
transform 1 0 36512 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_318
timestamp 1666464484
transform 1 0 36960 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_321
timestamp 1666464484
transform 1 0 37296 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_385
timestamp 1666464484
transform 1 0 44464 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_389
timestamp 1666464484
transform 1 0 44912 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_392
timestamp 1666464484
transform 1 0 45248 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_408
timestamp 1666464484
transform 1 0 47040 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_416
timestamp 1666464484
transform 1 0 47936 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_2
timestamp 1666464484
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_66
timestamp 1666464484
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_70
timestamp 1666464484
transform 1 0 9184 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_73
timestamp 1666464484
transform 1 0 9520 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_137
timestamp 1666464484
transform 1 0 16688 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_141
timestamp 1666464484
transform 1 0 17136 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_144
timestamp 1666464484
transform 1 0 17472 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_208
timestamp 1666464484
transform 1 0 24640 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_212
timestamp 1666464484
transform 1 0 25088 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_215
timestamp 1666464484
transform 1 0 25424 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_279
timestamp 1666464484
transform 1 0 32592 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_283
timestamp 1666464484
transform 1 0 33040 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_286
timestamp 1666464484
transform 1 0 33376 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_350
timestamp 1666464484
transform 1 0 40544 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_354
timestamp 1666464484
transform 1 0 40992 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_41_357
timestamp 1666464484
transform 1 0 41328 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_389
timestamp 1666464484
transform 1 0 44912 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_397
timestamp 1666464484
transform 1 0 45808 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_403
timestamp 1666464484
transform 1 0 46480 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_419
timestamp 1666464484
transform 1 0 48272 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_2
timestamp 1666464484
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_34
timestamp 1666464484
transform 1 0 5152 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_37
timestamp 1666464484
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_101
timestamp 1666464484
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_105
timestamp 1666464484
transform 1 0 13104 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_108
timestamp 1666464484
transform 1 0 13440 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_140
timestamp 1666464484
transform 1 0 17024 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_142
timestamp 1666464484
transform 1 0 17248 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_145
timestamp 1666464484
transform 1 0 17584 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_153
timestamp 1666464484
transform 1 0 18480 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_169
timestamp 1666464484
transform 1 0 20272 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_179
timestamp 1666464484
transform 1 0 21392 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_243
timestamp 1666464484
transform 1 0 28560 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_247
timestamp 1666464484
transform 1 0 29008 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_250
timestamp 1666464484
transform 1 0 29344 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_314
timestamp 1666464484
transform 1 0 36512 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_318
timestamp 1666464484
transform 1 0 36960 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_321
timestamp 1666464484
transform 1 0 37296 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_385
timestamp 1666464484
transform 1 0 44464 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_389
timestamp 1666464484
transform 1 0 44912 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_392
timestamp 1666464484
transform 1 0 45248 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_408
timestamp 1666464484
transform 1 0 47040 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_416
timestamp 1666464484
transform 1 0 47936 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_2
timestamp 1666464484
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_66
timestamp 1666464484
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_70
timestamp 1666464484
transform 1 0 9184 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_73
timestamp 1666464484
transform 1 0 9520 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_137
timestamp 1666464484
transform 1 0 16688 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_141
timestamp 1666464484
transform 1 0 17136 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_144
timestamp 1666464484
transform 1 0 17472 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_208
timestamp 1666464484
transform 1 0 24640 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_212
timestamp 1666464484
transform 1 0 25088 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_215
timestamp 1666464484
transform 1 0 25424 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_279
timestamp 1666464484
transform 1 0 32592 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_283
timestamp 1666464484
transform 1 0 33040 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_286
timestamp 1666464484
transform 1 0 33376 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_350
timestamp 1666464484
transform 1 0 40544 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_354
timestamp 1666464484
transform 1 0 40992 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_43_357
timestamp 1666464484
transform 1 0 41328 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_389
timestamp 1666464484
transform 1 0 44912 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_397
timestamp 1666464484
transform 1 0 45808 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_403
timestamp 1666464484
transform 1 0 46480 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_419
timestamp 1666464484
transform 1 0 48272 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_44_2
timestamp 1666464484
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_34
timestamp 1666464484
transform 1 0 5152 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_37
timestamp 1666464484
transform 1 0 5488 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_101
timestamp 1666464484
transform 1 0 12656 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_105
timestamp 1666464484
transform 1 0 13104 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_108
timestamp 1666464484
transform 1 0 13440 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_172
timestamp 1666464484
transform 1 0 20608 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_176
timestamp 1666464484
transform 1 0 21056 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_179
timestamp 1666464484
transform 1 0 21392 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_243
timestamp 1666464484
transform 1 0 28560 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_247
timestamp 1666464484
transform 1 0 29008 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_250
timestamp 1666464484
transform 1 0 29344 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_314
timestamp 1666464484
transform 1 0 36512 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_318
timestamp 1666464484
transform 1 0 36960 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_321
timestamp 1666464484
transform 1 0 37296 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_385
timestamp 1666464484
transform 1 0 44464 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_389
timestamp 1666464484
transform 1 0 44912 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_392
timestamp 1666464484
transform 1 0 45248 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_408
timestamp 1666464484
transform 1 0 47040 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_416
timestamp 1666464484
transform 1 0 47936 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_2
timestamp 1666464484
transform 1 0 1568 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_66
timestamp 1666464484
transform 1 0 8736 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_70
timestamp 1666464484
transform 1 0 9184 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_73
timestamp 1666464484
transform 1 0 9520 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_137
timestamp 1666464484
transform 1 0 16688 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_141
timestamp 1666464484
transform 1 0 17136 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_144
timestamp 1666464484
transform 1 0 17472 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_208
timestamp 1666464484
transform 1 0 24640 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_212
timestamp 1666464484
transform 1 0 25088 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_215
timestamp 1666464484
transform 1 0 25424 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_279
timestamp 1666464484
transform 1 0 32592 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_283
timestamp 1666464484
transform 1 0 33040 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_286
timestamp 1666464484
transform 1 0 33376 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_350
timestamp 1666464484
transform 1 0 40544 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_354
timestamp 1666464484
transform 1 0 40992 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_45_357
timestamp 1666464484
transform 1 0 41328 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_389
timestamp 1666464484
transform 1 0 44912 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_397
timestamp 1666464484
transform 1 0 45808 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_403
timestamp 1666464484
transform 1 0 46480 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_419
timestamp 1666464484
transform 1 0 48272 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_46_2
timestamp 1666464484
transform 1 0 1568 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_34
timestamp 1666464484
transform 1 0 5152 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_37
timestamp 1666464484
transform 1 0 5488 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_101
timestamp 1666464484
transform 1 0 12656 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_105
timestamp 1666464484
transform 1 0 13104 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_108
timestamp 1666464484
transform 1 0 13440 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_172
timestamp 1666464484
transform 1 0 20608 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_176
timestamp 1666464484
transform 1 0 21056 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_179
timestamp 1666464484
transform 1 0 21392 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_243
timestamp 1666464484
transform 1 0 28560 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_247
timestamp 1666464484
transform 1 0 29008 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_250
timestamp 1666464484
transform 1 0 29344 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_314
timestamp 1666464484
transform 1 0 36512 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_318
timestamp 1666464484
transform 1 0 36960 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_321
timestamp 1666464484
transform 1 0 37296 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_385
timestamp 1666464484
transform 1 0 44464 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_389
timestamp 1666464484
transform 1 0 44912 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_392
timestamp 1666464484
transform 1 0 45248 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_400
timestamp 1666464484
transform 1 0 46144 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_403
timestamp 1666464484
transform 1 0 46480 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_419
timestamp 1666464484
transform 1 0 48272 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_2
timestamp 1666464484
transform 1 0 1568 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_66
timestamp 1666464484
transform 1 0 8736 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_70
timestamp 1666464484
transform 1 0 9184 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_73
timestamp 1666464484
transform 1 0 9520 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_137
timestamp 1666464484
transform 1 0 16688 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_141
timestamp 1666464484
transform 1 0 17136 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_144
timestamp 1666464484
transform 1 0 17472 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_208
timestamp 1666464484
transform 1 0 24640 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_212
timestamp 1666464484
transform 1 0 25088 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_215
timestamp 1666464484
transform 1 0 25424 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_279
timestamp 1666464484
transform 1 0 32592 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_283
timestamp 1666464484
transform 1 0 33040 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_286
timestamp 1666464484
transform 1 0 33376 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_350
timestamp 1666464484
transform 1 0 40544 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_354
timestamp 1666464484
transform 1 0 40992 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_357
timestamp 1666464484
transform 1 0 41328 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_389
timestamp 1666464484
transform 1 0 44912 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_405
timestamp 1666464484
transform 1 0 46704 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_413
timestamp 1666464484
transform 1 0 47600 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_417
timestamp 1666464484
transform 1 0 48048 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_419
timestamp 1666464484
transform 1 0 48272 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_2
timestamp 1666464484
transform 1 0 1568 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_17
timestamp 1666464484
transform 1 0 3248 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_21
timestamp 1666464484
transform 1 0 3696 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_29
timestamp 1666464484
transform 1 0 4592 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_33
timestamp 1666464484
transform 1 0 5040 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_37
timestamp 1666464484
transform 1 0 5488 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_101
timestamp 1666464484
transform 1 0 12656 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_105
timestamp 1666464484
transform 1 0 13104 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_108
timestamp 1666464484
transform 1 0 13440 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_172
timestamp 1666464484
transform 1 0 20608 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_176
timestamp 1666464484
transform 1 0 21056 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_179
timestamp 1666464484
transform 1 0 21392 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_243
timestamp 1666464484
transform 1 0 28560 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_247
timestamp 1666464484
transform 1 0 29008 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_250
timestamp 1666464484
transform 1 0 29344 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_314
timestamp 1666464484
transform 1 0 36512 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_318
timestamp 1666464484
transform 1 0 36960 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_321
timestamp 1666464484
transform 1 0 37296 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_385
timestamp 1666464484
transform 1 0 44464 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_389
timestamp 1666464484
transform 1 0 44912 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_392
timestamp 1666464484
transform 1 0 45248 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_400
timestamp 1666464484
transform 1 0 46144 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_403
timestamp 1666464484
transform 1 0 46480 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_419
timestamp 1666464484
transform 1 0 48272 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_2
timestamp 1666464484
transform 1 0 1568 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_66
timestamp 1666464484
transform 1 0 8736 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_70
timestamp 1666464484
transform 1 0 9184 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_73
timestamp 1666464484
transform 1 0 9520 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_137
timestamp 1666464484
transform 1 0 16688 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_141
timestamp 1666464484
transform 1 0 17136 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_144
timestamp 1666464484
transform 1 0 17472 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_208
timestamp 1666464484
transform 1 0 24640 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_212
timestamp 1666464484
transform 1 0 25088 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_215
timestamp 1666464484
transform 1 0 25424 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_279
timestamp 1666464484
transform 1 0 32592 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_283
timestamp 1666464484
transform 1 0 33040 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_286
timestamp 1666464484
transform 1 0 33376 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_350
timestamp 1666464484
transform 1 0 40544 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_354
timestamp 1666464484
transform 1 0 40992 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_49_357
timestamp 1666464484
transform 1 0 41328 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_389
timestamp 1666464484
transform 1 0 44912 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_405
timestamp 1666464484
transform 1 0 46704 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_413
timestamp 1666464484
transform 1 0 47600 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_417
timestamp 1666464484
transform 1 0 48048 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_419
timestamp 1666464484
transform 1 0 48272 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_2
timestamp 1666464484
transform 1 0 1568 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_34
timestamp 1666464484
transform 1 0 5152 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_37
timestamp 1666464484
transform 1 0 5488 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_101
timestamp 1666464484
transform 1 0 12656 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_105
timestamp 1666464484
transform 1 0 13104 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_108
timestamp 1666464484
transform 1 0 13440 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_172
timestamp 1666464484
transform 1 0 20608 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_176
timestamp 1666464484
transform 1 0 21056 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_179
timestamp 1666464484
transform 1 0 21392 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_243
timestamp 1666464484
transform 1 0 28560 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_247
timestamp 1666464484
transform 1 0 29008 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_250
timestamp 1666464484
transform 1 0 29344 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_314
timestamp 1666464484
transform 1 0 36512 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_318
timestamp 1666464484
transform 1 0 36960 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_321
timestamp 1666464484
transform 1 0 37296 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_385
timestamp 1666464484
transform 1 0 44464 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_389
timestamp 1666464484
transform 1 0 44912 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_392
timestamp 1666464484
transform 1 0 45248 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_400
timestamp 1666464484
transform 1 0 46144 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_403
timestamp 1666464484
transform 1 0 46480 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_419
timestamp 1666464484
transform 1 0 48272 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_2
timestamp 1666464484
transform 1 0 1568 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_66
timestamp 1666464484
transform 1 0 8736 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_70
timestamp 1666464484
transform 1 0 9184 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_73
timestamp 1666464484
transform 1 0 9520 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_137
timestamp 1666464484
transform 1 0 16688 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_141
timestamp 1666464484
transform 1 0 17136 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_144
timestamp 1666464484
transform 1 0 17472 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_208
timestamp 1666464484
transform 1 0 24640 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_212
timestamp 1666464484
transform 1 0 25088 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_215
timestamp 1666464484
transform 1 0 25424 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_279
timestamp 1666464484
transform 1 0 32592 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_283
timestamp 1666464484
transform 1 0 33040 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_286
timestamp 1666464484
transform 1 0 33376 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_350
timestamp 1666464484
transform 1 0 40544 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_354
timestamp 1666464484
transform 1 0 40992 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_51_357
timestamp 1666464484
transform 1 0 41328 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_389
timestamp 1666464484
transform 1 0 44912 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_405
timestamp 1666464484
transform 1 0 46704 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_413
timestamp 1666464484
transform 1 0 47600 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_417
timestamp 1666464484
transform 1 0 48048 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_419
timestamp 1666464484
transform 1 0 48272 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_52_2
timestamp 1666464484
transform 1 0 1568 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_34
timestamp 1666464484
transform 1 0 5152 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_37
timestamp 1666464484
transform 1 0 5488 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_101
timestamp 1666464484
transform 1 0 12656 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_105
timestamp 1666464484
transform 1 0 13104 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_108
timestamp 1666464484
transform 1 0 13440 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_172
timestamp 1666464484
transform 1 0 20608 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_176
timestamp 1666464484
transform 1 0 21056 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_179
timestamp 1666464484
transform 1 0 21392 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_243
timestamp 1666464484
transform 1 0 28560 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_247
timestamp 1666464484
transform 1 0 29008 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_250
timestamp 1666464484
transform 1 0 29344 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_314
timestamp 1666464484
transform 1 0 36512 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_318
timestamp 1666464484
transform 1 0 36960 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_321
timestamp 1666464484
transform 1 0 37296 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_385
timestamp 1666464484
transform 1 0 44464 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_389
timestamp 1666464484
transform 1 0 44912 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_392
timestamp 1666464484
transform 1 0 45248 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_400
timestamp 1666464484
transform 1 0 46144 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_403
timestamp 1666464484
transform 1 0 46480 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_419
timestamp 1666464484
transform 1 0 48272 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_2
timestamp 1666464484
transform 1 0 1568 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_66
timestamp 1666464484
transform 1 0 8736 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_70
timestamp 1666464484
transform 1 0 9184 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_73
timestamp 1666464484
transform 1 0 9520 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_137
timestamp 1666464484
transform 1 0 16688 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_141
timestamp 1666464484
transform 1 0 17136 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_144
timestamp 1666464484
transform 1 0 17472 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_208
timestamp 1666464484
transform 1 0 24640 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_212
timestamp 1666464484
transform 1 0 25088 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_215
timestamp 1666464484
transform 1 0 25424 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_279
timestamp 1666464484
transform 1 0 32592 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_283
timestamp 1666464484
transform 1 0 33040 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_286
timestamp 1666464484
transform 1 0 33376 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_350
timestamp 1666464484
transform 1 0 40544 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_354
timestamp 1666464484
transform 1 0 40992 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_53_357
timestamp 1666464484
transform 1 0 41328 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_389
timestamp 1666464484
transform 1 0 44912 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_399
timestamp 1666464484
transform 1 0 46032 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_403
timestamp 1666464484
transform 1 0 46480 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_419
timestamp 1666464484
transform 1 0 48272 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_2
timestamp 1666464484
transform 1 0 1568 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_7
timestamp 1666464484
transform 1 0 2128 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_23
timestamp 1666464484
transform 1 0 3920 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_31
timestamp 1666464484
transform 1 0 4816 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_37
timestamp 1666464484
transform 1 0 5488 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_69
timestamp 1666464484
transform 1 0 9072 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_72
timestamp 1666464484
transform 1 0 9408 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_104
timestamp 1666464484
transform 1 0 12992 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_107
timestamp 1666464484
transform 1 0 13328 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_139
timestamp 1666464484
transform 1 0 16912 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_142
timestamp 1666464484
transform 1 0 17248 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_174
timestamp 1666464484
transform 1 0 20832 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_177
timestamp 1666464484
transform 1 0 21168 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_209
timestamp 1666464484
transform 1 0 24752 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_212
timestamp 1666464484
transform 1 0 25088 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_244
timestamp 1666464484
transform 1 0 28672 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_247
timestamp 1666464484
transform 1 0 29008 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_279
timestamp 1666464484
transform 1 0 32592 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_282
timestamp 1666464484
transform 1 0 32928 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_314
timestamp 1666464484
transform 1 0 36512 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_317
timestamp 1666464484
transform 1 0 36848 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_349
timestamp 1666464484
transform 1 0 40432 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_352
timestamp 1666464484
transform 1 0 40768 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_368
timestamp 1666464484
transform 1 0 42560 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_376
timestamp 1666464484
transform 1 0 43456 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_380
timestamp 1666464484
transform 1 0 43904 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_384
timestamp 1666464484
transform 1 0 44352 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_387
timestamp 1666464484
transform 1 0 44688 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_403
timestamp 1666464484
transform 1 0 46480 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_419
timestamp 1666464484
transform 1 0 48272 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1666464484
transform -1 0 48608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1666464484
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1666464484
transform -1 0 48608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1666464484
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1666464484
transform -1 0 48608 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1666464484
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1666464484
transform -1 0 48608 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1666464484
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1666464484
transform -1 0 48608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1666464484
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1666464484
transform -1 0 48608 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1666464484
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1666464484
transform -1 0 48608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1666464484
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1666464484
transform -1 0 48608 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1666464484
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1666464484
transform -1 0 48608 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1666464484
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1666464484
transform -1 0 48608 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1666464484
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1666464484
transform -1 0 48608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1666464484
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1666464484
transform -1 0 48608 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1666464484
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1666464484
transform -1 0 48608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1666464484
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1666464484
transform -1 0 48608 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1666464484
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1666464484
transform -1 0 48608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1666464484
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1666464484
transform -1 0 48608 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1666464484
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1666464484
transform -1 0 48608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_34
timestamp 1666464484
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_35
timestamp 1666464484
transform -1 0 48608 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_36
timestamp 1666464484
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_37
timestamp 1666464484
transform -1 0 48608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_38
timestamp 1666464484
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_39
timestamp 1666464484
transform -1 0 48608 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_40
timestamp 1666464484
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_41
timestamp 1666464484
transform -1 0 48608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_42
timestamp 1666464484
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_43
timestamp 1666464484
transform -1 0 48608 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_44
timestamp 1666464484
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_45
timestamp 1666464484
transform -1 0 48608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_46
timestamp 1666464484
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_47
timestamp 1666464484
transform -1 0 48608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_48
timestamp 1666464484
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_49
timestamp 1666464484
transform -1 0 48608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_50
timestamp 1666464484
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_51
timestamp 1666464484
transform -1 0 48608 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_52
timestamp 1666464484
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_53
timestamp 1666464484
transform -1 0 48608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_54
timestamp 1666464484
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_55
timestamp 1666464484
transform -1 0 48608 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_56
timestamp 1666464484
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_57
timestamp 1666464484
transform -1 0 48608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_58
timestamp 1666464484
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_59
timestamp 1666464484
transform -1 0 48608 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_60
timestamp 1666464484
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_61
timestamp 1666464484
transform -1 0 48608 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_62
timestamp 1666464484
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_63
timestamp 1666464484
transform -1 0 48608 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_64
timestamp 1666464484
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_65
timestamp 1666464484
transform -1 0 48608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_66
timestamp 1666464484
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_67
timestamp 1666464484
transform -1 0 48608 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_68
timestamp 1666464484
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_69
timestamp 1666464484
transform -1 0 48608 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_70
timestamp 1666464484
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_71
timestamp 1666464484
transform -1 0 48608 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_72
timestamp 1666464484
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_73
timestamp 1666464484
transform -1 0 48608 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_74
timestamp 1666464484
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_75
timestamp 1666464484
transform -1 0 48608 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_76
timestamp 1666464484
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_77
timestamp 1666464484
transform -1 0 48608 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_78
timestamp 1666464484
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_79
timestamp 1666464484
transform -1 0 48608 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_80
timestamp 1666464484
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_81
timestamp 1666464484
transform -1 0 48608 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_82
timestamp 1666464484
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_83
timestamp 1666464484
transform -1 0 48608 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_84
timestamp 1666464484
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_85
timestamp 1666464484
transform -1 0 48608 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_86
timestamp 1666464484
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_87
timestamp 1666464484
transform -1 0 48608 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_88
timestamp 1666464484
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_89
timestamp 1666464484
transform -1 0 48608 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_90
timestamp 1666464484
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_91
timestamp 1666464484
transform -1 0 48608 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_92
timestamp 1666464484
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_93
timestamp 1666464484
transform -1 0 48608 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_94
timestamp 1666464484
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_95
timestamp 1666464484
transform -1 0 48608 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_96
timestamp 1666464484
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_97
timestamp 1666464484
transform -1 0 48608 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_98
timestamp 1666464484
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_99
timestamp 1666464484
transform -1 0 48608 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_100
timestamp 1666464484
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_101
timestamp 1666464484
transform -1 0 48608 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_102
timestamp 1666464484
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_103
timestamp 1666464484
transform -1 0 48608 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_104
timestamp 1666464484
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_105
timestamp 1666464484
transform -1 0 48608 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_106
timestamp 1666464484
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_107
timestamp 1666464484
transform -1 0 48608 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_108
timestamp 1666464484
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_109
timestamp 1666464484
transform -1 0 48608 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_110 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_111
timestamp 1666464484
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_112
timestamp 1666464484
transform 1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_113
timestamp 1666464484
transform 1 0 17024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_114
timestamp 1666464484
transform 1 0 20944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_115
timestamp 1666464484
transform 1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_116
timestamp 1666464484
transform 1 0 28784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_117
timestamp 1666464484
transform 1 0 32704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_118
timestamp 1666464484
transform 1 0 36624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_119
timestamp 1666464484
transform 1 0 40544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_120
timestamp 1666464484
transform 1 0 44464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_121
timestamp 1666464484
transform 1 0 9296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_122
timestamp 1666464484
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_123
timestamp 1666464484
transform 1 0 25200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_124
timestamp 1666464484
transform 1 0 33152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_125
timestamp 1666464484
transform 1 0 41104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_126
timestamp 1666464484
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_127
timestamp 1666464484
transform 1 0 13216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_128
timestamp 1666464484
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_129
timestamp 1666464484
transform 1 0 29120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_130
timestamp 1666464484
transform 1 0 37072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_131
timestamp 1666464484
transform 1 0 45024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_132
timestamp 1666464484
transform 1 0 9296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_133
timestamp 1666464484
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_134
timestamp 1666464484
transform 1 0 25200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_135
timestamp 1666464484
transform 1 0 33152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_136
timestamp 1666464484
transform 1 0 41104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_137
timestamp 1666464484
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_138
timestamp 1666464484
transform 1 0 13216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_139
timestamp 1666464484
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_140
timestamp 1666464484
transform 1 0 29120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_141
timestamp 1666464484
transform 1 0 37072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_142
timestamp 1666464484
transform 1 0 45024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_143
timestamp 1666464484
transform 1 0 9296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_144
timestamp 1666464484
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_145
timestamp 1666464484
transform 1 0 25200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_146
timestamp 1666464484
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_147
timestamp 1666464484
transform 1 0 41104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_148
timestamp 1666464484
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_149
timestamp 1666464484
transform 1 0 13216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_150
timestamp 1666464484
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_151
timestamp 1666464484
transform 1 0 29120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_152
timestamp 1666464484
transform 1 0 37072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_153
timestamp 1666464484
transform 1 0 45024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_154
timestamp 1666464484
transform 1 0 9296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_155
timestamp 1666464484
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_156
timestamp 1666464484
transform 1 0 25200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_157
timestamp 1666464484
transform 1 0 33152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_158
timestamp 1666464484
transform 1 0 41104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_159
timestamp 1666464484
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_160
timestamp 1666464484
transform 1 0 13216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_161
timestamp 1666464484
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_162
timestamp 1666464484
transform 1 0 29120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_163
timestamp 1666464484
transform 1 0 37072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_164
timestamp 1666464484
transform 1 0 45024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_165
timestamp 1666464484
transform 1 0 9296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_166
timestamp 1666464484
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_167
timestamp 1666464484
transform 1 0 25200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_168
timestamp 1666464484
transform 1 0 33152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_169
timestamp 1666464484
transform 1 0 41104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_170
timestamp 1666464484
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_171
timestamp 1666464484
transform 1 0 13216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_172
timestamp 1666464484
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_173
timestamp 1666464484
transform 1 0 29120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_174
timestamp 1666464484
transform 1 0 37072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_175
timestamp 1666464484
transform 1 0 45024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_176
timestamp 1666464484
transform 1 0 9296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_177
timestamp 1666464484
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_178
timestamp 1666464484
transform 1 0 25200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_179
timestamp 1666464484
transform 1 0 33152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_180
timestamp 1666464484
transform 1 0 41104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_181
timestamp 1666464484
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_182
timestamp 1666464484
transform 1 0 13216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_183
timestamp 1666464484
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_184
timestamp 1666464484
transform 1 0 29120 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_185
timestamp 1666464484
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_186
timestamp 1666464484
transform 1 0 45024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_187
timestamp 1666464484
transform 1 0 9296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_188
timestamp 1666464484
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_189
timestamp 1666464484
transform 1 0 25200 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_190
timestamp 1666464484
transform 1 0 33152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_191
timestamp 1666464484
transform 1 0 41104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_192
timestamp 1666464484
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_193
timestamp 1666464484
transform 1 0 13216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_194
timestamp 1666464484
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_195
timestamp 1666464484
transform 1 0 29120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_196
timestamp 1666464484
transform 1 0 37072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_197
timestamp 1666464484
transform 1 0 45024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_198
timestamp 1666464484
transform 1 0 9296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_199
timestamp 1666464484
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_200
timestamp 1666464484
transform 1 0 25200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_201
timestamp 1666464484
transform 1 0 33152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_202
timestamp 1666464484
transform 1 0 41104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_203
timestamp 1666464484
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_204
timestamp 1666464484
transform 1 0 13216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_205
timestamp 1666464484
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_206
timestamp 1666464484
transform 1 0 29120 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_207
timestamp 1666464484
transform 1 0 37072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_208
timestamp 1666464484
transform 1 0 45024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_209
timestamp 1666464484
transform 1 0 9296 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_210
timestamp 1666464484
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_211
timestamp 1666464484
transform 1 0 25200 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_212
timestamp 1666464484
transform 1 0 33152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_213
timestamp 1666464484
transform 1 0 41104 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_214
timestamp 1666464484
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_215
timestamp 1666464484
transform 1 0 13216 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_216
timestamp 1666464484
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_217
timestamp 1666464484
transform 1 0 29120 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_218
timestamp 1666464484
transform 1 0 37072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_219
timestamp 1666464484
transform 1 0 45024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_220
timestamp 1666464484
transform 1 0 9296 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_221
timestamp 1666464484
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_222
timestamp 1666464484
transform 1 0 25200 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_223
timestamp 1666464484
transform 1 0 33152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_224
timestamp 1666464484
transform 1 0 41104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_225
timestamp 1666464484
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_226
timestamp 1666464484
transform 1 0 13216 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_227
timestamp 1666464484
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_228
timestamp 1666464484
transform 1 0 29120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_229
timestamp 1666464484
transform 1 0 37072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_230
timestamp 1666464484
transform 1 0 45024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_231
timestamp 1666464484
transform 1 0 9296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_232
timestamp 1666464484
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_233
timestamp 1666464484
transform 1 0 25200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_234
timestamp 1666464484
transform 1 0 33152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_235
timestamp 1666464484
transform 1 0 41104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_236
timestamp 1666464484
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_237
timestamp 1666464484
transform 1 0 13216 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_238
timestamp 1666464484
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_239
timestamp 1666464484
transform 1 0 29120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_240
timestamp 1666464484
transform 1 0 37072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_241
timestamp 1666464484
transform 1 0 45024 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_242
timestamp 1666464484
transform 1 0 9296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_243
timestamp 1666464484
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_244
timestamp 1666464484
transform 1 0 25200 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_245
timestamp 1666464484
transform 1 0 33152 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_246
timestamp 1666464484
transform 1 0 41104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_247
timestamp 1666464484
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_248
timestamp 1666464484
transform 1 0 13216 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_249
timestamp 1666464484
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_250
timestamp 1666464484
transform 1 0 29120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_251
timestamp 1666464484
transform 1 0 37072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_252
timestamp 1666464484
transform 1 0 45024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_253
timestamp 1666464484
transform 1 0 9296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_254
timestamp 1666464484
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_255
timestamp 1666464484
transform 1 0 25200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_256
timestamp 1666464484
transform 1 0 33152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_257
timestamp 1666464484
transform 1 0 41104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_258
timestamp 1666464484
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_259
timestamp 1666464484
transform 1 0 13216 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_260
timestamp 1666464484
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_261
timestamp 1666464484
transform 1 0 29120 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_262
timestamp 1666464484
transform 1 0 37072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_263
timestamp 1666464484
transform 1 0 45024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_264
timestamp 1666464484
transform 1 0 9296 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_265
timestamp 1666464484
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_266
timestamp 1666464484
transform 1 0 25200 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_267
timestamp 1666464484
transform 1 0 33152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_268
timestamp 1666464484
transform 1 0 41104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_269
timestamp 1666464484
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_270
timestamp 1666464484
transform 1 0 13216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_271
timestamp 1666464484
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_272
timestamp 1666464484
transform 1 0 29120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_273
timestamp 1666464484
transform 1 0 37072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_274
timestamp 1666464484
transform 1 0 45024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_275
timestamp 1666464484
transform 1 0 9296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_276
timestamp 1666464484
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_277
timestamp 1666464484
transform 1 0 25200 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_278
timestamp 1666464484
transform 1 0 33152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_279
timestamp 1666464484
transform 1 0 41104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_280
timestamp 1666464484
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_281
timestamp 1666464484
transform 1 0 13216 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_282
timestamp 1666464484
transform 1 0 21168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_283
timestamp 1666464484
transform 1 0 29120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_284
timestamp 1666464484
transform 1 0 37072 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_285
timestamp 1666464484
transform 1 0 45024 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_286
timestamp 1666464484
transform 1 0 9296 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_287
timestamp 1666464484
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_288
timestamp 1666464484
transform 1 0 25200 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_289
timestamp 1666464484
transform 1 0 33152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_290
timestamp 1666464484
transform 1 0 41104 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_291
timestamp 1666464484
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_292
timestamp 1666464484
transform 1 0 13216 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_293
timestamp 1666464484
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_294
timestamp 1666464484
transform 1 0 29120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_295
timestamp 1666464484
transform 1 0 37072 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_296
timestamp 1666464484
transform 1 0 45024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_297
timestamp 1666464484
transform 1 0 9296 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_298
timestamp 1666464484
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_299
timestamp 1666464484
transform 1 0 25200 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_300
timestamp 1666464484
transform 1 0 33152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_301
timestamp 1666464484
transform 1 0 41104 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_302
timestamp 1666464484
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_303
timestamp 1666464484
transform 1 0 13216 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_304
timestamp 1666464484
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_305
timestamp 1666464484
transform 1 0 29120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_306
timestamp 1666464484
transform 1 0 37072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_307
timestamp 1666464484
transform 1 0 45024 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_308
timestamp 1666464484
transform 1 0 9296 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_309
timestamp 1666464484
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_310
timestamp 1666464484
transform 1 0 25200 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_311
timestamp 1666464484
transform 1 0 33152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_312
timestamp 1666464484
transform 1 0 41104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_313
timestamp 1666464484
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_314
timestamp 1666464484
transform 1 0 13216 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_315
timestamp 1666464484
transform 1 0 21168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_316
timestamp 1666464484
transform 1 0 29120 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_317
timestamp 1666464484
transform 1 0 37072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_318
timestamp 1666464484
transform 1 0 45024 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_319
timestamp 1666464484
transform 1 0 9296 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_320
timestamp 1666464484
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_321
timestamp 1666464484
transform 1 0 25200 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_322
timestamp 1666464484
transform 1 0 33152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_323
timestamp 1666464484
transform 1 0 41104 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_324
timestamp 1666464484
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_325
timestamp 1666464484
transform 1 0 13216 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_326
timestamp 1666464484
transform 1 0 21168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_327
timestamp 1666464484
transform 1 0 29120 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_328
timestamp 1666464484
transform 1 0 37072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_329
timestamp 1666464484
transform 1 0 45024 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_330
timestamp 1666464484
transform 1 0 9296 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_331
timestamp 1666464484
transform 1 0 17248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_332
timestamp 1666464484
transform 1 0 25200 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_333
timestamp 1666464484
transform 1 0 33152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_334
timestamp 1666464484
transform 1 0 41104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_335
timestamp 1666464484
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_336
timestamp 1666464484
transform 1 0 13216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_337
timestamp 1666464484
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_338
timestamp 1666464484
transform 1 0 29120 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_339
timestamp 1666464484
transform 1 0 37072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_340
timestamp 1666464484
transform 1 0 45024 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_341
timestamp 1666464484
transform 1 0 9296 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_342
timestamp 1666464484
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_343
timestamp 1666464484
transform 1 0 25200 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_344
timestamp 1666464484
transform 1 0 33152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_345
timestamp 1666464484
transform 1 0 41104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_346
timestamp 1666464484
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_347
timestamp 1666464484
transform 1 0 13216 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_348
timestamp 1666464484
transform 1 0 21168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_349
timestamp 1666464484
transform 1 0 29120 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_350
timestamp 1666464484
transform 1 0 37072 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_351
timestamp 1666464484
transform 1 0 45024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_352
timestamp 1666464484
transform 1 0 9296 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_353
timestamp 1666464484
transform 1 0 17248 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_354
timestamp 1666464484
transform 1 0 25200 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_355
timestamp 1666464484
transform 1 0 33152 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_356
timestamp 1666464484
transform 1 0 41104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_357
timestamp 1666464484
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_358
timestamp 1666464484
transform 1 0 13216 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_359
timestamp 1666464484
transform 1 0 21168 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_360
timestamp 1666464484
transform 1 0 29120 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_361
timestamp 1666464484
transform 1 0 37072 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_362
timestamp 1666464484
transform 1 0 45024 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_363
timestamp 1666464484
transform 1 0 9296 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_364
timestamp 1666464484
transform 1 0 17248 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_365
timestamp 1666464484
transform 1 0 25200 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_366
timestamp 1666464484
transform 1 0 33152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_367
timestamp 1666464484
transform 1 0 41104 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_368
timestamp 1666464484
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_369
timestamp 1666464484
transform 1 0 13216 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_370
timestamp 1666464484
transform 1 0 21168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_371
timestamp 1666464484
transform 1 0 29120 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_372
timestamp 1666464484
transform 1 0 37072 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_373
timestamp 1666464484
transform 1 0 45024 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_374
timestamp 1666464484
transform 1 0 9296 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_375
timestamp 1666464484
transform 1 0 17248 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_376
timestamp 1666464484
transform 1 0 25200 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_377
timestamp 1666464484
transform 1 0 33152 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_378
timestamp 1666464484
transform 1 0 41104 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_379
timestamp 1666464484
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_380
timestamp 1666464484
transform 1 0 13216 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_381
timestamp 1666464484
transform 1 0 21168 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_382
timestamp 1666464484
transform 1 0 29120 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_383
timestamp 1666464484
transform 1 0 37072 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_384
timestamp 1666464484
transform 1 0 45024 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_385
timestamp 1666464484
transform 1 0 9296 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_386
timestamp 1666464484
transform 1 0 17248 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_387
timestamp 1666464484
transform 1 0 25200 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_388
timestamp 1666464484
transform 1 0 33152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_389
timestamp 1666464484
transform 1 0 41104 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_390
timestamp 1666464484
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_391
timestamp 1666464484
transform 1 0 13216 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_392
timestamp 1666464484
transform 1 0 21168 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_393
timestamp 1666464484
transform 1 0 29120 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_394
timestamp 1666464484
transform 1 0 37072 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_395
timestamp 1666464484
transform 1 0 45024 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_396
timestamp 1666464484
transform 1 0 9296 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_397
timestamp 1666464484
transform 1 0 17248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_398
timestamp 1666464484
transform 1 0 25200 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_399
timestamp 1666464484
transform 1 0 33152 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_400
timestamp 1666464484
transform 1 0 41104 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_401
timestamp 1666464484
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_402
timestamp 1666464484
transform 1 0 13216 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_403
timestamp 1666464484
transform 1 0 21168 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_404
timestamp 1666464484
transform 1 0 29120 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_405
timestamp 1666464484
transform 1 0 37072 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_406
timestamp 1666464484
transform 1 0 45024 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_407
timestamp 1666464484
transform 1 0 9296 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_408
timestamp 1666464484
transform 1 0 17248 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_409
timestamp 1666464484
transform 1 0 25200 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_410
timestamp 1666464484
transform 1 0 33152 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_411
timestamp 1666464484
transform 1 0 41104 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_412
timestamp 1666464484
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_413
timestamp 1666464484
transform 1 0 9184 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_414
timestamp 1666464484
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_415
timestamp 1666464484
transform 1 0 17024 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_416
timestamp 1666464484
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_417
timestamp 1666464484
transform 1 0 24864 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_418
timestamp 1666464484
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_419
timestamp 1666464484
transform 1 0 32704 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_420
timestamp 1666464484
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_421
timestamp 1666464484
transform 1 0 40544 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_422
timestamp 1666464484
transform 1 0 44464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _078_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 43568 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _079_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 37968 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _080_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 34048 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _081_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 39312 0 1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _082_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 41440 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _083_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 41664 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _084_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 42560 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _085_
timestamp 1666464484
transform -1 0 44016 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _086_
timestamp 1666464484
transform -1 0 40544 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _087_
timestamp 1666464484
transform -1 0 43456 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _088_
timestamp 1666464484
transform -1 0 40992 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _089_
timestamp 1666464484
transform -1 0 43792 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _090_
timestamp 1666464484
transform -1 0 43120 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _091_
timestamp 1666464484
transform -1 0 44912 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _092_
timestamp 1666464484
transform 1 0 41216 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _093_
timestamp 1666464484
transform -1 0 42896 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _094_
timestamp 1666464484
transform -1 0 42672 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _095_
timestamp 1666464484
transform -1 0 43232 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _096_
timestamp 1666464484
transform -1 0 43456 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _097_
timestamp 1666464484
transform 1 0 41440 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _098_
timestamp 1666464484
transform -1 0 40992 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _099_
timestamp 1666464484
transform 1 0 41440 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _100_
timestamp 1666464484
transform -1 0 40992 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _101_
timestamp 1666464484
transform -1 0 41328 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _102_
timestamp 1666464484
transform 1 0 38752 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _103_
timestamp 1666464484
transform -1 0 40208 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _104_
timestamp 1666464484
transform -1 0 39424 0 -1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _105_
timestamp 1666464484
transform -1 0 41104 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _106_
timestamp 1666464484
transform -1 0 38528 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _107_
timestamp 1666464484
transform -1 0 40208 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _108_
timestamp 1666464484
transform -1 0 39088 0 1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _109_
timestamp 1666464484
transform -1 0 39648 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _110_
timestamp 1666464484
transform -1 0 40768 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _111_
timestamp 1666464484
transform 1 0 35840 0 -1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _112_
timestamp 1666464484
transform -1 0 36736 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _113_
timestamp 1666464484
transform 1 0 34272 0 1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _114_
timestamp 1666464484
transform -1 0 35056 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _115_
timestamp 1666464484
transform -1 0 35616 0 -1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _116_
timestamp 1666464484
transform -1 0 38080 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _117_
timestamp 1666464484
transform -1 0 35392 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _118_
timestamp 1666464484
transform -1 0 35952 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _119_
timestamp 1666464484
transform -1 0 40992 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _120_
timestamp 1666464484
transform -1 0 41104 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _121_
timestamp 1666464484
transform 1 0 35168 0 -1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _122_
timestamp 1666464484
transform -1 0 35056 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _123_
timestamp 1666464484
transform 1 0 35280 0 1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _124_
timestamp 1666464484
transform -1 0 34160 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _125_
timestamp 1666464484
transform 1 0 37072 0 -1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _126_
timestamp 1666464484
transform -1 0 33712 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _127_
timestamp 1666464484
transform 1 0 36176 0 -1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _128_
timestamp 1666464484
transform -1 0 32816 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _129_
timestamp 1666464484
transform -1 0 40992 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _130_
timestamp 1666464484
transform 1 0 37408 0 1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _131_
timestamp 1666464484
transform -1 0 31472 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _132_
timestamp 1666464484
transform 1 0 36848 0 -1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _133_
timestamp 1666464484
transform -1 0 31472 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _134_
timestamp 1666464484
transform 1 0 37408 0 1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _135_
timestamp 1666464484
transform -1 0 32368 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _136_
timestamp 1666464484
transform 1 0 37296 0 -1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _137_
timestamp 1666464484
transform -1 0 31808 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _138_
timestamp 1666464484
transform -1 0 40432 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _139_
timestamp 1666464484
transform 1 0 37744 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _140_
timestamp 1666464484
transform -1 0 31696 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _141_
timestamp 1666464484
transform 1 0 37744 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _142_
timestamp 1666464484
transform -1 0 31584 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _143_
timestamp 1666464484
transform 1 0 37856 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _144_
timestamp 1666464484
transform -1 0 30688 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _145_
timestamp 1666464484
transform 1 0 37968 0 -1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _146_
timestamp 1666464484
transform 1 0 29008 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _147_
timestamp 1666464484
transform -1 0 39872 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _148_
timestamp 1666464484
transform 1 0 37744 0 1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _149_
timestamp 1666464484
transform 1 0 29456 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _150_
timestamp 1666464484
transform 1 0 37744 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _151_
timestamp 1666464484
transform -1 0 29680 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _152_
timestamp 1666464484
transform 1 0 37072 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _153_
timestamp 1666464484
transform -1 0 27664 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _154_
timestamp 1666464484
transform 1 0 29568 0 1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _155_
timestamp 1666464484
transform -1 0 28560 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _156_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 3360 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _157_
timestamp 1666464484
transform 1 0 5936 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _158_
timestamp 1666464484
transform 1 0 17248 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _159_
timestamp 1666464484
transform 1 0 3248 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _160_
timestamp 1666464484
transform 1 0 5600 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _161_
timestamp 1666464484
transform 1 0 13552 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _162_
timestamp 1666464484
transform 1 0 1904 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _163_
timestamp 1666464484
transform -1 0 5152 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _164_
timestamp 1666464484
transform 1 0 9856 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _165_
timestamp 1666464484
transform 1 0 29456 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _166_
timestamp 1666464484
transform 1 0 33712 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _167_
timestamp 1666464484
transform 1 0 34496 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _168_
timestamp 1666464484
transform 1 0 37408 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _169_
timestamp 1666464484
transform 1 0 35280 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _170_
timestamp 1666464484
transform 1 0 35504 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _171_
timestamp 1666464484
transform 1 0 35616 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _172_
timestamp 1666464484
transform 1 0 37408 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _173_
timestamp 1666464484
transform 1 0 35056 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _174_
timestamp 1666464484
transform 1 0 33712 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _175_
timestamp 1666464484
transform 1 0 32928 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _176_
timestamp 1666464484
transform 1 0 29792 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _177_
timestamp 1666464484
transform 1 0 25760 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _178_
timestamp 1666464484
transform 1 0 25536 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _179_
timestamp 1666464484
transform 1 0 25424 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _180_
timestamp 1666464484
transform 1 0 25536 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _181_
timestamp 1666464484
transform -1 0 23520 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _182_
timestamp 1666464484
transform 1 0 17808 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _183_
timestamp 1666464484
transform 1 0 16912 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _184_
timestamp 1666464484
transform 1 0 13888 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _185_
timestamp 1666464484
transform 1 0 16016 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _186_
timestamp 1666464484
transform 1 0 16464 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _187_
timestamp 1666464484
transform 1 0 17472 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _188_
timestamp 1666464484
transform 1 0 19376 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _189_
timestamp 1666464484
transform 1 0 24976 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _190_
timestamp 1666464484
transform 1 0 27328 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _191_
timestamp 1666464484
transform 1 0 29456 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _192_
timestamp 1666464484
transform 1 0 29456 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _193_
timestamp 1666464484
transform 1 0 29456 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _194_
timestamp 1666464484
transform 1 0 28336 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _195_
timestamp 1666464484
transform -1 0 24752 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _196_
timestamp 1666464484
transform 1 0 12432 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _205_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 37968 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _206_
timestamp 1666464484
transform -1 0 18480 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clock dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 19488 0 -1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_0__f_clock
timestamp 1666464484
transform -1 0 17024 0 -1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_1__f_clock
timestamp 1666464484
transform -1 0 17024 0 -1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_2__f_clock
timestamp 1666464484
transform 1 0 22848 0 1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_3__f_clock
timestamp 1666464484
transform 1 0 26656 0 -1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1666464484
transform 1 0 1680 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1666464484
transform 1 0 1680 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1666464484
transform 1 0 1680 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output4
timestamp 1666464484
transform 1 0 47600 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output5 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 46704 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output6
timestamp 1666464484
transform 1 0 46704 0 -1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output7
timestamp 1666464484
transform 1 0 46704 0 1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output8
timestamp 1666464484
transform 1 0 46704 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output9
timestamp 1666464484
transform 1 0 46704 0 1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output10
timestamp 1666464484
transform 1 0 46704 0 1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output11
timestamp 1666464484
transform 1 0 46704 0 1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output12
timestamp 1666464484
transform 1 0 46704 0 1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output13
timestamp 1666464484
transform 1 0 46704 0 1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output14
timestamp 1666464484
transform 1 0 46704 0 -1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output15
timestamp 1666464484
transform 1 0 46704 0 -1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output16
timestamp 1666464484
transform 1 0 46704 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output17
timestamp 1666464484
transform 1 0 46704 0 -1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output18
timestamp 1666464484
transform 1 0 46704 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output19
timestamp 1666464484
transform 1 0 46704 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output20
timestamp 1666464484
transform 1 0 46704 0 -1 37632
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output21
timestamp 1666464484
transform 1 0 46704 0 -1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output22
timestamp 1666464484
transform 1 0 46704 0 1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output23
timestamp 1666464484
transform 1 0 46704 0 1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output24
timestamp 1666464484
transform 1 0 46704 0 1 42336
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output25
timestamp 1666464484
transform 1 0 46704 0 1 43904
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output26
timestamp 1666464484
transform 1 0 46704 0 1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output27
timestamp 1666464484
transform 1 0 46704 0 1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output28
timestamp 1666464484
transform 1 0 46704 0 -1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output29
timestamp 1666464484
transform 1 0 44912 0 1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output30
timestamp 1666464484
transform 1 0 46704 0 1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output31
timestamp 1666464484
transform 1 0 46704 0 -1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output32
timestamp 1666464484
transform 1 0 46704 0 -1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output33
timestamp 1666464484
transform 1 0 46704 0 -1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output34
timestamp 1666464484
transform 1 0 46704 0 -1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output35
timestamp 1666464484
transform 1 0 46704 0 -1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output36
timestamp 1666464484
transform 1 0 46704 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output37
timestamp 1666464484
transform -1 0 3248 0 1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spi_core_38 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 8960 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spi_core_39
timestamp 1666464484
transform -1 0 14448 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spi_core_40
timestamp 1666464484
transform -1 0 19936 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spi_core_41
timestamp 1666464484
transform 1 0 24304 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spi_core_42
timestamp 1666464484
transform -1 0 2128 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spi_core_43
timestamp 1666464484
transform -1 0 2128 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spi_core_44
timestamp 1666464484
transform -1 0 2128 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  spi_core_45 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 2128 0 1 45472
box -86 -86 534 870
<< labels >>
flabel metal2 s 2856 -960 3080 480 0 FreeSans 896 90 0 0 clock
port 0 nsew signal input
flabel metal3 s 49520 1512 50960 1736 0 FreeSans 896 0 0 0 clock_out
port 1 nsew signal tristate
flabel metal3 s 49520 2968 50960 3192 0 FreeSans 896 0 0 0 data_out[0]
port 2 nsew signal tristate
flabel metal3 s 49520 17528 50960 17752 0 FreeSans 896 0 0 0 data_out[10]
port 3 nsew signal tristate
flabel metal3 s 49520 18984 50960 19208 0 FreeSans 896 0 0 0 data_out[11]
port 4 nsew signal tristate
flabel metal3 s 49520 20440 50960 20664 0 FreeSans 896 0 0 0 data_out[12]
port 5 nsew signal tristate
flabel metal3 s 49520 21896 50960 22120 0 FreeSans 896 0 0 0 data_out[13]
port 6 nsew signal tristate
flabel metal3 s 49520 23352 50960 23576 0 FreeSans 896 0 0 0 data_out[14]
port 7 nsew signal tristate
flabel metal3 s 49520 24808 50960 25032 0 FreeSans 896 0 0 0 data_out[15]
port 8 nsew signal tristate
flabel metal3 s 49520 26264 50960 26488 0 FreeSans 896 0 0 0 data_out[16]
port 9 nsew signal tristate
flabel metal3 s 49520 27720 50960 27944 0 FreeSans 896 0 0 0 data_out[17]
port 10 nsew signal tristate
flabel metal3 s 49520 29176 50960 29400 0 FreeSans 896 0 0 0 data_out[18]
port 11 nsew signal tristate
flabel metal3 s 49520 30632 50960 30856 0 FreeSans 896 0 0 0 data_out[19]
port 12 nsew signal tristate
flabel metal3 s 49520 4424 50960 4648 0 FreeSans 896 0 0 0 data_out[1]
port 13 nsew signal tristate
flabel metal3 s 49520 32088 50960 32312 0 FreeSans 896 0 0 0 data_out[20]
port 14 nsew signal tristate
flabel metal3 s 49520 33544 50960 33768 0 FreeSans 896 0 0 0 data_out[21]
port 15 nsew signal tristate
flabel metal3 s 49520 35000 50960 35224 0 FreeSans 896 0 0 0 data_out[22]
port 16 nsew signal tristate
flabel metal3 s 49520 36456 50960 36680 0 FreeSans 896 0 0 0 data_out[23]
port 17 nsew signal tristate
flabel metal3 s 49520 37912 50960 38136 0 FreeSans 896 0 0 0 data_out[24]
port 18 nsew signal tristate
flabel metal3 s 49520 39368 50960 39592 0 FreeSans 896 0 0 0 data_out[25]
port 19 nsew signal tristate
flabel metal3 s 49520 40824 50960 41048 0 FreeSans 896 0 0 0 data_out[26]
port 20 nsew signal tristate
flabel metal3 s 49520 42280 50960 42504 0 FreeSans 896 0 0 0 data_out[27]
port 21 nsew signal tristate
flabel metal3 s 49520 43736 50960 43960 0 FreeSans 896 0 0 0 data_out[28]
port 22 nsew signal tristate
flabel metal3 s 49520 45192 50960 45416 0 FreeSans 896 0 0 0 data_out[29]
port 23 nsew signal tristate
flabel metal3 s 49520 5880 50960 6104 0 FreeSans 896 0 0 0 data_out[2]
port 24 nsew signal tristate
flabel metal3 s 49520 46648 50960 46872 0 FreeSans 896 0 0 0 data_out[30]
port 25 nsew signal tristate
flabel metal3 s 49520 48104 50960 48328 0 FreeSans 896 0 0 0 data_out[31]
port 26 nsew signal tristate
flabel metal3 s 49520 7336 50960 7560 0 FreeSans 896 0 0 0 data_out[3]
port 27 nsew signal tristate
flabel metal3 s 49520 8792 50960 9016 0 FreeSans 896 0 0 0 data_out[4]
port 28 nsew signal tristate
flabel metal3 s 49520 10248 50960 10472 0 FreeSans 896 0 0 0 data_out[5]
port 29 nsew signal tristate
flabel metal3 s 49520 11704 50960 11928 0 FreeSans 896 0 0 0 data_out[6]
port 30 nsew signal tristate
flabel metal3 s 49520 13160 50960 13384 0 FreeSans 896 0 0 0 data_out[7]
port 31 nsew signal tristate
flabel metal3 s 49520 14616 50960 14840 0 FreeSans 896 0 0 0 data_out[8]
port 32 nsew signal tristate
flabel metal3 s 49520 16072 50960 16296 0 FreeSans 896 0 0 0 data_out[9]
port 33 nsew signal tristate
flabel metal2 s 30296 -960 30520 480 0 FreeSans 896 90 0 0 la_data_in[0]
port 34 nsew signal input
flabel metal2 s 35784 -960 36008 480 0 FreeSans 896 90 0 0 la_data_in[1]
port 35 nsew signal input
flabel metal2 s 41272 -960 41496 480 0 FreeSans 896 90 0 0 la_data_in[2]
port 36 nsew signal input
flabel metal2 s 46760 -960 46984 480 0 FreeSans 896 90 0 0 la_data_in[3]
port 37 nsew signal input
flabel metal2 s 8344 -960 8568 480 0 FreeSans 896 90 0 0 la_oenb[0]
port 38 nsew signal tristate
flabel metal2 s 13832 -960 14056 480 0 FreeSans 896 90 0 0 la_oenb[1]
port 39 nsew signal tristate
flabel metal2 s 19320 -960 19544 480 0 FreeSans 896 90 0 0 la_oenb[2]
port 40 nsew signal tristate
flabel metal2 s 24808 -960 25032 480 0 FreeSans 896 90 0 0 la_oenb[3]
port 41 nsew signal tristate
flabel metal3 s -960 40264 480 40488 0 FreeSans 896 0 0 0 miso
port 42 nsew signal tristate
flabel metal3 s -960 46424 480 46648 0 FreeSans 896 0 0 0 miso_oeb
port 43 nsew signal tristate
flabel metal3 s -960 15624 480 15848 0 FreeSans 896 0 0 0 mosi
port 44 nsew signal input
flabel metal3 s -960 21784 480 22008 0 FreeSans 896 0 0 0 mosi_oeb
port 45 nsew signal tristate
flabel metal3 s -960 3304 480 3528 0 FreeSans 896 0 0 0 sclk
port 46 nsew signal input
flabel metal3 s -960 9464 480 9688 0 FreeSans 896 0 0 0 sclk_oeb
port 47 nsew signal tristate
flabel metal3 s -960 27944 480 28168 0 FreeSans 896 0 0 0 ss_n
port 48 nsew signal input
flabel metal3 s -960 34104 480 34328 0 FreeSans 896 0 0 0 ss_n_oeb
port 49 nsew signal tristate
flabel metal4 s 2034 3076 2654 46316 0 FreeSans 2560 90 0 0 vccd1
port 50 nsew power bidirectional
flabel metal4 s 38034 3076 38654 46316 0 FreeSans 2560 90 0 0 vccd1
port 50 nsew power bidirectional
flabel metal4 s 5754 3076 6374 46316 0 FreeSans 2560 90 0 0 vssd1
port 51 nsew ground bidirectional
flabel metal4 s 41754 3076 42374 46316 0 FreeSans 2560 90 0 0 vssd1
port 51 nsew ground bidirectional
rlabel metal1 24976 46256 24976 46256 0 vccd1
rlabel metal1 24976 45472 24976 45472 0 vssd1
rlabel metal2 33096 5600 33096 5600 0 _000_
rlabel metal2 34664 4928 34664 4928 0 _001_
rlabel metal2 35448 3920 35448 3920 0 _002_
rlabel metal2 44408 5600 44408 5600 0 _003_
rlabel metal2 37576 8176 37576 8176 0 _004_
rlabel metal2 36456 7616 36456 7616 0 _005_
rlabel metal2 36568 10192 36568 10192 0 _006_
rlabel metal2 38360 11536 38360 11536 0 _007_
rlabel metal2 36008 13272 36008 13272 0 _008_
rlabel metal2 37688 11088 37688 11088 0 _009_
rlabel metal3 35224 11480 35224 11480 0 _010_
rlabel metal2 33544 9296 33544 9296 0 _011_
rlabel metal3 28168 6552 28168 6552 0 _012_
rlabel metal2 26488 4480 26488 4480 0 _013_
rlabel metal3 28056 3416 28056 3416 0 _014_
rlabel metal3 27776 5880 27776 5880 0 _015_
rlabel metal2 24248 4592 24248 4592 0 _016_
rlabel metal3 22176 10024 22176 10024 0 _017_
rlabel metal2 17864 8064 17864 8064 0 _018_
rlabel metal3 16240 10696 16240 10696 0 _019_
rlabel metal3 25564 12712 25564 12712 0 _020_
rlabel metal3 18760 9688 18760 9688 0 _021_
rlabel metal3 26320 12376 26320 12376 0 _022_
rlabel metal3 27104 10808 27104 10808 0 _023_
rlabel metal3 29904 11480 29904 11480 0 _024_
rlabel metal3 29680 15848 29680 15848 0 _025_
rlabel metal2 30352 11480 30352 11480 0 _026_
rlabel metal2 30464 9912 30464 9912 0 _027_
rlabel metal3 30184 16296 30184 16296 0 _028_
rlabel metal2 29232 18536 29232 18536 0 _029_
rlabel metal2 23800 13664 23800 13664 0 _030_
rlabel metal3 14896 5992 14896 5992 0 _031_
rlabel metal2 38864 14728 38864 14728 0 _032_
rlabel metal3 36288 15288 36288 15288 0 _033_
rlabel metal2 36120 15792 36120 15792 0 _034_
rlabel metal2 34608 14728 34608 14728 0 _035_
rlabel metal2 35336 16520 35336 16520 0 _036_
rlabel metal2 35112 17360 35112 17360 0 _037_
rlabel metal2 39760 27832 39760 27832 0 _038_
rlabel metal2 40376 19656 40376 19656 0 _039_
rlabel metal2 35448 17472 35448 17472 0 _040_
rlabel metal2 35560 17920 35560 17920 0 _041_
rlabel metal2 37296 17080 37296 17080 0 _042_
rlabel metal3 34552 18312 34552 18312 0 _043_
rlabel metal2 40320 23576 40320 23576 0 _044_
rlabel metal3 34496 19096 34496 19096 0 _045_
rlabel metal3 34216 18536 34216 18536 0 _046_
rlabel metal2 32200 19544 32200 19544 0 _047_
rlabel metal3 34776 17752 34776 17752 0 _048_
rlabel metal2 39536 26936 39536 26936 0 _049_
rlabel metal3 34944 17080 34944 17080 0 _050_
rlabel metal2 31864 17248 31864 17248 0 _051_
rlabel metal2 30520 19712 30520 19712 0 _052_
rlabel metal2 30072 16520 30072 16520 0 _053_
rlabel metal2 38808 27496 38808 27496 0 _054_
rlabel metal3 30072 17640 30072 17640 0 _055_
rlabel metal2 29792 18648 29792 18648 0 _056_
rlabel metal2 27944 20776 27944 20776 0 _057_
rlabel metal3 29120 21000 29120 21000 0 _058_
rlabel metal2 41384 5040 41384 5040 0 _059_
rlabel metal2 39928 21000 39928 21000 0 _060_
rlabel metal2 34328 20048 34328 20048 0 _061_
rlabel metal3 41216 20664 41216 20664 0 _062_
rlabel metal2 41664 15848 41664 15848 0 _063_
rlabel metal2 41496 9464 41496 9464 0 _064_
rlabel metal3 43008 5320 43008 5320 0 _065_
rlabel metal3 41776 4984 41776 4984 0 _066_
rlabel metal3 42112 6664 42112 6664 0 _067_
rlabel metal3 43736 5880 43736 5880 0 _068_
rlabel metal3 41832 8232 41832 8232 0 _069_
rlabel metal2 42560 6664 42560 6664 0 _070_
rlabel metal2 43008 8344 43008 8344 0 _071_
rlabel metal2 41664 10808 41664 10808 0 _072_
rlabel metal3 41272 12040 41272 12040 0 _073_
rlabel metal2 37688 14112 37688 14112 0 _074_
rlabel metal3 39480 13944 39480 13944 0 _075_
rlabel metal3 39984 15512 39984 15512 0 _076_
rlabel metal2 38248 14336 38248 14336 0 _077_
rlabel metal3 28728 7448 28728 7448 0 clknet_0_clock
rlabel metal2 6216 7392 6216 7392 0 clknet_2_0__leaf_clock
rlabel metal2 6832 10472 6832 10472 0 clknet_2_1__leaf_clock
rlabel metal2 29736 5040 29736 5040 0 clknet_2_2__leaf_clock
rlabel metal3 24864 11368 24864 11368 0 clknet_2_3__leaf_clock
rlabel metal2 3080 4718 3080 4718 0 clock
rlabel metal3 48818 1624 48818 1624 0 clock_out
rlabel metal3 48650 3080 48650 3080 0 data_out[0]
rlabel metal2 47880 17976 47880 17976 0 data_out[10]
rlabel metal3 48650 19096 48650 19096 0 data_out[11]
rlabel metal3 48650 20552 48650 20552 0 data_out[12]
rlabel metal3 48650 22008 48650 22008 0 data_out[13]
rlabel metal3 48650 23464 48650 23464 0 data_out[14]
rlabel metal3 48650 24920 48650 24920 0 data_out[15]
rlabel metal3 48650 26376 48650 26376 0 data_out[16]
rlabel metal3 48706 27832 48706 27832 0 data_out[17]
rlabel metal3 48706 29288 48706 29288 0 data_out[18]
rlabel metal2 47880 30800 47880 30800 0 data_out[19]
rlabel metal3 49098 4536 49098 4536 0 data_out[1]
rlabel metal2 47880 32312 47880 32312 0 data_out[20]
rlabel metal2 47880 33824 47880 33824 0 data_out[21]
rlabel metal2 47880 35448 47880 35448 0 data_out[22]
rlabel metal2 47880 36848 47880 36848 0 data_out[23]
rlabel metal3 48720 38696 48720 38696 0 data_out[24]
rlabel metal3 48650 39480 48650 39480 0 data_out[25]
rlabel metal3 48650 40936 48650 40936 0 data_out[26]
rlabel metal3 48650 42392 48650 42392 0 data_out[27]
rlabel metal3 48650 43848 48650 43848 0 data_out[28]
rlabel metal3 48650 45304 48650 45304 0 data_out[29]
rlabel metal3 48650 5992 48650 5992 0 data_out[2]
rlabel metal2 47880 45864 47880 45864 0 data_out[30]
rlabel metal2 46088 47096 46088 47096 0 data_out[31]
rlabel metal3 48650 7448 48650 7448 0 data_out[3]
rlabel metal3 48706 8904 48706 8904 0 data_out[4]
rlabel metal2 47880 10416 47880 10416 0 data_out[5]
rlabel metal2 47880 11928 47880 11928 0 data_out[6]
rlabel metal2 47880 13552 47880 13552 0 data_out[7]
rlabel metal3 48706 14728 48706 14728 0 data_out[8]
rlabel metal3 48664 16856 48664 16856 0 data_out[9]
rlabel metal3 1302 40488 1302 40488 0 miso
rlabel metal2 1848 15568 1848 15568 0 mosi
rlabel metal3 6664 7560 6664 7560 0 mosi_reg\[0\]
rlabel metal2 22904 6216 22904 6216 0 mosi_reg\[1\]
rlabel metal2 20328 6048 20328 6048 0 mosi_reg\[2\]
rlabel metal2 2968 9856 2968 9856 0 net1
rlabel metal2 28560 11928 28560 11928 0 net10
rlabel metal2 28784 5768 28784 5768 0 net11
rlabel metal2 20440 4312 20440 4312 0 net12
rlabel metal3 46032 28616 46032 28616 0 net13
rlabel metal2 46872 29344 46872 29344 0 net14
rlabel metal2 46424 30912 46424 30912 0 net15
rlabel metal3 38360 6552 38360 6552 0 net16
rlabel metal2 23688 16408 23688 16408 0 net17
rlabel metal2 46368 33992 46368 33992 0 net18
rlabel metal2 20552 16464 20552 16464 0 net19
rlabel metal2 2520 3304 2520 3304 0 net2
rlabel metal2 22456 15904 22456 15904 0 net20
rlabel metal2 46872 38752 46872 38752 0 net21
rlabel metal3 46144 31080 46144 31080 0 net22
rlabel metal2 46256 40936 46256 40936 0 net23
rlabel metal2 46312 42224 46312 42224 0 net24
rlabel metal2 46592 44296 46592 44296 0 net25
rlabel metal2 45864 45360 45864 45360 0 net26
rlabel metal2 37688 5264 37688 5264 0 net27
rlabel metal2 46424 44744 46424 44744 0 net28
rlabel metal2 45080 45752 45080 45752 0 net29
rlabel metal2 2520 28392 2520 28392 0 net3
rlabel metal2 46312 7952 46312 7952 0 net30
rlabel metal2 38360 6272 38360 6272 0 net31
rlabel metal2 38584 7896 38584 7896 0 net32
rlabel metal3 39816 10472 39816 10472 0 net33
rlabel metal3 46592 13720 46592 13720 0 net34
rlabel metal2 38584 13104 38584 13104 0 net35
rlabel metal2 36792 14672 36792 14672 0 net36
rlabel metal2 3080 41048 3080 41048 0 net37
rlabel metal2 8568 1862 8568 1862 0 net38
rlabel metal2 14056 1862 14056 1862 0 net39
rlabel metal3 47488 4536 47488 4536 0 net4
rlabel metal2 19544 1862 19544 1862 0 net40
rlabel metal2 24696 3304 24696 3304 0 net41
rlabel metal3 1134 22008 1134 22008 0 net42
rlabel metal2 1848 9352 1848 9352 0 net43
rlabel metal3 1134 34328 1134 34328 0 net44
rlabel metal2 1848 46256 1848 46256 0 net45
rlabel metal2 32536 4984 32536 4984 0 net5
rlabel metal2 37912 14280 37912 14280 0 net6
rlabel metal2 36456 13552 36456 13552 0 net7
rlabel metal2 28840 10248 28840 10248 0 net8
rlabel metal1 29568 3752 29568 3752 0 net9
rlabel metal3 1134 3528 1134 3528 0 sclk
rlabel metal2 4200 8372 4200 8372 0 sclk_reg\[0\]
rlabel metal2 2072 8232 2072 8232 0 sclk_reg\[1\]
rlabel metal2 12936 15288 12936 15288 0 sclk_reg\[2\]
rlabel metal3 1134 28056 1134 28056 0 ss_n
rlabel metal2 6328 10080 6328 10080 0 ss_n_reg\[0\]
rlabel metal2 13048 7504 13048 7504 0 ss_n_reg\[1\]
rlabel metal2 16632 6720 16632 6720 0 ss_n_reg\[2\]
<< properties >>
string FIXED_BBOX 0 0 50000 50000
<< end >>

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO driver_core
  CLASS BLOCK ;
  FOREIGN driver_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 720.000 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 687.680 0.000 688.240 4.000 ;
    END
  END clock
  PIN clock_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 706.720 0.000 707.280 4.000 ;
    END
  END clock_a
  PIN col_select_a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 573.440 0.000 574.000 4.000 ;
    END
  END col_select_a[0]
  PIN col_select_a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 592.480 0.000 593.040 4.000 ;
    END
  END col_select_a[1]
  PIN col_select_a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 611.520 0.000 612.080 4.000 ;
    END
  END col_select_a[2]
  PIN col_select_a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 630.560 0.000 631.120 4.000 ;
    END
  END col_select_a[3]
  PIN col_select_a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 649.600 0.000 650.160 4.000 ;
    END
  END col_select_a[4]
  PIN col_select_a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 668.640 0.000 669.200 4.000 ;
    END
  END col_select_a[5]
  PIN data_in_a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 59.360 0.000 59.920 4.000 ;
    END
  END data_in_a[0]
  PIN data_in_a[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 249.760 0.000 250.320 4.000 ;
    END
  END data_in_a[10]
  PIN data_in_a[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 268.800 0.000 269.360 4.000 ;
    END
  END data_in_a[11]
  PIN data_in_a[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 287.840 0.000 288.400 4.000 ;
    END
  END data_in_a[12]
  PIN data_in_a[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 306.880 0.000 307.440 4.000 ;
    END
  END data_in_a[13]
  PIN data_in_a[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 325.920 0.000 326.480 4.000 ;
    END
  END data_in_a[14]
  PIN data_in_a[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 344.960 0.000 345.520 4.000 ;
    END
  END data_in_a[15]
  PIN data_in_a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 78.400 0.000 78.960 4.000 ;
    END
  END data_in_a[1]
  PIN data_in_a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 0.000 98.000 4.000 ;
    END
  END data_in_a[2]
  PIN data_in_a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 116.480 0.000 117.040 4.000 ;
    END
  END data_in_a[3]
  PIN data_in_a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 135.520 0.000 136.080 4.000 ;
    END
  END data_in_a[4]
  PIN data_in_a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 154.560 0.000 155.120 4.000 ;
    END
  END data_in_a[5]
  PIN data_in_a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 173.600 0.000 174.160 4.000 ;
    END
  END data_in_a[6]
  PIN data_in_a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 192.640 0.000 193.200 4.000 ;
    END
  END data_in_a[7]
  PIN data_in_a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 211.680 0.000 212.240 4.000 ;
    END
  END data_in_a[8]
  PIN data_in_a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 230.720 0.000 231.280 4.000 ;
    END
  END data_in_a[9]
  PIN driver_io[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 21.280 0.000 21.840 4.000 ;
    END
  END driver_io[0]
  PIN driver_io[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 40.320 0.000 40.880 4.000 ;
    END
  END driver_io[1]
  PIN inverter_select_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 878.080 0.000 878.640 4.000 ;
    END
  END inverter_select_a
  PIN mem_address_a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 364.000 0.000 364.560 4.000 ;
    END
  END mem_address_a[0]
  PIN mem_address_a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 383.040 0.000 383.600 4.000 ;
    END
  END mem_address_a[1]
  PIN mem_address_a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 402.080 0.000 402.640 4.000 ;
    END
  END mem_address_a[2]
  PIN mem_address_a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 421.120 0.000 421.680 4.000 ;
    END
  END mem_address_a[3]
  PIN mem_address_a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 440.160 0.000 440.720 4.000 ;
    END
  END mem_address_a[4]
  PIN mem_address_a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 459.200 0.000 459.760 4.000 ;
    END
  END mem_address_a[5]
  PIN mem_address_a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 478.240 0.000 478.800 4.000 ;
    END
  END mem_address_a[6]
  PIN mem_address_a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 497.280 0.000 497.840 4.000 ;
    END
  END mem_address_a[7]
  PIN mem_address_a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 516.320 0.000 516.880 4.000 ;
    END
  END mem_address_a[8]
  PIN mem_address_a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 535.360 0.000 535.920 4.000 ;
    END
  END mem_address_a[9]
  PIN mem_write_n_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 554.400 0.000 554.960 4.000 ;
    END
  END mem_write_n_a
  PIN output_active_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 859.040 0.000 859.600 4.000 ;
    END
  END output_active_a
  PIN row_col_select_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 840.000 0.000 840.560 4.000 ;
    END
  END row_col_select_a
  PIN row_select_a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 725.760 0.000 726.320 4.000 ;
    END
  END row_select_a[0]
  PIN row_select_a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 744.800 0.000 745.360 4.000 ;
    END
  END row_select_a[1]
  PIN row_select_a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 763.840 0.000 764.400 4.000 ;
    END
  END row_select_a[2]
  PIN row_select_a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 782.880 0.000 783.440 4.000 ;
    END
  END row_select_a[3]
  PIN row_select_a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 801.920 0.000 802.480 4.000 ;
    END
  END row_select_a[4]
  PIN row_select_a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 820.960 0.000 821.520 4.000 ;
    END
  END row_select_a[5]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 10.920 15.380 12.520 701.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 100.920 15.380 102.520 701.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 190.920 15.380 192.520 701.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 280.920 15.380 282.520 701.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 370.920 15.380 372.520 701.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 460.920 15.380 462.520 701.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 550.920 15.380 552.520 701.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 640.920 15.380 642.520 701.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 730.920 15.380 732.520 701.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 820.920 15.380 822.520 701.980 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 55.920 15.380 57.520 701.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 145.920 15.380 147.520 701.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 235.920 15.380 237.520 701.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 325.920 15.380 327.520 701.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 415.920 15.380 417.520 701.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 505.920 15.380 507.520 701.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 595.920 15.380 597.520 701.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 685.920 15.380 687.520 701.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 775.920 15.380 777.520 701.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 865.920 15.380 867.520 701.980 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 893.200 701.980 ;
      LAYER Metal2 ;
        RECT 7.980 4.300 894.740 701.870 ;
        RECT 7.980 2.890 20.980 4.300 ;
        RECT 22.140 2.890 40.020 4.300 ;
        RECT 41.180 2.890 59.060 4.300 ;
        RECT 60.220 2.890 78.100 4.300 ;
        RECT 79.260 2.890 97.140 4.300 ;
        RECT 98.300 2.890 116.180 4.300 ;
        RECT 117.340 2.890 135.220 4.300 ;
        RECT 136.380 2.890 154.260 4.300 ;
        RECT 155.420 2.890 173.300 4.300 ;
        RECT 174.460 2.890 192.340 4.300 ;
        RECT 193.500 2.890 211.380 4.300 ;
        RECT 212.540 2.890 230.420 4.300 ;
        RECT 231.580 2.890 249.460 4.300 ;
        RECT 250.620 2.890 268.500 4.300 ;
        RECT 269.660 2.890 287.540 4.300 ;
        RECT 288.700 2.890 306.580 4.300 ;
        RECT 307.740 2.890 325.620 4.300 ;
        RECT 326.780 2.890 344.660 4.300 ;
        RECT 345.820 2.890 363.700 4.300 ;
        RECT 364.860 2.890 382.740 4.300 ;
        RECT 383.900 2.890 401.780 4.300 ;
        RECT 402.940 2.890 420.820 4.300 ;
        RECT 421.980 2.890 439.860 4.300 ;
        RECT 441.020 2.890 458.900 4.300 ;
        RECT 460.060 2.890 477.940 4.300 ;
        RECT 479.100 2.890 496.980 4.300 ;
        RECT 498.140 2.890 516.020 4.300 ;
        RECT 517.180 2.890 535.060 4.300 ;
        RECT 536.220 2.890 554.100 4.300 ;
        RECT 555.260 2.890 573.140 4.300 ;
        RECT 574.300 2.890 592.180 4.300 ;
        RECT 593.340 2.890 611.220 4.300 ;
        RECT 612.380 2.890 630.260 4.300 ;
        RECT 631.420 2.890 649.300 4.300 ;
        RECT 650.460 2.890 668.340 4.300 ;
        RECT 669.500 2.890 687.380 4.300 ;
        RECT 688.540 2.890 706.420 4.300 ;
        RECT 707.580 2.890 725.460 4.300 ;
        RECT 726.620 2.890 744.500 4.300 ;
        RECT 745.660 2.890 763.540 4.300 ;
        RECT 764.700 2.890 782.580 4.300 ;
        RECT 783.740 2.890 801.620 4.300 ;
        RECT 802.780 2.890 820.660 4.300 ;
        RECT 821.820 2.890 839.700 4.300 ;
        RECT 840.860 2.890 858.740 4.300 ;
        RECT 859.900 2.890 877.780 4.300 ;
        RECT 878.940 2.890 894.740 4.300 ;
      LAYER Metal3 ;
        RECT 7.930 2.940 894.790 701.820 ;
      LAYER Metal4 ;
        RECT 55.020 15.080 55.620 681.430 ;
        RECT 57.820 15.080 100.620 681.430 ;
        RECT 102.820 15.080 145.620 681.430 ;
        RECT 147.820 15.080 190.620 681.430 ;
        RECT 192.820 15.080 235.620 681.430 ;
        RECT 237.820 15.080 280.620 681.430 ;
        RECT 282.820 15.080 325.620 681.430 ;
        RECT 327.820 15.080 370.620 681.430 ;
        RECT 372.820 15.080 415.620 681.430 ;
        RECT 417.820 15.080 460.620 681.430 ;
        RECT 462.820 15.080 505.620 681.430 ;
        RECT 507.820 15.080 550.620 681.430 ;
        RECT 552.820 15.080 595.620 681.430 ;
        RECT 597.820 15.080 640.620 681.430 ;
        RECT 642.820 15.080 685.620 681.430 ;
        RECT 687.820 15.080 730.620 681.430 ;
        RECT 732.820 15.080 775.620 681.430 ;
        RECT 777.820 15.080 820.620 681.430 ;
        RECT 822.820 15.080 865.620 681.430 ;
        RECT 867.820 15.080 884.660 681.430 ;
        RECT 55.020 4.570 884.660 15.080 ;
  END
END driver_core
END LIBRARY


magic
tech gf180mcuC
magscale 1 5
timestamp 1670293816
<< obsm1 >>
rect 672 1538 79296 21489
<< metal2 >>
rect 616 22600 672 23000
rect 1288 22600 1344 23000
rect 1960 22600 2016 23000
rect 2632 22600 2688 23000
rect 3304 22600 3360 23000
rect 3976 22600 4032 23000
rect 4648 22600 4704 23000
rect 5320 22600 5376 23000
rect 5992 22600 6048 23000
rect 6664 22600 6720 23000
rect 7336 22600 7392 23000
rect 8008 22600 8064 23000
rect 8680 22600 8736 23000
rect 9352 22600 9408 23000
rect 10024 22600 10080 23000
rect 10696 22600 10752 23000
rect 11368 22600 11424 23000
rect 12040 22600 12096 23000
rect 12712 22600 12768 23000
rect 13384 22600 13440 23000
rect 14056 22600 14112 23000
rect 14728 22600 14784 23000
rect 15400 22600 15456 23000
rect 16072 22600 16128 23000
rect 16744 22600 16800 23000
rect 17416 22600 17472 23000
rect 18088 22600 18144 23000
rect 18760 22600 18816 23000
rect 19432 22600 19488 23000
rect 20104 22600 20160 23000
rect 20776 22600 20832 23000
rect 21448 22600 21504 23000
rect 22120 22600 22176 23000
rect 22792 22600 22848 23000
rect 23464 22600 23520 23000
rect 24136 22600 24192 23000
rect 24808 22600 24864 23000
rect 25480 22600 25536 23000
rect 26152 22600 26208 23000
rect 26824 22600 26880 23000
rect 27496 22600 27552 23000
rect 28168 22600 28224 23000
rect 28840 22600 28896 23000
rect 29512 22600 29568 23000
rect 30184 22600 30240 23000
rect 30856 22600 30912 23000
rect 31528 22600 31584 23000
rect 32200 22600 32256 23000
rect 32872 22600 32928 23000
rect 33544 22600 33600 23000
rect 34216 22600 34272 23000
rect 34888 22600 34944 23000
rect 35560 22600 35616 23000
rect 36232 22600 36288 23000
rect 36904 22600 36960 23000
rect 37576 22600 37632 23000
rect 38248 22600 38304 23000
rect 38920 22600 38976 23000
rect 39592 22600 39648 23000
rect 40264 22600 40320 23000
rect 40936 22600 40992 23000
rect 41608 22600 41664 23000
rect 42280 22600 42336 23000
rect 42952 22600 43008 23000
rect 43624 22600 43680 23000
rect 44296 22600 44352 23000
rect 44968 22600 45024 23000
rect 45640 22600 45696 23000
rect 46312 22600 46368 23000
rect 46984 22600 47040 23000
rect 47656 22600 47712 23000
rect 48328 22600 48384 23000
rect 49000 22600 49056 23000
rect 49672 22600 49728 23000
rect 50344 22600 50400 23000
rect 51016 22600 51072 23000
rect 51688 22600 51744 23000
rect 52360 22600 52416 23000
rect 53032 22600 53088 23000
rect 53704 22600 53760 23000
rect 54376 22600 54432 23000
rect 55048 22600 55104 23000
rect 55720 22600 55776 23000
rect 56392 22600 56448 23000
rect 57064 22600 57120 23000
rect 57736 22600 57792 23000
rect 58408 22600 58464 23000
rect 59080 22600 59136 23000
rect 59752 22600 59808 23000
rect 60424 22600 60480 23000
rect 61096 22600 61152 23000
rect 61768 22600 61824 23000
rect 62440 22600 62496 23000
rect 63112 22600 63168 23000
rect 63784 22600 63840 23000
rect 64456 22600 64512 23000
rect 65128 22600 65184 23000
rect 65800 22600 65856 23000
rect 66472 22600 66528 23000
rect 67144 22600 67200 23000
rect 67816 22600 67872 23000
rect 68488 22600 68544 23000
rect 69160 22600 69216 23000
rect 69832 22600 69888 23000
rect 70504 22600 70560 23000
rect 71176 22600 71232 23000
rect 71848 22600 71904 23000
rect 72520 22600 72576 23000
rect 73192 22600 73248 23000
rect 73864 22600 73920 23000
rect 74536 22600 74592 23000
rect 75208 22600 75264 23000
rect 75880 22600 75936 23000
rect 76552 22600 76608 23000
rect 77224 22600 77280 23000
rect 77896 22600 77952 23000
rect 78568 22600 78624 23000
rect 79240 22600 79296 23000
rect 2296 0 2352 400
rect 3472 0 3528 400
rect 4648 0 4704 400
rect 5824 0 5880 400
rect 7000 0 7056 400
rect 8176 0 8232 400
rect 9352 0 9408 400
rect 10528 0 10584 400
rect 11704 0 11760 400
rect 12880 0 12936 400
rect 14056 0 14112 400
rect 15232 0 15288 400
rect 16408 0 16464 400
rect 17584 0 17640 400
rect 18760 0 18816 400
rect 19936 0 19992 400
rect 21112 0 21168 400
rect 22288 0 22344 400
rect 23464 0 23520 400
rect 24640 0 24696 400
rect 25816 0 25872 400
rect 26992 0 27048 400
rect 28168 0 28224 400
rect 29344 0 29400 400
rect 30520 0 30576 400
rect 31696 0 31752 400
rect 32872 0 32928 400
rect 34048 0 34104 400
rect 35224 0 35280 400
rect 36400 0 36456 400
rect 37576 0 37632 400
rect 38752 0 38808 400
rect 39928 0 39984 400
rect 41104 0 41160 400
rect 42280 0 42336 400
rect 43456 0 43512 400
rect 44632 0 44688 400
rect 45808 0 45864 400
rect 46984 0 47040 400
rect 48160 0 48216 400
rect 49336 0 49392 400
rect 50512 0 50568 400
rect 51688 0 51744 400
rect 52864 0 52920 400
rect 54040 0 54096 400
rect 55216 0 55272 400
rect 56392 0 56448 400
rect 57568 0 57624 400
rect 58744 0 58800 400
rect 59920 0 59976 400
rect 61096 0 61152 400
rect 62272 0 62328 400
rect 63448 0 63504 400
rect 64624 0 64680 400
rect 65800 0 65856 400
rect 66976 0 67032 400
rect 68152 0 68208 400
rect 69328 0 69384 400
rect 70504 0 70560 400
rect 71680 0 71736 400
rect 72856 0 72912 400
rect 74032 0 74088 400
rect 75208 0 75264 400
rect 76384 0 76440 400
rect 77560 0 77616 400
<< obsm2 >>
rect 702 22570 1258 22666
rect 1374 22570 1930 22666
rect 2046 22570 2602 22666
rect 2718 22570 3274 22666
rect 3390 22570 3946 22666
rect 4062 22570 4618 22666
rect 4734 22570 5290 22666
rect 5406 22570 5962 22666
rect 6078 22570 6634 22666
rect 6750 22570 7306 22666
rect 7422 22570 7978 22666
rect 8094 22570 8650 22666
rect 8766 22570 9322 22666
rect 9438 22570 9994 22666
rect 10110 22570 10666 22666
rect 10782 22570 11338 22666
rect 11454 22570 12010 22666
rect 12126 22570 12682 22666
rect 12798 22570 13354 22666
rect 13470 22570 14026 22666
rect 14142 22570 14698 22666
rect 14814 22570 15370 22666
rect 15486 22570 16042 22666
rect 16158 22570 16714 22666
rect 16830 22570 17386 22666
rect 17502 22570 18058 22666
rect 18174 22570 18730 22666
rect 18846 22570 19402 22666
rect 19518 22570 20074 22666
rect 20190 22570 20746 22666
rect 20862 22570 21418 22666
rect 21534 22570 22090 22666
rect 22206 22570 22762 22666
rect 22878 22570 23434 22666
rect 23550 22570 24106 22666
rect 24222 22570 24778 22666
rect 24894 22570 25450 22666
rect 25566 22570 26122 22666
rect 26238 22570 26794 22666
rect 26910 22570 27466 22666
rect 27582 22570 28138 22666
rect 28254 22570 28810 22666
rect 28926 22570 29482 22666
rect 29598 22570 30154 22666
rect 30270 22570 30826 22666
rect 30942 22570 31498 22666
rect 31614 22570 32170 22666
rect 32286 22570 32842 22666
rect 32958 22570 33514 22666
rect 33630 22570 34186 22666
rect 34302 22570 34858 22666
rect 34974 22570 35530 22666
rect 35646 22570 36202 22666
rect 36318 22570 36874 22666
rect 36990 22570 37546 22666
rect 37662 22570 38218 22666
rect 38334 22570 38890 22666
rect 39006 22570 39562 22666
rect 39678 22570 40234 22666
rect 40350 22570 40906 22666
rect 41022 22570 41578 22666
rect 41694 22570 42250 22666
rect 42366 22570 42922 22666
rect 43038 22570 43594 22666
rect 43710 22570 44266 22666
rect 44382 22570 44938 22666
rect 45054 22570 45610 22666
rect 45726 22570 46282 22666
rect 46398 22570 46954 22666
rect 47070 22570 47626 22666
rect 47742 22570 48298 22666
rect 48414 22570 48970 22666
rect 49086 22570 49642 22666
rect 49758 22570 50314 22666
rect 50430 22570 50986 22666
rect 51102 22570 51658 22666
rect 51774 22570 52330 22666
rect 52446 22570 53002 22666
rect 53118 22570 53674 22666
rect 53790 22570 54346 22666
rect 54462 22570 55018 22666
rect 55134 22570 55690 22666
rect 55806 22570 56362 22666
rect 56478 22570 57034 22666
rect 57150 22570 57706 22666
rect 57822 22570 58378 22666
rect 58494 22570 59050 22666
rect 59166 22570 59722 22666
rect 59838 22570 60394 22666
rect 60510 22570 61066 22666
rect 61182 22570 61738 22666
rect 61854 22570 62410 22666
rect 62526 22570 63082 22666
rect 63198 22570 63754 22666
rect 63870 22570 64426 22666
rect 64542 22570 65098 22666
rect 65214 22570 65770 22666
rect 65886 22570 66442 22666
rect 66558 22570 67114 22666
rect 67230 22570 67786 22666
rect 67902 22570 68458 22666
rect 68574 22570 69130 22666
rect 69246 22570 69802 22666
rect 69918 22570 70474 22666
rect 70590 22570 71146 22666
rect 71262 22570 71818 22666
rect 71934 22570 72490 22666
rect 72606 22570 73162 22666
rect 73278 22570 73834 22666
rect 73950 22570 74506 22666
rect 74622 22570 75178 22666
rect 75294 22570 75850 22666
rect 75966 22570 76522 22666
rect 76638 22570 77194 22666
rect 77310 22570 77866 22666
rect 77982 22570 78538 22666
rect 78654 22570 79210 22666
rect 79326 22570 79394 22666
rect 630 430 79394 22570
rect 630 350 2266 430
rect 2382 350 3442 430
rect 3558 350 4618 430
rect 4734 350 5794 430
rect 5910 350 6970 430
rect 7086 350 8146 430
rect 8262 350 9322 430
rect 9438 350 10498 430
rect 10614 350 11674 430
rect 11790 350 12850 430
rect 12966 350 14026 430
rect 14142 350 15202 430
rect 15318 350 16378 430
rect 16494 350 17554 430
rect 17670 350 18730 430
rect 18846 350 19906 430
rect 20022 350 21082 430
rect 21198 350 22258 430
rect 22374 350 23434 430
rect 23550 350 24610 430
rect 24726 350 25786 430
rect 25902 350 26962 430
rect 27078 350 28138 430
rect 28254 350 29314 430
rect 29430 350 30490 430
rect 30606 350 31666 430
rect 31782 350 32842 430
rect 32958 350 34018 430
rect 34134 350 35194 430
rect 35310 350 36370 430
rect 36486 350 37546 430
rect 37662 350 38722 430
rect 38838 350 39898 430
rect 40014 350 41074 430
rect 41190 350 42250 430
rect 42366 350 43426 430
rect 43542 350 44602 430
rect 44718 350 45778 430
rect 45894 350 46954 430
rect 47070 350 48130 430
rect 48246 350 49306 430
rect 49422 350 50482 430
rect 50598 350 51658 430
rect 51774 350 52834 430
rect 52950 350 54010 430
rect 54126 350 55186 430
rect 55302 350 56362 430
rect 56478 350 57538 430
rect 57654 350 58714 430
rect 58830 350 59890 430
rect 60006 350 61066 430
rect 61182 350 62242 430
rect 62358 350 63418 430
rect 63534 350 64594 430
rect 64710 350 65770 430
rect 65886 350 66946 430
rect 67062 350 68122 430
rect 68238 350 69298 430
rect 69414 350 70474 430
rect 70590 350 71650 430
rect 71766 350 72826 430
rect 72942 350 74002 430
rect 74118 350 75178 430
rect 75294 350 76354 430
rect 76470 350 77530 430
rect 77646 350 79394 430
<< metal3 >>
rect 0 22176 400 22232
rect 0 21504 400 21560
rect 0 20832 400 20888
rect 0 20160 400 20216
rect 0 19488 400 19544
rect 0 18816 400 18872
rect 0 18144 400 18200
rect 0 17472 400 17528
rect 0 16800 400 16856
rect 0 16128 400 16184
rect 0 15456 400 15512
rect 0 14784 400 14840
rect 0 14112 400 14168
rect 0 13440 400 13496
rect 0 12768 400 12824
rect 0 12096 400 12152
rect 0 11424 400 11480
rect 0 10752 400 10808
rect 0 10080 400 10136
rect 0 9408 400 9464
rect 0 8736 400 8792
rect 0 8064 400 8120
rect 0 7392 400 7448
rect 0 6720 400 6776
rect 0 6048 400 6104
rect 0 5376 400 5432
rect 0 4704 400 4760
rect 0 4032 400 4088
rect 0 3360 400 3416
rect 0 2688 400 2744
rect 0 2016 400 2072
rect 0 1344 400 1400
rect 0 672 400 728
<< obsm3 >>
rect 350 22262 79399 22610
rect 430 22146 79399 22262
rect 350 21590 79399 22146
rect 430 21474 79399 21590
rect 350 20918 79399 21474
rect 430 20802 79399 20918
rect 350 20246 79399 20802
rect 430 20130 79399 20246
rect 350 19574 79399 20130
rect 430 19458 79399 19574
rect 350 18902 79399 19458
rect 430 18786 79399 18902
rect 350 18230 79399 18786
rect 430 18114 79399 18230
rect 350 17558 79399 18114
rect 430 17442 79399 17558
rect 350 16886 79399 17442
rect 430 16770 79399 16886
rect 350 16214 79399 16770
rect 430 16098 79399 16214
rect 350 15542 79399 16098
rect 430 15426 79399 15542
rect 350 14870 79399 15426
rect 430 14754 79399 14870
rect 350 14198 79399 14754
rect 430 14082 79399 14198
rect 350 13526 79399 14082
rect 430 13410 79399 13526
rect 350 12854 79399 13410
rect 430 12738 79399 12854
rect 350 12182 79399 12738
rect 430 12066 79399 12182
rect 350 11510 79399 12066
rect 430 11394 79399 11510
rect 350 10838 79399 11394
rect 430 10722 79399 10838
rect 350 10166 79399 10722
rect 430 10050 79399 10166
rect 350 9494 79399 10050
rect 430 9378 79399 9494
rect 350 8822 79399 9378
rect 430 8706 79399 8822
rect 350 8150 79399 8706
rect 430 8034 79399 8150
rect 350 7478 79399 8034
rect 430 7362 79399 7478
rect 350 6806 79399 7362
rect 430 6690 79399 6806
rect 350 6134 79399 6690
rect 430 6018 79399 6134
rect 350 5462 79399 6018
rect 430 5346 79399 5462
rect 350 4790 79399 5346
rect 430 4674 79399 4790
rect 350 4118 79399 4674
rect 430 4002 79399 4118
rect 350 3446 79399 4002
rect 430 3330 79399 3446
rect 350 2774 79399 3330
rect 430 2658 79399 2774
rect 350 2102 79399 2658
rect 430 1986 79399 2102
rect 350 1430 79399 1986
rect 430 1314 79399 1430
rect 350 758 79399 1314
rect 430 642 79399 758
rect 350 462 79399 642
<< metal4 >>
rect 2224 1538 2384 21198
rect 9904 1538 10064 21198
rect 17584 1538 17744 21198
rect 25264 1538 25424 21198
rect 32944 1538 33104 21198
rect 40624 1538 40784 21198
rect 48304 1538 48464 21198
rect 55984 1538 56144 21198
rect 63664 1538 63824 21198
rect 71344 1538 71504 21198
rect 79024 1538 79184 21198
<< obsm4 >>
rect 15302 4825 17554 19591
rect 17774 4825 25234 19591
rect 25454 4825 32914 19591
rect 33134 4825 40594 19591
rect 40814 4825 48274 19591
rect 48494 4825 55954 19591
rect 56174 4825 63634 19591
rect 63854 4825 71314 19591
rect 71534 4825 74802 19591
<< labels >>
rlabel metal2 s 77560 0 77616 400 6 clock
port 1 nsew signal input
rlabel metal2 s 22120 22600 22176 23000 6 clock_out[0]
port 2 nsew signal output
rlabel metal2 s 22792 22600 22848 23000 6 clock_out[1]
port 3 nsew signal output
rlabel metal2 s 23464 22600 23520 23000 6 clock_out[2]
port 4 nsew signal output
rlabel metal2 s 24136 22600 24192 23000 6 clock_out[3]
port 5 nsew signal output
rlabel metal2 s 24808 22600 24864 23000 6 clock_out[4]
port 6 nsew signal output
rlabel metal2 s 25480 22600 25536 23000 6 clock_out[5]
port 7 nsew signal output
rlabel metal2 s 26152 22600 26208 23000 6 clock_out[6]
port 8 nsew signal output
rlabel metal2 s 26824 22600 26880 23000 6 clock_out[7]
port 9 nsew signal output
rlabel metal2 s 27496 22600 27552 23000 6 clock_out[8]
port 10 nsew signal output
rlabel metal2 s 28168 22600 28224 23000 6 clock_out[9]
port 11 nsew signal output
rlabel metal2 s 40936 22600 40992 23000 6 col_select_left[0]
port 12 nsew signal output
rlabel metal2 s 41608 22600 41664 23000 6 col_select_left[1]
port 13 nsew signal output
rlabel metal2 s 42280 22600 42336 23000 6 col_select_left[2]
port 14 nsew signal output
rlabel metal2 s 42952 22600 43008 23000 6 col_select_left[3]
port 15 nsew signal output
rlabel metal2 s 43624 22600 43680 23000 6 col_select_left[4]
port 16 nsew signal output
rlabel metal2 s 44296 22600 44352 23000 6 col_select_left[5]
port 17 nsew signal output
rlabel metal2 s 36904 22600 36960 23000 6 col_select_right[0]
port 18 nsew signal output
rlabel metal2 s 37576 22600 37632 23000 6 col_select_right[1]
port 19 nsew signal output
rlabel metal2 s 38248 22600 38304 23000 6 col_select_right[2]
port 20 nsew signal output
rlabel metal2 s 38920 22600 38976 23000 6 col_select_right[3]
port 21 nsew signal output
rlabel metal2 s 39592 22600 39648 23000 6 col_select_right[4]
port 22 nsew signal output
rlabel metal2 s 40264 22600 40320 23000 6 col_select_right[5]
port 23 nsew signal output
rlabel metal2 s 55720 22600 55776 23000 6 data_out_left[0]
port 24 nsew signal output
rlabel metal2 s 62440 22600 62496 23000 6 data_out_left[10]
port 25 nsew signal output
rlabel metal2 s 63112 22600 63168 23000 6 data_out_left[11]
port 26 nsew signal output
rlabel metal2 s 63784 22600 63840 23000 6 data_out_left[12]
port 27 nsew signal output
rlabel metal2 s 64456 22600 64512 23000 6 data_out_left[13]
port 28 nsew signal output
rlabel metal2 s 65128 22600 65184 23000 6 data_out_left[14]
port 29 nsew signal output
rlabel metal2 s 65800 22600 65856 23000 6 data_out_left[15]
port 30 nsew signal output
rlabel metal2 s 56392 22600 56448 23000 6 data_out_left[1]
port 31 nsew signal output
rlabel metal2 s 57064 22600 57120 23000 6 data_out_left[2]
port 32 nsew signal output
rlabel metal2 s 57736 22600 57792 23000 6 data_out_left[3]
port 33 nsew signal output
rlabel metal2 s 58408 22600 58464 23000 6 data_out_left[4]
port 34 nsew signal output
rlabel metal2 s 59080 22600 59136 23000 6 data_out_left[5]
port 35 nsew signal output
rlabel metal2 s 59752 22600 59808 23000 6 data_out_left[6]
port 36 nsew signal output
rlabel metal2 s 60424 22600 60480 23000 6 data_out_left[7]
port 37 nsew signal output
rlabel metal2 s 61096 22600 61152 23000 6 data_out_left[8]
port 38 nsew signal output
rlabel metal2 s 61768 22600 61824 23000 6 data_out_left[9]
port 39 nsew signal output
rlabel metal2 s 44968 22600 45024 23000 6 data_out_right[0]
port 40 nsew signal output
rlabel metal2 s 51688 22600 51744 23000 6 data_out_right[10]
port 41 nsew signal output
rlabel metal2 s 52360 22600 52416 23000 6 data_out_right[11]
port 42 nsew signal output
rlabel metal2 s 53032 22600 53088 23000 6 data_out_right[12]
port 43 nsew signal output
rlabel metal2 s 53704 22600 53760 23000 6 data_out_right[13]
port 44 nsew signal output
rlabel metal2 s 54376 22600 54432 23000 6 data_out_right[14]
port 45 nsew signal output
rlabel metal2 s 55048 22600 55104 23000 6 data_out_right[15]
port 46 nsew signal output
rlabel metal2 s 45640 22600 45696 23000 6 data_out_right[1]
port 47 nsew signal output
rlabel metal2 s 46312 22600 46368 23000 6 data_out_right[2]
port 48 nsew signal output
rlabel metal2 s 46984 22600 47040 23000 6 data_out_right[3]
port 49 nsew signal output
rlabel metal2 s 47656 22600 47712 23000 6 data_out_right[4]
port 50 nsew signal output
rlabel metal2 s 48328 22600 48384 23000 6 data_out_right[5]
port 51 nsew signal output
rlabel metal2 s 49000 22600 49056 23000 6 data_out_right[6]
port 52 nsew signal output
rlabel metal2 s 49672 22600 49728 23000 6 data_out_right[7]
port 53 nsew signal output
rlabel metal2 s 50344 22600 50400 23000 6 data_out_right[8]
port 54 nsew signal output
rlabel metal2 s 51016 22600 51072 23000 6 data_out_right[9]
port 55 nsew signal output
rlabel metal2 s 73192 22600 73248 23000 6 inverter_select[0]
port 56 nsew signal output
rlabel metal2 s 73864 22600 73920 23000 6 inverter_select[1]
port 57 nsew signal output
rlabel metal2 s 74536 22600 74592 23000 6 inverter_select[2]
port 58 nsew signal output
rlabel metal2 s 75208 22600 75264 23000 6 inverter_select[3]
port 59 nsew signal output
rlabel metal2 s 75880 22600 75936 23000 6 inverter_select[4]
port 60 nsew signal output
rlabel metal2 s 76552 22600 76608 23000 6 inverter_select[5]
port 61 nsew signal output
rlabel metal2 s 77224 22600 77280 23000 6 inverter_select[6]
port 62 nsew signal output
rlabel metal2 s 77896 22600 77952 23000 6 inverter_select[7]
port 63 nsew signal output
rlabel metal2 s 78568 22600 78624 23000 6 inverter_select[8]
port 64 nsew signal output
rlabel metal2 s 79240 22600 79296 23000 6 inverter_select[9]
port 65 nsew signal output
rlabel metal2 s 7000 0 7056 400 6 io_control_trigger_in
port 66 nsew signal input
rlabel metal2 s 8176 0 8232 400 6 io_control_trigger_oeb
port 67 nsew signal output
rlabel metal2 s 11704 0 11760 400 6 io_driver_io_oeb[0]
port 68 nsew signal output
rlabel metal2 s 23464 0 23520 400 6 io_driver_io_oeb[10]
port 69 nsew signal output
rlabel metal2 s 24640 0 24696 400 6 io_driver_io_oeb[11]
port 70 nsew signal output
rlabel metal2 s 25816 0 25872 400 6 io_driver_io_oeb[12]
port 71 nsew signal output
rlabel metal2 s 26992 0 27048 400 6 io_driver_io_oeb[13]
port 72 nsew signal output
rlabel metal2 s 28168 0 28224 400 6 io_driver_io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 29344 0 29400 400 6 io_driver_io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 30520 0 30576 400 6 io_driver_io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 31696 0 31752 400 6 io_driver_io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 32872 0 32928 400 6 io_driver_io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 34048 0 34104 400 6 io_driver_io_oeb[19]
port 78 nsew signal output
rlabel metal2 s 12880 0 12936 400 6 io_driver_io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 14056 0 14112 400 6 io_driver_io_oeb[2]
port 80 nsew signal output
rlabel metal2 s 15232 0 15288 400 6 io_driver_io_oeb[3]
port 81 nsew signal output
rlabel metal2 s 16408 0 16464 400 6 io_driver_io_oeb[4]
port 82 nsew signal output
rlabel metal2 s 17584 0 17640 400 6 io_driver_io_oeb[5]
port 83 nsew signal output
rlabel metal2 s 18760 0 18816 400 6 io_driver_io_oeb[6]
port 84 nsew signal output
rlabel metal2 s 19936 0 19992 400 6 io_driver_io_oeb[7]
port 85 nsew signal output
rlabel metal2 s 21112 0 21168 400 6 io_driver_io_oeb[8]
port 86 nsew signal output
rlabel metal2 s 22288 0 22344 400 6 io_driver_io_oeb[9]
port 87 nsew signal output
rlabel metal2 s 4648 0 4704 400 6 io_latch_data_in
port 88 nsew signal input
rlabel metal2 s 5824 0 5880 400 6 io_latch_data_oeb
port 89 nsew signal output
rlabel metal2 s 2296 0 2352 400 6 io_reset_n_in
port 90 nsew signal input
rlabel metal2 s 3472 0 3528 400 6 io_reset_n_oeb
port 91 nsew signal output
rlabel metal2 s 10528 0 10584 400 6 io_update_cycle_complete_oeb
port 92 nsew signal output
rlabel metal2 s 9352 0 9408 400 6 io_update_cycle_complete_out
port 93 nsew signal output
rlabel metal2 s 56392 0 56448 400 6 la_data_in[0]
port 94 nsew signal input
rlabel metal2 s 68152 0 68208 400 6 la_data_in[10]
port 95 nsew signal input
rlabel metal2 s 69328 0 69384 400 6 la_data_in[11]
port 96 nsew signal input
rlabel metal2 s 70504 0 70560 400 6 la_data_in[12]
port 97 nsew signal input
rlabel metal2 s 71680 0 71736 400 6 la_data_in[13]
port 98 nsew signal input
rlabel metal2 s 72856 0 72912 400 6 la_data_in[14]
port 99 nsew signal input
rlabel metal2 s 74032 0 74088 400 6 la_data_in[15]
port 100 nsew signal input
rlabel metal2 s 75208 0 75264 400 6 la_data_in[16]
port 101 nsew signal input
rlabel metal2 s 76384 0 76440 400 6 la_data_in[17]
port 102 nsew signal input
rlabel metal2 s 57568 0 57624 400 6 la_data_in[1]
port 103 nsew signal input
rlabel metal2 s 58744 0 58800 400 6 la_data_in[2]
port 104 nsew signal input
rlabel metal2 s 59920 0 59976 400 6 la_data_in[3]
port 105 nsew signal input
rlabel metal2 s 61096 0 61152 400 6 la_data_in[4]
port 106 nsew signal input
rlabel metal2 s 62272 0 62328 400 6 la_data_in[5]
port 107 nsew signal input
rlabel metal2 s 63448 0 63504 400 6 la_data_in[6]
port 108 nsew signal input
rlabel metal2 s 64624 0 64680 400 6 la_data_in[7]
port 109 nsew signal input
rlabel metal2 s 65800 0 65856 400 6 la_data_in[8]
port 110 nsew signal input
rlabel metal2 s 66976 0 67032 400 6 la_data_in[9]
port 111 nsew signal input
rlabel metal2 s 35224 0 35280 400 6 la_oenb[0]
port 112 nsew signal input
rlabel metal2 s 46984 0 47040 400 6 la_oenb[10]
port 113 nsew signal input
rlabel metal2 s 48160 0 48216 400 6 la_oenb[11]
port 114 nsew signal input
rlabel metal2 s 49336 0 49392 400 6 la_oenb[12]
port 115 nsew signal input
rlabel metal2 s 50512 0 50568 400 6 la_oenb[13]
port 116 nsew signal input
rlabel metal2 s 51688 0 51744 400 6 la_oenb[14]
port 117 nsew signal input
rlabel metal2 s 52864 0 52920 400 6 la_oenb[15]
port 118 nsew signal input
rlabel metal2 s 54040 0 54096 400 6 la_oenb[16]
port 119 nsew signal input
rlabel metal2 s 55216 0 55272 400 6 la_oenb[17]
port 120 nsew signal input
rlabel metal2 s 36400 0 36456 400 6 la_oenb[1]
port 121 nsew signal input
rlabel metal2 s 37576 0 37632 400 6 la_oenb[2]
port 122 nsew signal input
rlabel metal2 s 38752 0 38808 400 6 la_oenb[3]
port 123 nsew signal input
rlabel metal2 s 39928 0 39984 400 6 la_oenb[4]
port 124 nsew signal input
rlabel metal2 s 41104 0 41160 400 6 la_oenb[5]
port 125 nsew signal input
rlabel metal2 s 42280 0 42336 400 6 la_oenb[6]
port 126 nsew signal input
rlabel metal2 s 43456 0 43512 400 6 la_oenb[7]
port 127 nsew signal input
rlabel metal2 s 44632 0 44688 400 6 la_oenb[8]
port 128 nsew signal input
rlabel metal2 s 45808 0 45864 400 6 la_oenb[9]
port 129 nsew signal input
rlabel metal2 s 8680 22600 8736 23000 6 mem_address_left[0]
port 130 nsew signal output
rlabel metal2 s 9352 22600 9408 23000 6 mem_address_left[1]
port 131 nsew signal output
rlabel metal2 s 10024 22600 10080 23000 6 mem_address_left[2]
port 132 nsew signal output
rlabel metal2 s 10696 22600 10752 23000 6 mem_address_left[3]
port 133 nsew signal output
rlabel metal2 s 11368 22600 11424 23000 6 mem_address_left[4]
port 134 nsew signal output
rlabel metal2 s 12040 22600 12096 23000 6 mem_address_left[5]
port 135 nsew signal output
rlabel metal2 s 12712 22600 12768 23000 6 mem_address_left[6]
port 136 nsew signal output
rlabel metal2 s 13384 22600 13440 23000 6 mem_address_left[7]
port 137 nsew signal output
rlabel metal2 s 14056 22600 14112 23000 6 mem_address_left[8]
port 138 nsew signal output
rlabel metal2 s 14728 22600 14784 23000 6 mem_address_left[9]
port 139 nsew signal output
rlabel metal2 s 1960 22600 2016 23000 6 mem_address_right[0]
port 140 nsew signal output
rlabel metal2 s 2632 22600 2688 23000 6 mem_address_right[1]
port 141 nsew signal output
rlabel metal2 s 3304 22600 3360 23000 6 mem_address_right[2]
port 142 nsew signal output
rlabel metal2 s 3976 22600 4032 23000 6 mem_address_right[3]
port 143 nsew signal output
rlabel metal2 s 4648 22600 4704 23000 6 mem_address_right[4]
port 144 nsew signal output
rlabel metal2 s 5320 22600 5376 23000 6 mem_address_right[5]
port 145 nsew signal output
rlabel metal2 s 5992 22600 6048 23000 6 mem_address_right[6]
port 146 nsew signal output
rlabel metal2 s 6664 22600 6720 23000 6 mem_address_right[7]
port 147 nsew signal output
rlabel metal2 s 7336 22600 7392 23000 6 mem_address_right[8]
port 148 nsew signal output
rlabel metal2 s 8008 22600 8064 23000 6 mem_address_right[9]
port 149 nsew signal output
rlabel metal2 s 15400 22600 15456 23000 6 mem_write_n[0]
port 150 nsew signal output
rlabel metal2 s 16072 22600 16128 23000 6 mem_write_n[1]
port 151 nsew signal output
rlabel metal2 s 16744 22600 16800 23000 6 mem_write_n[2]
port 152 nsew signal output
rlabel metal2 s 17416 22600 17472 23000 6 mem_write_n[3]
port 153 nsew signal output
rlabel metal2 s 18088 22600 18144 23000 6 mem_write_n[4]
port 154 nsew signal output
rlabel metal2 s 18760 22600 18816 23000 6 mem_write_n[5]
port 155 nsew signal output
rlabel metal2 s 19432 22600 19488 23000 6 mem_write_n[6]
port 156 nsew signal output
rlabel metal2 s 20104 22600 20160 23000 6 mem_write_n[7]
port 157 nsew signal output
rlabel metal2 s 20776 22600 20832 23000 6 mem_write_n[8]
port 158 nsew signal output
rlabel metal2 s 21448 22600 21504 23000 6 mem_write_n[9]
port 159 nsew signal output
rlabel metal2 s 1288 22600 1344 23000 6 output_active_left
port 160 nsew signal output
rlabel metal2 s 616 22600 672 23000 6 output_active_right
port 161 nsew signal output
rlabel metal2 s 66472 22600 66528 23000 6 row_col_select[0]
port 162 nsew signal output
rlabel metal2 s 67144 22600 67200 23000 6 row_col_select[1]
port 163 nsew signal output
rlabel metal2 s 67816 22600 67872 23000 6 row_col_select[2]
port 164 nsew signal output
rlabel metal2 s 68488 22600 68544 23000 6 row_col_select[3]
port 165 nsew signal output
rlabel metal2 s 69160 22600 69216 23000 6 row_col_select[4]
port 166 nsew signal output
rlabel metal2 s 69832 22600 69888 23000 6 row_col_select[5]
port 167 nsew signal output
rlabel metal2 s 70504 22600 70560 23000 6 row_col_select[6]
port 168 nsew signal output
rlabel metal2 s 71176 22600 71232 23000 6 row_col_select[7]
port 169 nsew signal output
rlabel metal2 s 71848 22600 71904 23000 6 row_col_select[8]
port 170 nsew signal output
rlabel metal2 s 72520 22600 72576 23000 6 row_col_select[9]
port 171 nsew signal output
rlabel metal2 s 32872 22600 32928 23000 6 row_select_left[0]
port 172 nsew signal output
rlabel metal2 s 33544 22600 33600 23000 6 row_select_left[1]
port 173 nsew signal output
rlabel metal2 s 34216 22600 34272 23000 6 row_select_left[2]
port 174 nsew signal output
rlabel metal2 s 34888 22600 34944 23000 6 row_select_left[3]
port 175 nsew signal output
rlabel metal2 s 35560 22600 35616 23000 6 row_select_left[4]
port 176 nsew signal output
rlabel metal2 s 36232 22600 36288 23000 6 row_select_left[5]
port 177 nsew signal output
rlabel metal2 s 28840 22600 28896 23000 6 row_select_right[0]
port 178 nsew signal output
rlabel metal2 s 29512 22600 29568 23000 6 row_select_right[1]
port 179 nsew signal output
rlabel metal2 s 30184 22600 30240 23000 6 row_select_right[2]
port 180 nsew signal output
rlabel metal2 s 30856 22600 30912 23000 6 row_select_right[3]
port 181 nsew signal output
rlabel metal2 s 31528 22600 31584 23000 6 row_select_right[4]
port 182 nsew signal output
rlabel metal2 s 32200 22600 32256 23000 6 row_select_right[5]
port 183 nsew signal output
rlabel metal3 s 0 1344 400 1400 6 spi_data[0]
port 184 nsew signal input
rlabel metal3 s 0 8064 400 8120 6 spi_data[10]
port 185 nsew signal input
rlabel metal3 s 0 8736 400 8792 6 spi_data[11]
port 186 nsew signal input
rlabel metal3 s 0 9408 400 9464 6 spi_data[12]
port 187 nsew signal input
rlabel metal3 s 0 10080 400 10136 6 spi_data[13]
port 188 nsew signal input
rlabel metal3 s 0 10752 400 10808 6 spi_data[14]
port 189 nsew signal input
rlabel metal3 s 0 11424 400 11480 6 spi_data[15]
port 190 nsew signal input
rlabel metal3 s 0 12096 400 12152 6 spi_data[16]
port 191 nsew signal input
rlabel metal3 s 0 12768 400 12824 6 spi_data[17]
port 192 nsew signal input
rlabel metal3 s 0 13440 400 13496 6 spi_data[18]
port 193 nsew signal input
rlabel metal3 s 0 14112 400 14168 6 spi_data[19]
port 194 nsew signal input
rlabel metal3 s 0 2016 400 2072 6 spi_data[1]
port 195 nsew signal input
rlabel metal3 s 0 14784 400 14840 6 spi_data[20]
port 196 nsew signal input
rlabel metal3 s 0 15456 400 15512 6 spi_data[21]
port 197 nsew signal input
rlabel metal3 s 0 16128 400 16184 6 spi_data[22]
port 198 nsew signal input
rlabel metal3 s 0 16800 400 16856 6 spi_data[23]
port 199 nsew signal input
rlabel metal3 s 0 17472 400 17528 6 spi_data[24]
port 200 nsew signal input
rlabel metal3 s 0 18144 400 18200 6 spi_data[25]
port 201 nsew signal input
rlabel metal3 s 0 18816 400 18872 6 spi_data[26]
port 202 nsew signal input
rlabel metal3 s 0 19488 400 19544 6 spi_data[27]
port 203 nsew signal input
rlabel metal3 s 0 20160 400 20216 6 spi_data[28]
port 204 nsew signal input
rlabel metal3 s 0 20832 400 20888 6 spi_data[29]
port 205 nsew signal input
rlabel metal3 s 0 2688 400 2744 6 spi_data[2]
port 206 nsew signal input
rlabel metal3 s 0 21504 400 21560 6 spi_data[30]
port 207 nsew signal input
rlabel metal3 s 0 22176 400 22232 6 spi_data[31]
port 208 nsew signal input
rlabel metal3 s 0 3360 400 3416 6 spi_data[3]
port 209 nsew signal input
rlabel metal3 s 0 4032 400 4088 6 spi_data[4]
port 210 nsew signal input
rlabel metal3 s 0 4704 400 4760 6 spi_data[5]
port 211 nsew signal input
rlabel metal3 s 0 5376 400 5432 6 spi_data[6]
port 212 nsew signal input
rlabel metal3 s 0 6048 400 6104 6 spi_data[7]
port 213 nsew signal input
rlabel metal3 s 0 6720 400 6776 6 spi_data[8]
port 214 nsew signal input
rlabel metal3 s 0 7392 400 7448 6 spi_data[9]
port 215 nsew signal input
rlabel metal3 s 0 672 400 728 6 spi_data_clock
port 216 nsew signal input
rlabel metal4 s 2224 1538 2384 21198 6 vdd
port 217 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 21198 6 vdd
port 217 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 21198 6 vdd
port 217 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 21198 6 vdd
port 217 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 21198 6 vdd
port 217 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 21198 6 vdd
port 217 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 21198 6 vss
port 218 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 21198 6 vss
port 218 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 21198 6 vss
port 218 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 21198 6 vss
port 218 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 21198 6 vss
port 218 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 80000 23000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4693172
string GDS_FILE /home/jasteve4/Documents/MicroMotorController/openlane/controller_core/runs/22_12_05_21_28/results/signoff/controller_core.magic.gds
string GDS_START 291382
<< end >>


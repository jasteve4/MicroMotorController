VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO spi_core
  CLASS BLOCK ;
  FOREIGN spi_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 250.000 BY 250.000 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 14.560 0.000 15.120 4.000 ;
    END
  END clock
  PIN clock_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 7.840 250.000 8.400 ;
    END
  END clock_out
  PIN data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 15.120 250.000 15.680 ;
    END
  END data_out[0]
  PIN data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 87.920 250.000 88.480 ;
    END
  END data_out[10]
  PIN data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 95.200 250.000 95.760 ;
    END
  END data_out[11]
  PIN data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 102.480 250.000 103.040 ;
    END
  END data_out[12]
  PIN data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 109.760 250.000 110.320 ;
    END
  END data_out[13]
  PIN data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 117.040 250.000 117.600 ;
    END
  END data_out[14]
  PIN data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 124.320 250.000 124.880 ;
    END
  END data_out[15]
  PIN data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 131.600 250.000 132.160 ;
    END
  END data_out[16]
  PIN data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 138.880 250.000 139.440 ;
    END
  END data_out[17]
  PIN data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 146.160 250.000 146.720 ;
    END
  END data_out[18]
  PIN data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 153.440 250.000 154.000 ;
    END
  END data_out[19]
  PIN data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 22.400 250.000 22.960 ;
    END
  END data_out[1]
  PIN data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 160.720 250.000 161.280 ;
    END
  END data_out[20]
  PIN data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 168.000 250.000 168.560 ;
    END
  END data_out[21]
  PIN data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 175.280 250.000 175.840 ;
    END
  END data_out[22]
  PIN data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 182.560 250.000 183.120 ;
    END
  END data_out[23]
  PIN data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 189.840 250.000 190.400 ;
    END
  END data_out[24]
  PIN data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 197.120 250.000 197.680 ;
    END
  END data_out[25]
  PIN data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 204.400 250.000 204.960 ;
    END
  END data_out[26]
  PIN data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 211.680 250.000 212.240 ;
    END
  END data_out[27]
  PIN data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 218.960 250.000 219.520 ;
    END
  END data_out[28]
  PIN data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 226.240 250.000 226.800 ;
    END
  END data_out[29]
  PIN data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 29.680 250.000 30.240 ;
    END
  END data_out[2]
  PIN data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 233.520 250.000 234.080 ;
    END
  END data_out[30]
  PIN data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 240.800 250.000 241.360 ;
    END
  END data_out[31]
  PIN data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 36.960 250.000 37.520 ;
    END
  END data_out[3]
  PIN data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 44.240 250.000 44.800 ;
    END
  END data_out[4]
  PIN data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 51.520 250.000 52.080 ;
    END
  END data_out[5]
  PIN data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 58.800 250.000 59.360 ;
    END
  END data_out[6]
  PIN data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 66.080 250.000 66.640 ;
    END
  END data_out[7]
  PIN data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 73.360 250.000 73.920 ;
    END
  END data_out[8]
  PIN data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 80.640 250.000 81.200 ;
    END
  END data_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 151.760 0.000 152.320 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 179.200 0.000 179.760 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 206.640 0.000 207.200 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 234.080 0.000 234.640 4.000 ;
    END
  END la_data_in[3]
  PIN la_oenb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 42.000 0.000 42.560 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 69.440 0.000 70.000 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 96.880 0.000 97.440 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 0.000 124.880 4.000 ;
    END
  END la_oenb[3]
  PIN miso
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 201.600 4.000 202.160 ;
    END
  END miso
  PIN miso_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 232.400 4.000 232.960 ;
    END
  END miso_oeb
  PIN mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 78.400 4.000 78.960 ;
    END
  END mosi
  PIN mosi_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 109.200 4.000 109.760 ;
    END
  END mosi_oeb
  PIN sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 16.800 4.000 17.360 ;
    END
  END sclk
  PIN sclk_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 47.600 4.000 48.160 ;
    END
  END sclk_oeb
  PIN ss_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 140.000 4.000 140.560 ;
    END
  END ss_n
  PIN ss_n_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 170.800 4.000 171.360 ;
    END
  END ss_n_oeb
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 231.580 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 231.580 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 231.580 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 243.040 231.580 ;
      LAYER Metal2 ;
        RECT 9.100 4.300 240.660 241.270 ;
        RECT 9.100 4.000 14.260 4.300 ;
        RECT 15.420 4.000 41.700 4.300 ;
        RECT 42.860 4.000 69.140 4.300 ;
        RECT 70.300 4.000 96.580 4.300 ;
        RECT 97.740 4.000 124.020 4.300 ;
        RECT 125.180 4.000 151.460 4.300 ;
        RECT 152.620 4.000 178.900 4.300 ;
        RECT 180.060 4.000 206.340 4.300 ;
        RECT 207.500 4.000 233.780 4.300 ;
        RECT 234.940 4.000 240.660 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 240.500 245.700 241.220 ;
        RECT 4.000 234.380 246.820 240.500 ;
        RECT 4.000 233.260 245.700 234.380 ;
        RECT 4.300 233.220 245.700 233.260 ;
        RECT 4.300 232.100 246.820 233.220 ;
        RECT 4.000 227.100 246.820 232.100 ;
        RECT 4.000 225.940 245.700 227.100 ;
        RECT 4.000 219.820 246.820 225.940 ;
        RECT 4.000 218.660 245.700 219.820 ;
        RECT 4.000 212.540 246.820 218.660 ;
        RECT 4.000 211.380 245.700 212.540 ;
        RECT 4.000 205.260 246.820 211.380 ;
        RECT 4.000 204.100 245.700 205.260 ;
        RECT 4.000 202.460 246.820 204.100 ;
        RECT 4.300 201.300 246.820 202.460 ;
        RECT 4.000 197.980 246.820 201.300 ;
        RECT 4.000 196.820 245.700 197.980 ;
        RECT 4.000 190.700 246.820 196.820 ;
        RECT 4.000 189.540 245.700 190.700 ;
        RECT 4.000 183.420 246.820 189.540 ;
        RECT 4.000 182.260 245.700 183.420 ;
        RECT 4.000 176.140 246.820 182.260 ;
        RECT 4.000 174.980 245.700 176.140 ;
        RECT 4.000 171.660 246.820 174.980 ;
        RECT 4.300 170.500 246.820 171.660 ;
        RECT 4.000 168.860 246.820 170.500 ;
        RECT 4.000 167.700 245.700 168.860 ;
        RECT 4.000 161.580 246.820 167.700 ;
        RECT 4.000 160.420 245.700 161.580 ;
        RECT 4.000 154.300 246.820 160.420 ;
        RECT 4.000 153.140 245.700 154.300 ;
        RECT 4.000 147.020 246.820 153.140 ;
        RECT 4.000 145.860 245.700 147.020 ;
        RECT 4.000 140.860 246.820 145.860 ;
        RECT 4.300 139.740 246.820 140.860 ;
        RECT 4.300 139.700 245.700 139.740 ;
        RECT 4.000 138.580 245.700 139.700 ;
        RECT 4.000 132.460 246.820 138.580 ;
        RECT 4.000 131.300 245.700 132.460 ;
        RECT 4.000 125.180 246.820 131.300 ;
        RECT 4.000 124.020 245.700 125.180 ;
        RECT 4.000 117.900 246.820 124.020 ;
        RECT 4.000 116.740 245.700 117.900 ;
        RECT 4.000 110.620 246.820 116.740 ;
        RECT 4.000 110.060 245.700 110.620 ;
        RECT 4.300 109.460 245.700 110.060 ;
        RECT 4.300 108.900 246.820 109.460 ;
        RECT 4.000 103.340 246.820 108.900 ;
        RECT 4.000 102.180 245.700 103.340 ;
        RECT 4.000 96.060 246.820 102.180 ;
        RECT 4.000 94.900 245.700 96.060 ;
        RECT 4.000 88.780 246.820 94.900 ;
        RECT 4.000 87.620 245.700 88.780 ;
        RECT 4.000 81.500 246.820 87.620 ;
        RECT 4.000 80.340 245.700 81.500 ;
        RECT 4.000 79.260 246.820 80.340 ;
        RECT 4.300 78.100 246.820 79.260 ;
        RECT 4.000 74.220 246.820 78.100 ;
        RECT 4.000 73.060 245.700 74.220 ;
        RECT 4.000 66.940 246.820 73.060 ;
        RECT 4.000 65.780 245.700 66.940 ;
        RECT 4.000 59.660 246.820 65.780 ;
        RECT 4.000 58.500 245.700 59.660 ;
        RECT 4.000 52.380 246.820 58.500 ;
        RECT 4.000 51.220 245.700 52.380 ;
        RECT 4.000 48.460 246.820 51.220 ;
        RECT 4.300 47.300 246.820 48.460 ;
        RECT 4.000 45.100 246.820 47.300 ;
        RECT 4.000 43.940 245.700 45.100 ;
        RECT 4.000 37.820 246.820 43.940 ;
        RECT 4.000 36.660 245.700 37.820 ;
        RECT 4.000 30.540 246.820 36.660 ;
        RECT 4.000 29.380 245.700 30.540 ;
        RECT 4.000 23.260 246.820 29.380 ;
        RECT 4.000 22.100 245.700 23.260 ;
        RECT 4.000 17.660 246.820 22.100 ;
        RECT 4.300 16.500 246.820 17.660 ;
        RECT 4.000 15.980 246.820 16.500 ;
        RECT 4.000 14.820 245.700 15.980 ;
        RECT 4.000 8.700 246.820 14.820 ;
        RECT 4.000 7.980 245.700 8.700 ;
  END
END spi_core
END LIBRARY


magic
tech gf180mcuC
magscale 1 5
timestamp 1670294109
<< obsm1 >>
rect 672 1538 24304 23158
<< metal2 >>
rect 6216 0 6272 400
rect 18704 0 18760 400
<< obsm2 >>
rect 854 430 22442 23147
rect 854 350 6186 430
rect 6302 350 18674 430
rect 18790 350 22442 430
<< metal3 >>
rect 0 20720 400 20776
rect 0 12432 400 12488
rect 24600 12432 25000 12488
rect 0 4144 400 4200
<< obsm3 >>
rect 400 20806 24600 23142
rect 430 20690 24600 20806
rect 400 12518 24600 20690
rect 430 12402 24570 12518
rect 400 4230 24600 12402
rect 430 4114 24600 4230
rect 400 1554 24600 4114
<< metal4 >>
rect 2224 1538 2384 23158
rect 9904 1538 10064 23158
rect 17584 1538 17744 23158
<< labels >>
rlabel metal3 s 0 4144 400 4200 6 clock_out_a
port 1 nsew signal output
rlabel metal3 s 0 12432 400 12488 6 clock_out_b
port 2 nsew signal output
rlabel metal3 s 0 20720 400 20776 6 clock_out_c
port 3 nsew signal output
rlabel metal2 s 6216 0 6272 400 6 core_clock
port 4 nsew signal input
rlabel metal3 s 24600 12432 25000 12488 6 io_clock
port 5 nsew signal input
rlabel metal2 s 18704 0 18760 400 6 la_oenb
port 6 nsew signal input
rlabel metal4 s 2224 1538 2384 23158 6 vdd
port 7 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 23158 6 vdd
port 7 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 23158 6 vss
port 8 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 25000 25000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 300606
string GDS_FILE /home/jasteve4/Documents/MicroMotorController/openlane/clock_mux/runs/22_12_05_21_34/results/signoff/clock_mux.magic.gds
string GDS_START 83520
<< end >>


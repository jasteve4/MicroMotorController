VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO controller_core
  CLASS BLOCK ;
  FOREIGN controller_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 800.000 BY 230.000 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 775.600 0.000 776.160 4.000 ;
    END
  END clock
  PIN clock_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 221.200 226.000 221.760 230.000 ;
    END
  END clock_out[0]
  PIN clock_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 227.920 226.000 228.480 230.000 ;
    END
  END clock_out[1]
  PIN clock_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 234.640 226.000 235.200 230.000 ;
    END
  END clock_out[2]
  PIN clock_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 241.360 226.000 241.920 230.000 ;
    END
  END clock_out[3]
  PIN clock_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 248.080 226.000 248.640 230.000 ;
    END
  END clock_out[4]
  PIN clock_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 254.800 226.000 255.360 230.000 ;
    END
  END clock_out[5]
  PIN clock_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 261.520 226.000 262.080 230.000 ;
    END
  END clock_out[6]
  PIN clock_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 268.240 226.000 268.800 230.000 ;
    END
  END clock_out[7]
  PIN clock_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 274.960 226.000 275.520 230.000 ;
    END
  END clock_out[8]
  PIN clock_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 281.680 226.000 282.240 230.000 ;
    END
  END clock_out[9]
  PIN col_select_left[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 409.360 226.000 409.920 230.000 ;
    END
  END col_select_left[0]
  PIN col_select_left[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 416.080 226.000 416.640 230.000 ;
    END
  END col_select_left[1]
  PIN col_select_left[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 422.800 226.000 423.360 230.000 ;
    END
  END col_select_left[2]
  PIN col_select_left[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 429.520 226.000 430.080 230.000 ;
    END
  END col_select_left[3]
  PIN col_select_left[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 436.240 226.000 436.800 230.000 ;
    END
  END col_select_left[4]
  PIN col_select_left[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 442.960 226.000 443.520 230.000 ;
    END
  END col_select_left[5]
  PIN col_select_right[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 369.040 226.000 369.600 230.000 ;
    END
  END col_select_right[0]
  PIN col_select_right[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 375.760 226.000 376.320 230.000 ;
    END
  END col_select_right[1]
  PIN col_select_right[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 382.480 226.000 383.040 230.000 ;
    END
  END col_select_right[2]
  PIN col_select_right[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 389.200 226.000 389.760 230.000 ;
    END
  END col_select_right[3]
  PIN col_select_right[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 395.920 226.000 396.480 230.000 ;
    END
  END col_select_right[4]
  PIN col_select_right[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 402.640 226.000 403.200 230.000 ;
    END
  END col_select_right[5]
  PIN data_out_left[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 557.200 226.000 557.760 230.000 ;
    END
  END data_out_left[0]
  PIN data_out_left[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 624.400 226.000 624.960 230.000 ;
    END
  END data_out_left[10]
  PIN data_out_left[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 631.120 226.000 631.680 230.000 ;
    END
  END data_out_left[11]
  PIN data_out_left[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 637.840 226.000 638.400 230.000 ;
    END
  END data_out_left[12]
  PIN data_out_left[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 644.560 226.000 645.120 230.000 ;
    END
  END data_out_left[13]
  PIN data_out_left[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 651.280 226.000 651.840 230.000 ;
    END
  END data_out_left[14]
  PIN data_out_left[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 658.000 226.000 658.560 230.000 ;
    END
  END data_out_left[15]
  PIN data_out_left[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 563.920 226.000 564.480 230.000 ;
    END
  END data_out_left[1]
  PIN data_out_left[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 570.640 226.000 571.200 230.000 ;
    END
  END data_out_left[2]
  PIN data_out_left[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 577.360 226.000 577.920 230.000 ;
    END
  END data_out_left[3]
  PIN data_out_left[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 584.080 226.000 584.640 230.000 ;
    END
  END data_out_left[4]
  PIN data_out_left[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 590.800 226.000 591.360 230.000 ;
    END
  END data_out_left[5]
  PIN data_out_left[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 597.520 226.000 598.080 230.000 ;
    END
  END data_out_left[6]
  PIN data_out_left[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 604.240 226.000 604.800 230.000 ;
    END
  END data_out_left[7]
  PIN data_out_left[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 610.960 226.000 611.520 230.000 ;
    END
  END data_out_left[8]
  PIN data_out_left[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 617.680 226.000 618.240 230.000 ;
    END
  END data_out_left[9]
  PIN data_out_right[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 449.680 226.000 450.240 230.000 ;
    END
  END data_out_right[0]
  PIN data_out_right[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 516.880 226.000 517.440 230.000 ;
    END
  END data_out_right[10]
  PIN data_out_right[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 523.600 226.000 524.160 230.000 ;
    END
  END data_out_right[11]
  PIN data_out_right[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 530.320 226.000 530.880 230.000 ;
    END
  END data_out_right[12]
  PIN data_out_right[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 537.040 226.000 537.600 230.000 ;
    END
  END data_out_right[13]
  PIN data_out_right[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 543.760 226.000 544.320 230.000 ;
    END
  END data_out_right[14]
  PIN data_out_right[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 550.480 226.000 551.040 230.000 ;
    END
  END data_out_right[15]
  PIN data_out_right[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 456.400 226.000 456.960 230.000 ;
    END
  END data_out_right[1]
  PIN data_out_right[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 463.120 226.000 463.680 230.000 ;
    END
  END data_out_right[2]
  PIN data_out_right[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 469.840 226.000 470.400 230.000 ;
    END
  END data_out_right[3]
  PIN data_out_right[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 476.560 226.000 477.120 230.000 ;
    END
  END data_out_right[4]
  PIN data_out_right[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 483.280 226.000 483.840 230.000 ;
    END
  END data_out_right[5]
  PIN data_out_right[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 490.000 226.000 490.560 230.000 ;
    END
  END data_out_right[6]
  PIN data_out_right[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 496.720 226.000 497.280 230.000 ;
    END
  END data_out_right[7]
  PIN data_out_right[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 503.440 226.000 504.000 230.000 ;
    END
  END data_out_right[8]
  PIN data_out_right[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 510.160 226.000 510.720 230.000 ;
    END
  END data_out_right[9]
  PIN inverter_select[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 731.920 226.000 732.480 230.000 ;
    END
  END inverter_select[0]
  PIN inverter_select[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 738.640 226.000 739.200 230.000 ;
    END
  END inverter_select[1]
  PIN inverter_select[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 745.360 226.000 745.920 230.000 ;
    END
  END inverter_select[2]
  PIN inverter_select[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 752.080 226.000 752.640 230.000 ;
    END
  END inverter_select[3]
  PIN inverter_select[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 758.800 226.000 759.360 230.000 ;
    END
  END inverter_select[4]
  PIN inverter_select[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 765.520 226.000 766.080 230.000 ;
    END
  END inverter_select[5]
  PIN inverter_select[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 772.240 226.000 772.800 230.000 ;
    END
  END inverter_select[6]
  PIN inverter_select[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 778.960 226.000 779.520 230.000 ;
    END
  END inverter_select[7]
  PIN inverter_select[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 785.680 226.000 786.240 230.000 ;
    END
  END inverter_select[8]
  PIN inverter_select[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 792.400 226.000 792.960 230.000 ;
    END
  END inverter_select[9]
  PIN io_control_trigger_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 70.000 0.000 70.560 4.000 ;
    END
  END io_control_trigger_in
  PIN io_control_trigger_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 81.760 0.000 82.320 4.000 ;
    END
  END io_control_trigger_oeb
  PIN io_driver_io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 117.040 0.000 117.600 4.000 ;
    END
  END io_driver_io_oeb[0]
  PIN io_driver_io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 234.640 0.000 235.200 4.000 ;
    END
  END io_driver_io_oeb[10]
  PIN io_driver_io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 246.400 0.000 246.960 4.000 ;
    END
  END io_driver_io_oeb[11]
  PIN io_driver_io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 258.160 0.000 258.720 4.000 ;
    END
  END io_driver_io_oeb[12]
  PIN io_driver_io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 269.920 0.000 270.480 4.000 ;
    END
  END io_driver_io_oeb[13]
  PIN io_driver_io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 281.680 0.000 282.240 4.000 ;
    END
  END io_driver_io_oeb[14]
  PIN io_driver_io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 293.440 0.000 294.000 4.000 ;
    END
  END io_driver_io_oeb[15]
  PIN io_driver_io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 305.200 0.000 305.760 4.000 ;
    END
  END io_driver_io_oeb[16]
  PIN io_driver_io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 316.960 0.000 317.520 4.000 ;
    END
  END io_driver_io_oeb[17]
  PIN io_driver_io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 328.720 0.000 329.280 4.000 ;
    END
  END io_driver_io_oeb[18]
  PIN io_driver_io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 340.480 0.000 341.040 4.000 ;
    END
  END io_driver_io_oeb[19]
  PIN io_driver_io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 128.800 0.000 129.360 4.000 ;
    END
  END io_driver_io_oeb[1]
  PIN io_driver_io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 140.560 0.000 141.120 4.000 ;
    END
  END io_driver_io_oeb[2]
  PIN io_driver_io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 152.320 0.000 152.880 4.000 ;
    END
  END io_driver_io_oeb[3]
  PIN io_driver_io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 164.080 0.000 164.640 4.000 ;
    END
  END io_driver_io_oeb[4]
  PIN io_driver_io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 175.840 0.000 176.400 4.000 ;
    END
  END io_driver_io_oeb[5]
  PIN io_driver_io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 187.600 0.000 188.160 4.000 ;
    END
  END io_driver_io_oeb[6]
  PIN io_driver_io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 199.360 0.000 199.920 4.000 ;
    END
  END io_driver_io_oeb[7]
  PIN io_driver_io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 211.120 0.000 211.680 4.000 ;
    END
  END io_driver_io_oeb[8]
  PIN io_driver_io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 222.880 0.000 223.440 4.000 ;
    END
  END io_driver_io_oeb[9]
  PIN io_latch_data_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 46.480 0.000 47.040 4.000 ;
    END
  END io_latch_data_in
  PIN io_latch_data_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 58.240 0.000 58.800 4.000 ;
    END
  END io_latch_data_oeb
  PIN io_reset_n_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 22.960 0.000 23.520 4.000 ;
    END
  END io_reset_n_in
  PIN io_reset_n_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 34.720 0.000 35.280 4.000 ;
    END
  END io_reset_n_oeb
  PIN io_update_cycle_complete_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 105.280 0.000 105.840 4.000 ;
    END
  END io_update_cycle_complete_oeb
  PIN io_update_cycle_complete_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 93.520 0.000 94.080 4.000 ;
    END
  END io_update_cycle_complete_out
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 563.920 0.000 564.480 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 681.520 0.000 682.080 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 693.280 0.000 693.840 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 705.040 0.000 705.600 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 716.800 0.000 717.360 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 728.560 0.000 729.120 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 740.320 0.000 740.880 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 752.080 0.000 752.640 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 763.840 0.000 764.400 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 575.680 0.000 576.240 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 587.440 0.000 588.000 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 599.200 0.000 599.760 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 610.960 0.000 611.520 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 622.720 0.000 623.280 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 634.480 0.000 635.040 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 646.240 0.000 646.800 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 658.000 0.000 658.560 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 669.760 0.000 670.320 4.000 ;
    END
  END la_data_in[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 352.240 0.000 352.800 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 469.840 0.000 470.400 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 481.600 0.000 482.160 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 493.360 0.000 493.920 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 505.120 0.000 505.680 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 516.880 0.000 517.440 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 528.640 0.000 529.200 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 540.400 0.000 540.960 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 552.160 0.000 552.720 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 364.000 0.000 364.560 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 375.760 0.000 376.320 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 387.520 0.000 388.080 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 399.280 0.000 399.840 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 411.040 0.000 411.600 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 422.800 0.000 423.360 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 434.560 0.000 435.120 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 446.320 0.000 446.880 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 458.080 0.000 458.640 4.000 ;
    END
  END la_oenb[9]
  PIN mem_address_left[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 86.800 226.000 87.360 230.000 ;
    END
  END mem_address_left[0]
  PIN mem_address_left[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 93.520 226.000 94.080 230.000 ;
    END
  END mem_address_left[1]
  PIN mem_address_left[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 100.240 226.000 100.800 230.000 ;
    END
  END mem_address_left[2]
  PIN mem_address_left[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 106.960 226.000 107.520 230.000 ;
    END
  END mem_address_left[3]
  PIN mem_address_left[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 113.680 226.000 114.240 230.000 ;
    END
  END mem_address_left[4]
  PIN mem_address_left[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 120.400 226.000 120.960 230.000 ;
    END
  END mem_address_left[5]
  PIN mem_address_left[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 127.120 226.000 127.680 230.000 ;
    END
  END mem_address_left[6]
  PIN mem_address_left[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 133.840 226.000 134.400 230.000 ;
    END
  END mem_address_left[7]
  PIN mem_address_left[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 140.560 226.000 141.120 230.000 ;
    END
  END mem_address_left[8]
  PIN mem_address_left[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 147.280 226.000 147.840 230.000 ;
    END
  END mem_address_left[9]
  PIN mem_address_right[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 19.600 226.000 20.160 230.000 ;
    END
  END mem_address_right[0]
  PIN mem_address_right[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.320 226.000 26.880 230.000 ;
    END
  END mem_address_right[1]
  PIN mem_address_right[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 33.040 226.000 33.600 230.000 ;
    END
  END mem_address_right[2]
  PIN mem_address_right[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 39.760 226.000 40.320 230.000 ;
    END
  END mem_address_right[3]
  PIN mem_address_right[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 46.480 226.000 47.040 230.000 ;
    END
  END mem_address_right[4]
  PIN mem_address_right[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 53.200 226.000 53.760 230.000 ;
    END
  END mem_address_right[5]
  PIN mem_address_right[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 59.920 226.000 60.480 230.000 ;
    END
  END mem_address_right[6]
  PIN mem_address_right[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 66.640 226.000 67.200 230.000 ;
    END
  END mem_address_right[7]
  PIN mem_address_right[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 73.360 226.000 73.920 230.000 ;
    END
  END mem_address_right[8]
  PIN mem_address_right[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 80.080 226.000 80.640 230.000 ;
    END
  END mem_address_right[9]
  PIN mem_write_n[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 154.000 226.000 154.560 230.000 ;
    END
  END mem_write_n[0]
  PIN mem_write_n[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 160.720 226.000 161.280 230.000 ;
    END
  END mem_write_n[1]
  PIN mem_write_n[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 167.440 226.000 168.000 230.000 ;
    END
  END mem_write_n[2]
  PIN mem_write_n[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 174.160 226.000 174.720 230.000 ;
    END
  END mem_write_n[3]
  PIN mem_write_n[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 180.880 226.000 181.440 230.000 ;
    END
  END mem_write_n[4]
  PIN mem_write_n[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 187.600 226.000 188.160 230.000 ;
    END
  END mem_write_n[5]
  PIN mem_write_n[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 194.320 226.000 194.880 230.000 ;
    END
  END mem_write_n[6]
  PIN mem_write_n[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 201.040 226.000 201.600 230.000 ;
    END
  END mem_write_n[7]
  PIN mem_write_n[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 207.760 226.000 208.320 230.000 ;
    END
  END mem_write_n[8]
  PIN mem_write_n[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 214.480 226.000 215.040 230.000 ;
    END
  END mem_write_n[9]
  PIN output_active_left
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 12.880 226.000 13.440 230.000 ;
    END
  END output_active_left
  PIN output_active_right
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 6.160 226.000 6.720 230.000 ;
    END
  END output_active_right
  PIN row_col_select[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 664.720 226.000 665.280 230.000 ;
    END
  END row_col_select[0]
  PIN row_col_select[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 671.440 226.000 672.000 230.000 ;
    END
  END row_col_select[1]
  PIN row_col_select[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 678.160 226.000 678.720 230.000 ;
    END
  END row_col_select[2]
  PIN row_col_select[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 684.880 226.000 685.440 230.000 ;
    END
  END row_col_select[3]
  PIN row_col_select[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 691.600 226.000 692.160 230.000 ;
    END
  END row_col_select[4]
  PIN row_col_select[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 698.320 226.000 698.880 230.000 ;
    END
  END row_col_select[5]
  PIN row_col_select[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 705.040 226.000 705.600 230.000 ;
    END
  END row_col_select[6]
  PIN row_col_select[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 711.760 226.000 712.320 230.000 ;
    END
  END row_col_select[7]
  PIN row_col_select[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 718.480 226.000 719.040 230.000 ;
    END
  END row_col_select[8]
  PIN row_col_select[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 725.200 226.000 725.760 230.000 ;
    END
  END row_col_select[9]
  PIN row_select_left[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 328.720 226.000 329.280 230.000 ;
    END
  END row_select_left[0]
  PIN row_select_left[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 335.440 226.000 336.000 230.000 ;
    END
  END row_select_left[1]
  PIN row_select_left[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 342.160 226.000 342.720 230.000 ;
    END
  END row_select_left[2]
  PIN row_select_left[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 348.880 226.000 349.440 230.000 ;
    END
  END row_select_left[3]
  PIN row_select_left[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 355.600 226.000 356.160 230.000 ;
    END
  END row_select_left[4]
  PIN row_select_left[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 362.320 226.000 362.880 230.000 ;
    END
  END row_select_left[5]
  PIN row_select_right[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 288.400 226.000 288.960 230.000 ;
    END
  END row_select_right[0]
  PIN row_select_right[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 295.120 226.000 295.680 230.000 ;
    END
  END row_select_right[1]
  PIN row_select_right[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 301.840 226.000 302.400 230.000 ;
    END
  END row_select_right[2]
  PIN row_select_right[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 308.560 226.000 309.120 230.000 ;
    END
  END row_select_right[3]
  PIN row_select_right[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 315.280 226.000 315.840 230.000 ;
    END
  END row_select_right[4]
  PIN row_select_right[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 322.000 226.000 322.560 230.000 ;
    END
  END row_select_right[5]
  PIN spi_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 13.440 4.000 14.000 ;
    END
  END spi_data[0]
  PIN spi_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 80.640 4.000 81.200 ;
    END
  END spi_data[10]
  PIN spi_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 87.360 4.000 87.920 ;
    END
  END spi_data[11]
  PIN spi_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 94.080 4.000 94.640 ;
    END
  END spi_data[12]
  PIN spi_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 100.800 4.000 101.360 ;
    END
  END spi_data[13]
  PIN spi_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 107.520 4.000 108.080 ;
    END
  END spi_data[14]
  PIN spi_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 114.240 4.000 114.800 ;
    END
  END spi_data[15]
  PIN spi_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 120.960 4.000 121.520 ;
    END
  END spi_data[16]
  PIN spi_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 127.680 4.000 128.240 ;
    END
  END spi_data[17]
  PIN spi_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 134.400 4.000 134.960 ;
    END
  END spi_data[18]
  PIN spi_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 141.120 4.000 141.680 ;
    END
  END spi_data[19]
  PIN spi_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 20.160 4.000 20.720 ;
    END
  END spi_data[1]
  PIN spi_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 147.840 4.000 148.400 ;
    END
  END spi_data[20]
  PIN spi_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 154.560 4.000 155.120 ;
    END
  END spi_data[21]
  PIN spi_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 161.280 4.000 161.840 ;
    END
  END spi_data[22]
  PIN spi_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 168.000 4.000 168.560 ;
    END
  END spi_data[23]
  PIN spi_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 174.720 4.000 175.280 ;
    END
  END spi_data[24]
  PIN spi_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 181.440 4.000 182.000 ;
    END
  END spi_data[25]
  PIN spi_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 188.160 4.000 188.720 ;
    END
  END spi_data[26]
  PIN spi_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 194.880 4.000 195.440 ;
    END
  END spi_data[27]
  PIN spi_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 201.600 4.000 202.160 ;
    END
  END spi_data[28]
  PIN spi_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 208.320 4.000 208.880 ;
    END
  END spi_data[29]
  PIN spi_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 26.880 4.000 27.440 ;
    END
  END spi_data[2]
  PIN spi_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 215.040 4.000 215.600 ;
    END
  END spi_data[30]
  PIN spi_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 221.760 4.000 222.320 ;
    END
  END spi_data[31]
  PIN spi_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 33.600 4.000 34.160 ;
    END
  END spi_data[3]
  PIN spi_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 40.320 4.000 40.880 ;
    END
  END spi_data[4]
  PIN spi_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 47.040 4.000 47.600 ;
    END
  END spi_data[5]
  PIN spi_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 53.760 4.000 54.320 ;
    END
  END spi_data[6]
  PIN spi_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 60.480 4.000 61.040 ;
    END
  END spi_data[7]
  PIN spi_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 67.200 4.000 67.760 ;
    END
  END spi_data[8]
  PIN spi_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 73.920 4.000 74.480 ;
    END
  END spi_data[9]
  PIN spi_data_clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 6.720 4.000 7.280 ;
    END
  END spi_data_clock
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 211.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 211.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 211.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 211.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 211.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 211.980 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 211.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 211.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 211.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 211.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 211.980 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 792.960 214.890 ;
      LAYER Metal2 ;
        RECT 7.020 225.700 12.580 226.660 ;
        RECT 13.740 225.700 19.300 226.660 ;
        RECT 20.460 225.700 26.020 226.660 ;
        RECT 27.180 225.700 32.740 226.660 ;
        RECT 33.900 225.700 39.460 226.660 ;
        RECT 40.620 225.700 46.180 226.660 ;
        RECT 47.340 225.700 52.900 226.660 ;
        RECT 54.060 225.700 59.620 226.660 ;
        RECT 60.780 225.700 66.340 226.660 ;
        RECT 67.500 225.700 73.060 226.660 ;
        RECT 74.220 225.700 79.780 226.660 ;
        RECT 80.940 225.700 86.500 226.660 ;
        RECT 87.660 225.700 93.220 226.660 ;
        RECT 94.380 225.700 99.940 226.660 ;
        RECT 101.100 225.700 106.660 226.660 ;
        RECT 107.820 225.700 113.380 226.660 ;
        RECT 114.540 225.700 120.100 226.660 ;
        RECT 121.260 225.700 126.820 226.660 ;
        RECT 127.980 225.700 133.540 226.660 ;
        RECT 134.700 225.700 140.260 226.660 ;
        RECT 141.420 225.700 146.980 226.660 ;
        RECT 148.140 225.700 153.700 226.660 ;
        RECT 154.860 225.700 160.420 226.660 ;
        RECT 161.580 225.700 167.140 226.660 ;
        RECT 168.300 225.700 173.860 226.660 ;
        RECT 175.020 225.700 180.580 226.660 ;
        RECT 181.740 225.700 187.300 226.660 ;
        RECT 188.460 225.700 194.020 226.660 ;
        RECT 195.180 225.700 200.740 226.660 ;
        RECT 201.900 225.700 207.460 226.660 ;
        RECT 208.620 225.700 214.180 226.660 ;
        RECT 215.340 225.700 220.900 226.660 ;
        RECT 222.060 225.700 227.620 226.660 ;
        RECT 228.780 225.700 234.340 226.660 ;
        RECT 235.500 225.700 241.060 226.660 ;
        RECT 242.220 225.700 247.780 226.660 ;
        RECT 248.940 225.700 254.500 226.660 ;
        RECT 255.660 225.700 261.220 226.660 ;
        RECT 262.380 225.700 267.940 226.660 ;
        RECT 269.100 225.700 274.660 226.660 ;
        RECT 275.820 225.700 281.380 226.660 ;
        RECT 282.540 225.700 288.100 226.660 ;
        RECT 289.260 225.700 294.820 226.660 ;
        RECT 295.980 225.700 301.540 226.660 ;
        RECT 302.700 225.700 308.260 226.660 ;
        RECT 309.420 225.700 314.980 226.660 ;
        RECT 316.140 225.700 321.700 226.660 ;
        RECT 322.860 225.700 328.420 226.660 ;
        RECT 329.580 225.700 335.140 226.660 ;
        RECT 336.300 225.700 341.860 226.660 ;
        RECT 343.020 225.700 348.580 226.660 ;
        RECT 349.740 225.700 355.300 226.660 ;
        RECT 356.460 225.700 362.020 226.660 ;
        RECT 363.180 225.700 368.740 226.660 ;
        RECT 369.900 225.700 375.460 226.660 ;
        RECT 376.620 225.700 382.180 226.660 ;
        RECT 383.340 225.700 388.900 226.660 ;
        RECT 390.060 225.700 395.620 226.660 ;
        RECT 396.780 225.700 402.340 226.660 ;
        RECT 403.500 225.700 409.060 226.660 ;
        RECT 410.220 225.700 415.780 226.660 ;
        RECT 416.940 225.700 422.500 226.660 ;
        RECT 423.660 225.700 429.220 226.660 ;
        RECT 430.380 225.700 435.940 226.660 ;
        RECT 437.100 225.700 442.660 226.660 ;
        RECT 443.820 225.700 449.380 226.660 ;
        RECT 450.540 225.700 456.100 226.660 ;
        RECT 457.260 225.700 462.820 226.660 ;
        RECT 463.980 225.700 469.540 226.660 ;
        RECT 470.700 225.700 476.260 226.660 ;
        RECT 477.420 225.700 482.980 226.660 ;
        RECT 484.140 225.700 489.700 226.660 ;
        RECT 490.860 225.700 496.420 226.660 ;
        RECT 497.580 225.700 503.140 226.660 ;
        RECT 504.300 225.700 509.860 226.660 ;
        RECT 511.020 225.700 516.580 226.660 ;
        RECT 517.740 225.700 523.300 226.660 ;
        RECT 524.460 225.700 530.020 226.660 ;
        RECT 531.180 225.700 536.740 226.660 ;
        RECT 537.900 225.700 543.460 226.660 ;
        RECT 544.620 225.700 550.180 226.660 ;
        RECT 551.340 225.700 556.900 226.660 ;
        RECT 558.060 225.700 563.620 226.660 ;
        RECT 564.780 225.700 570.340 226.660 ;
        RECT 571.500 225.700 577.060 226.660 ;
        RECT 578.220 225.700 583.780 226.660 ;
        RECT 584.940 225.700 590.500 226.660 ;
        RECT 591.660 225.700 597.220 226.660 ;
        RECT 598.380 225.700 603.940 226.660 ;
        RECT 605.100 225.700 610.660 226.660 ;
        RECT 611.820 225.700 617.380 226.660 ;
        RECT 618.540 225.700 624.100 226.660 ;
        RECT 625.260 225.700 630.820 226.660 ;
        RECT 631.980 225.700 637.540 226.660 ;
        RECT 638.700 225.700 644.260 226.660 ;
        RECT 645.420 225.700 650.980 226.660 ;
        RECT 652.140 225.700 657.700 226.660 ;
        RECT 658.860 225.700 664.420 226.660 ;
        RECT 665.580 225.700 671.140 226.660 ;
        RECT 672.300 225.700 677.860 226.660 ;
        RECT 679.020 225.700 684.580 226.660 ;
        RECT 685.740 225.700 691.300 226.660 ;
        RECT 692.460 225.700 698.020 226.660 ;
        RECT 699.180 225.700 704.740 226.660 ;
        RECT 705.900 225.700 711.460 226.660 ;
        RECT 712.620 225.700 718.180 226.660 ;
        RECT 719.340 225.700 724.900 226.660 ;
        RECT 726.060 225.700 731.620 226.660 ;
        RECT 732.780 225.700 738.340 226.660 ;
        RECT 739.500 225.700 745.060 226.660 ;
        RECT 746.220 225.700 751.780 226.660 ;
        RECT 752.940 225.700 758.500 226.660 ;
        RECT 759.660 225.700 765.220 226.660 ;
        RECT 766.380 225.700 771.940 226.660 ;
        RECT 773.100 225.700 778.660 226.660 ;
        RECT 779.820 225.700 785.380 226.660 ;
        RECT 786.540 225.700 792.100 226.660 ;
        RECT 793.260 225.700 793.940 226.660 ;
        RECT 6.300 4.300 793.940 225.700 ;
        RECT 6.300 3.500 22.660 4.300 ;
        RECT 23.820 3.500 34.420 4.300 ;
        RECT 35.580 3.500 46.180 4.300 ;
        RECT 47.340 3.500 57.940 4.300 ;
        RECT 59.100 3.500 69.700 4.300 ;
        RECT 70.860 3.500 81.460 4.300 ;
        RECT 82.620 3.500 93.220 4.300 ;
        RECT 94.380 3.500 104.980 4.300 ;
        RECT 106.140 3.500 116.740 4.300 ;
        RECT 117.900 3.500 128.500 4.300 ;
        RECT 129.660 3.500 140.260 4.300 ;
        RECT 141.420 3.500 152.020 4.300 ;
        RECT 153.180 3.500 163.780 4.300 ;
        RECT 164.940 3.500 175.540 4.300 ;
        RECT 176.700 3.500 187.300 4.300 ;
        RECT 188.460 3.500 199.060 4.300 ;
        RECT 200.220 3.500 210.820 4.300 ;
        RECT 211.980 3.500 222.580 4.300 ;
        RECT 223.740 3.500 234.340 4.300 ;
        RECT 235.500 3.500 246.100 4.300 ;
        RECT 247.260 3.500 257.860 4.300 ;
        RECT 259.020 3.500 269.620 4.300 ;
        RECT 270.780 3.500 281.380 4.300 ;
        RECT 282.540 3.500 293.140 4.300 ;
        RECT 294.300 3.500 304.900 4.300 ;
        RECT 306.060 3.500 316.660 4.300 ;
        RECT 317.820 3.500 328.420 4.300 ;
        RECT 329.580 3.500 340.180 4.300 ;
        RECT 341.340 3.500 351.940 4.300 ;
        RECT 353.100 3.500 363.700 4.300 ;
        RECT 364.860 3.500 375.460 4.300 ;
        RECT 376.620 3.500 387.220 4.300 ;
        RECT 388.380 3.500 398.980 4.300 ;
        RECT 400.140 3.500 410.740 4.300 ;
        RECT 411.900 3.500 422.500 4.300 ;
        RECT 423.660 3.500 434.260 4.300 ;
        RECT 435.420 3.500 446.020 4.300 ;
        RECT 447.180 3.500 457.780 4.300 ;
        RECT 458.940 3.500 469.540 4.300 ;
        RECT 470.700 3.500 481.300 4.300 ;
        RECT 482.460 3.500 493.060 4.300 ;
        RECT 494.220 3.500 504.820 4.300 ;
        RECT 505.980 3.500 516.580 4.300 ;
        RECT 517.740 3.500 528.340 4.300 ;
        RECT 529.500 3.500 540.100 4.300 ;
        RECT 541.260 3.500 551.860 4.300 ;
        RECT 553.020 3.500 563.620 4.300 ;
        RECT 564.780 3.500 575.380 4.300 ;
        RECT 576.540 3.500 587.140 4.300 ;
        RECT 588.300 3.500 598.900 4.300 ;
        RECT 600.060 3.500 610.660 4.300 ;
        RECT 611.820 3.500 622.420 4.300 ;
        RECT 623.580 3.500 634.180 4.300 ;
        RECT 635.340 3.500 645.940 4.300 ;
        RECT 647.100 3.500 657.700 4.300 ;
        RECT 658.860 3.500 669.460 4.300 ;
        RECT 670.620 3.500 681.220 4.300 ;
        RECT 682.380 3.500 692.980 4.300 ;
        RECT 694.140 3.500 704.740 4.300 ;
        RECT 705.900 3.500 716.500 4.300 ;
        RECT 717.660 3.500 728.260 4.300 ;
        RECT 729.420 3.500 740.020 4.300 ;
        RECT 741.180 3.500 751.780 4.300 ;
        RECT 752.940 3.500 763.540 4.300 ;
        RECT 764.700 3.500 775.300 4.300 ;
        RECT 776.460 3.500 793.940 4.300 ;
      LAYER Metal3 ;
        RECT 3.500 222.620 793.990 226.100 ;
        RECT 4.300 221.460 793.990 222.620 ;
        RECT 3.500 215.900 793.990 221.460 ;
        RECT 4.300 214.740 793.990 215.900 ;
        RECT 3.500 209.180 793.990 214.740 ;
        RECT 4.300 208.020 793.990 209.180 ;
        RECT 3.500 202.460 793.990 208.020 ;
        RECT 4.300 201.300 793.990 202.460 ;
        RECT 3.500 195.740 793.990 201.300 ;
        RECT 4.300 194.580 793.990 195.740 ;
        RECT 3.500 189.020 793.990 194.580 ;
        RECT 4.300 187.860 793.990 189.020 ;
        RECT 3.500 182.300 793.990 187.860 ;
        RECT 4.300 181.140 793.990 182.300 ;
        RECT 3.500 175.580 793.990 181.140 ;
        RECT 4.300 174.420 793.990 175.580 ;
        RECT 3.500 168.860 793.990 174.420 ;
        RECT 4.300 167.700 793.990 168.860 ;
        RECT 3.500 162.140 793.990 167.700 ;
        RECT 4.300 160.980 793.990 162.140 ;
        RECT 3.500 155.420 793.990 160.980 ;
        RECT 4.300 154.260 793.990 155.420 ;
        RECT 3.500 148.700 793.990 154.260 ;
        RECT 4.300 147.540 793.990 148.700 ;
        RECT 3.500 141.980 793.990 147.540 ;
        RECT 4.300 140.820 793.990 141.980 ;
        RECT 3.500 135.260 793.990 140.820 ;
        RECT 4.300 134.100 793.990 135.260 ;
        RECT 3.500 128.540 793.990 134.100 ;
        RECT 4.300 127.380 793.990 128.540 ;
        RECT 3.500 121.820 793.990 127.380 ;
        RECT 4.300 120.660 793.990 121.820 ;
        RECT 3.500 115.100 793.990 120.660 ;
        RECT 4.300 113.940 793.990 115.100 ;
        RECT 3.500 108.380 793.990 113.940 ;
        RECT 4.300 107.220 793.990 108.380 ;
        RECT 3.500 101.660 793.990 107.220 ;
        RECT 4.300 100.500 793.990 101.660 ;
        RECT 3.500 94.940 793.990 100.500 ;
        RECT 4.300 93.780 793.990 94.940 ;
        RECT 3.500 88.220 793.990 93.780 ;
        RECT 4.300 87.060 793.990 88.220 ;
        RECT 3.500 81.500 793.990 87.060 ;
        RECT 4.300 80.340 793.990 81.500 ;
        RECT 3.500 74.780 793.990 80.340 ;
        RECT 4.300 73.620 793.990 74.780 ;
        RECT 3.500 68.060 793.990 73.620 ;
        RECT 4.300 66.900 793.990 68.060 ;
        RECT 3.500 61.340 793.990 66.900 ;
        RECT 4.300 60.180 793.990 61.340 ;
        RECT 3.500 54.620 793.990 60.180 ;
        RECT 4.300 53.460 793.990 54.620 ;
        RECT 3.500 47.900 793.990 53.460 ;
        RECT 4.300 46.740 793.990 47.900 ;
        RECT 3.500 41.180 793.990 46.740 ;
        RECT 4.300 40.020 793.990 41.180 ;
        RECT 3.500 34.460 793.990 40.020 ;
        RECT 4.300 33.300 793.990 34.460 ;
        RECT 3.500 27.740 793.990 33.300 ;
        RECT 4.300 26.580 793.990 27.740 ;
        RECT 3.500 21.020 793.990 26.580 ;
        RECT 4.300 19.860 793.990 21.020 ;
        RECT 3.500 14.300 793.990 19.860 ;
        RECT 4.300 13.140 793.990 14.300 ;
        RECT 3.500 7.580 793.990 13.140 ;
        RECT 4.300 6.420 793.990 7.580 ;
        RECT 3.500 4.620 793.990 6.420 ;
      LAYER Metal4 ;
        RECT 153.020 48.250 175.540 195.910 ;
        RECT 177.740 48.250 252.340 195.910 ;
        RECT 254.540 48.250 329.140 195.910 ;
        RECT 331.340 48.250 405.940 195.910 ;
        RECT 408.140 48.250 482.740 195.910 ;
        RECT 484.940 48.250 559.540 195.910 ;
        RECT 561.740 48.250 636.340 195.910 ;
        RECT 638.540 48.250 713.140 195.910 ;
        RECT 715.340 48.250 748.020 195.910 ;
  END
END controller_core
END LIBRARY


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2960.200 BY 2960.200 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 1202.040 2965.000 1203.160 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2255.960 2957.800 2257.080 2965.000 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1928.920 2957.800 1930.040 2965.000 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1601.880 2957.800 1603.000 2965.000 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1274.840 2957.800 1275.960 2965.000 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 947.800 2957.800 948.920 2965.000 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 620.760 2957.800 621.880 2965.000 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 293.720 2957.800 294.840 2965.000 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2919.000 2.400 2920.120 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2701.720 2.400 2702.840 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2484.440 2.400 2485.560 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 1423.800 2965.000 1424.920 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2267.160 2.400 2268.280 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2049.880 2.400 2051.000 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1832.600 2.400 1833.720 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1615.320 2.400 1616.440 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1398.040 2.400 1399.160 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1180.760 2.400 1181.880 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 963.480 2.400 964.600 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 746.200 2.400 747.320 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 528.920 2.400 530.040 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 1645.560 2965.000 1646.680 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 1867.320 2965.000 1868.440 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 2089.080 2965.000 2090.200 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 2310.840 2965.000 2311.960 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 2532.600 2965.000 2533.720 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 2754.360 2965.000 2755.480 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2910.040 2957.800 2911.160 2965.000 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2583.000 2957.800 2584.120 2965.000 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 37.800 2965.000 38.920 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 1922.760 2965.000 1923.880 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 2144.520 2965.000 2145.640 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 2366.280 2965.000 2367.400 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 2588.040 2965.000 2589.160 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 2809.800 2965.000 2810.920 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2828.280 2957.800 2829.400 2965.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2501.240 2957.800 2502.360 2965.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2174.200 2957.800 2175.320 2965.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1847.160 2957.800 1848.280 2965.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1520.120 2957.800 1521.240 2965.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 204.120 2965.000 205.240 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1193.080 2957.800 1194.200 2965.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 866.040 2957.800 867.160 2965.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 539.000 2957.800 540.120 2965.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 211.960 2957.800 213.080 2965.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2864.680 2.400 2865.800 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2647.400 2.400 2648.520 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2430.120 2.400 2431.240 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2212.840 2.400 2213.960 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1995.560 2.400 1996.680 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1778.280 2.400 1779.400 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 370.440 2965.000 371.560 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1561.000 2.400 1562.120 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1343.720 2.400 1344.840 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1126.440 2.400 1127.560 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 909.160 2.400 910.280 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 691.880 2.400 693.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 474.600 2.400 475.720 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 311.640 2.400 312.760 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 148.680 2.400 149.800 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 536.760 2965.000 537.880 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 703.080 2965.000 704.200 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 869.400 2965.000 870.520 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 1035.720 2965.000 1036.840 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 1257.480 2965.000 1258.600 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 1479.240 2965.000 1480.360 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 1701.000 2965.000 1702.120 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 148.680 2965.000 149.800 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 2033.640 2965.000 2034.760 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 2255.400 2965.000 2256.520 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 2477.160 2965.000 2478.280 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 2698.920 2965.000 2700.040 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 2920.680 2965.000 2921.800 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2664.760 2957.800 2665.880 2965.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2337.720 2957.800 2338.840 2965.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2010.680 2957.800 2011.800 2965.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1683.640 2957.800 1684.760 2965.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1356.600 2957.800 1357.720 2965.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 315.000 2965.000 316.120 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1029.560 2957.800 1030.680 2965.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 702.520 2957.800 703.640 2965.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 375.480 2957.800 376.600 2965.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 48.440 2957.800 49.560 2965.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2756.040 2.400 2757.160 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2538.760 2.400 2539.880 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2321.480 2.400 2322.600 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2104.200 2.400 2105.320 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1886.920 2.400 1888.040 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1669.640 2.400 1670.760 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 481.320 2965.000 482.440 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1452.360 2.400 1453.480 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1235.080 2.400 1236.200 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1017.800 2.400 1018.920 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 800.520 2.400 801.640 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 583.240 2.400 584.360 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 365.960 2.400 367.080 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 203.000 2.400 204.120 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 40.040 2.400 41.160 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 647.640 2965.000 648.760 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 813.960 2965.000 815.080 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 980.280 2965.000 981.400 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 1146.600 2965.000 1147.720 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 1368.360 2965.000 1369.480 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 1590.120 2965.000 1591.240 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 1811.880 2965.000 1813.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 93.240 2965.000 94.360 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 1978.200 2965.000 1979.320 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 2199.960 2965.000 2201.080 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 2421.720 2965.000 2422.840 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 2643.480 2965.000 2644.600 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 2865.240 2965.000 2866.360 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2746.520 2957.800 2747.640 2965.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2419.480 2957.800 2420.600 2965.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2092.440 2957.800 2093.560 2965.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1765.400 2957.800 1766.520 2965.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1438.360 2957.800 1439.480 2965.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 259.560 2965.000 260.680 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1111.320 2957.800 1112.440 2965.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 784.280 2957.800 785.400 2965.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 457.240 2957.800 458.360 2965.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 130.200 2957.800 131.320 2965.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2810.360 2.400 2811.480 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2593.080 2.400 2594.200 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2375.800 2.400 2376.920 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2158.520 2.400 2159.640 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1941.240 2.400 1942.360 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1723.960 2.400 1725.080 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 425.880 2965.000 427.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1506.680 2.400 1507.800 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1289.400 2.400 1290.520 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1072.120 2.400 1073.240 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 854.840 2.400 855.960 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 637.560 2.400 638.680 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 420.280 2.400 421.400 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 257.320 2.400 258.440 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 94.360 2.400 95.480 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 592.200 2965.000 593.320 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 758.520 2965.000 759.640 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 924.840 2965.000 925.960 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 1091.160 2965.000 1092.280 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 1312.920 2965.000 1314.040 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 1534.680 2965.000 1535.800 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2957.800 1756.440 2965.000 1757.560 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 692.440 -4.800 693.560 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2372.440 -4.800 2373.560 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2389.240 -4.800 2390.360 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2406.040 -4.800 2407.160 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2422.840 -4.800 2423.960 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2439.640 -4.800 2440.760 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2456.440 -4.800 2457.560 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2473.240 -4.800 2474.360 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2490.040 -4.800 2491.160 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2506.840 -4.800 2507.960 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2523.640 -4.800 2524.760 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 860.440 -4.800 861.560 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2540.440 -4.800 2541.560 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2557.240 -4.800 2558.360 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2574.040 -4.800 2575.160 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2590.840 -4.800 2591.960 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2607.640 -4.800 2608.760 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2624.440 -4.800 2625.560 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2641.240 -4.800 2642.360 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2658.040 -4.800 2659.160 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2674.840 -4.800 2675.960 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2691.640 -4.800 2692.760 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 877.240 -4.800 878.360 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2708.440 -4.800 2709.560 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2725.240 -4.800 2726.360 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2742.040 -4.800 2743.160 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2758.840 -4.800 2759.960 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2775.640 -4.800 2776.760 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2792.440 -4.800 2793.560 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2809.240 -4.800 2810.360 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2826.040 -4.800 2827.160 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 894.040 -4.800 895.160 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 910.840 -4.800 911.960 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 927.640 -4.800 928.760 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 944.440 -4.800 945.560 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 961.240 -4.800 962.360 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 978.040 -4.800 979.160 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 994.840 -4.800 995.960 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1011.640 -4.800 1012.760 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 709.240 -4.800 710.360 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1028.440 -4.800 1029.560 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1045.240 -4.800 1046.360 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1062.040 -4.800 1063.160 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1078.840 -4.800 1079.960 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1095.640 -4.800 1096.760 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1112.440 -4.800 1113.560 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1129.240 -4.800 1130.360 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1146.040 -4.800 1147.160 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1162.840 -4.800 1163.960 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1179.640 -4.800 1180.760 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 726.040 -4.800 727.160 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1196.440 -4.800 1197.560 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1213.240 -4.800 1214.360 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1230.040 -4.800 1231.160 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1246.840 -4.800 1247.960 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1263.640 -4.800 1264.760 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1280.440 -4.800 1281.560 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1297.240 -4.800 1298.360 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1314.040 -4.800 1315.160 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1330.840 -4.800 1331.960 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1347.640 -4.800 1348.760 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 742.840 -4.800 743.960 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1364.440 -4.800 1365.560 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1381.240 -4.800 1382.360 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1398.040 -4.800 1399.160 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1414.840 -4.800 1415.960 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1431.640 -4.800 1432.760 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1448.440 -4.800 1449.560 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1465.240 -4.800 1466.360 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1482.040 -4.800 1483.160 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1498.840 -4.800 1499.960 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1515.640 -4.800 1516.760 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 759.640 -4.800 760.760 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1532.440 -4.800 1533.560 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1549.240 -4.800 1550.360 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1566.040 -4.800 1567.160 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1582.840 -4.800 1583.960 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1599.640 -4.800 1600.760 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1616.440 -4.800 1617.560 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1633.240 -4.800 1634.360 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1650.040 -4.800 1651.160 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1666.840 -4.800 1667.960 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1683.640 -4.800 1684.760 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 776.440 -4.800 777.560 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1700.440 -4.800 1701.560 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1717.240 -4.800 1718.360 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1734.040 -4.800 1735.160 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1750.840 -4.800 1751.960 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1767.640 -4.800 1768.760 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1784.440 -4.800 1785.560 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1801.240 -4.800 1802.360 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1818.040 -4.800 1819.160 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1834.840 -4.800 1835.960 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1851.640 -4.800 1852.760 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 793.240 -4.800 794.360 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1868.440 -4.800 1869.560 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1885.240 -4.800 1886.360 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1902.040 -4.800 1903.160 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1918.840 -4.800 1919.960 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1935.640 -4.800 1936.760 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1952.440 -4.800 1953.560 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1969.240 -4.800 1970.360 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1986.040 -4.800 1987.160 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2002.840 -4.800 2003.960 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2019.640 -4.800 2020.760 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 810.040 -4.800 811.160 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2036.440 -4.800 2037.560 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2053.240 -4.800 2054.360 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2070.040 -4.800 2071.160 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2086.840 -4.800 2087.960 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2103.640 -4.800 2104.760 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2120.440 -4.800 2121.560 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2137.240 -4.800 2138.360 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2154.040 -4.800 2155.160 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2170.840 -4.800 2171.960 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2187.640 -4.800 2188.760 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 826.840 -4.800 827.960 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2204.440 -4.800 2205.560 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2221.240 -4.800 2222.360 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2238.040 -4.800 2239.160 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2254.840 -4.800 2255.960 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2271.640 -4.800 2272.760 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2288.440 -4.800 2289.560 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2305.240 -4.800 2306.360 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2322.040 -4.800 2323.160 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2338.840 -4.800 2339.960 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2355.640 -4.800 2356.760 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 843.640 -4.800 844.760 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 698.040 -4.800 699.160 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2378.040 -4.800 2379.160 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2394.840 -4.800 2395.960 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2411.640 -4.800 2412.760 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2428.440 -4.800 2429.560 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2445.240 -4.800 2446.360 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2462.040 -4.800 2463.160 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2478.840 -4.800 2479.960 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2495.640 -4.800 2496.760 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2512.440 -4.800 2513.560 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2529.240 -4.800 2530.360 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 866.040 -4.800 867.160 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2546.040 -4.800 2547.160 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2562.840 -4.800 2563.960 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2579.640 -4.800 2580.760 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2596.440 -4.800 2597.560 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2613.240 -4.800 2614.360 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2630.040 -4.800 2631.160 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2646.840 -4.800 2647.960 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2663.640 -4.800 2664.760 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2680.440 -4.800 2681.560 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2697.240 -4.800 2698.360 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 882.840 -4.800 883.960 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2714.040 -4.800 2715.160 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2730.840 -4.800 2731.960 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2747.640 -4.800 2748.760 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2764.440 -4.800 2765.560 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2781.240 -4.800 2782.360 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2798.040 -4.800 2799.160 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2814.840 -4.800 2815.960 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2831.640 -4.800 2832.760 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 899.640 -4.800 900.760 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 916.440 -4.800 917.560 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 933.240 -4.800 934.360 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 950.040 -4.800 951.160 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 966.840 -4.800 967.960 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 983.640 -4.800 984.760 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1000.440 -4.800 1001.560 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1017.240 -4.800 1018.360 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 714.840 -4.800 715.960 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1034.040 -4.800 1035.160 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1050.840 -4.800 1051.960 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1067.640 -4.800 1068.760 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1084.440 -4.800 1085.560 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1101.240 -4.800 1102.360 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1118.040 -4.800 1119.160 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1134.840 -4.800 1135.960 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1151.640 -4.800 1152.760 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1168.440 -4.800 1169.560 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1185.240 -4.800 1186.360 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 731.640 -4.800 732.760 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1202.040 -4.800 1203.160 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1218.840 -4.800 1219.960 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1235.640 -4.800 1236.760 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1252.440 -4.800 1253.560 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1269.240 -4.800 1270.360 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1286.040 -4.800 1287.160 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1302.840 -4.800 1303.960 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1319.640 -4.800 1320.760 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1336.440 -4.800 1337.560 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1353.240 -4.800 1354.360 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 748.440 -4.800 749.560 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1370.040 -4.800 1371.160 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1386.840 -4.800 1387.960 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1403.640 -4.800 1404.760 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1420.440 -4.800 1421.560 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1437.240 -4.800 1438.360 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1454.040 -4.800 1455.160 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1470.840 -4.800 1471.960 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1487.640 -4.800 1488.760 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1504.440 -4.800 1505.560 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1521.240 -4.800 1522.360 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 765.240 -4.800 766.360 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1538.040 -4.800 1539.160 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1554.840 -4.800 1555.960 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1571.640 -4.800 1572.760 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1588.440 -4.800 1589.560 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1605.240 -4.800 1606.360 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1622.040 -4.800 1623.160 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1638.840 -4.800 1639.960 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1655.640 -4.800 1656.760 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1672.440 -4.800 1673.560 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1689.240 -4.800 1690.360 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 782.040 -4.800 783.160 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1706.040 -4.800 1707.160 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1722.840 -4.800 1723.960 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1739.640 -4.800 1740.760 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1756.440 -4.800 1757.560 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1773.240 -4.800 1774.360 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1790.040 -4.800 1791.160 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1806.840 -4.800 1807.960 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1823.640 -4.800 1824.760 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1840.440 -4.800 1841.560 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1857.240 -4.800 1858.360 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 798.840 -4.800 799.960 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1874.040 -4.800 1875.160 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1890.840 -4.800 1891.960 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1907.640 -4.800 1908.760 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1924.440 -4.800 1925.560 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1941.240 -4.800 1942.360 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1958.040 -4.800 1959.160 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1974.840 -4.800 1975.960 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1991.640 -4.800 1992.760 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2008.440 -4.800 2009.560 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2025.240 -4.800 2026.360 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 815.640 -4.800 816.760 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2042.040 -4.800 2043.160 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2058.840 -4.800 2059.960 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2075.640 -4.800 2076.760 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2092.440 -4.800 2093.560 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2109.240 -4.800 2110.360 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2126.040 -4.800 2127.160 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2142.840 -4.800 2143.960 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2159.640 -4.800 2160.760 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2176.440 -4.800 2177.560 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2193.240 -4.800 2194.360 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 832.440 -4.800 833.560 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2210.040 -4.800 2211.160 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2226.840 -4.800 2227.960 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2243.640 -4.800 2244.760 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2260.440 -4.800 2261.560 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2277.240 -4.800 2278.360 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2294.040 -4.800 2295.160 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2310.840 -4.800 2311.960 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2327.640 -4.800 2328.760 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2344.440 -4.800 2345.560 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2361.240 -4.800 2362.360 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 849.240 -4.800 850.360 2.400 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 703.640 -4.800 704.760 2.400 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2383.640 -4.800 2384.760 2.400 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2400.440 -4.800 2401.560 2.400 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2417.240 -4.800 2418.360 2.400 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2434.040 -4.800 2435.160 2.400 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2450.840 -4.800 2451.960 2.400 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2467.640 -4.800 2468.760 2.400 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2484.440 -4.800 2485.560 2.400 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2501.240 -4.800 2502.360 2.400 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2518.040 -4.800 2519.160 2.400 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2534.840 -4.800 2535.960 2.400 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 871.640 -4.800 872.760 2.400 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2551.640 -4.800 2552.760 2.400 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2568.440 -4.800 2569.560 2.400 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2585.240 -4.800 2586.360 2.400 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2602.040 -4.800 2603.160 2.400 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2618.840 -4.800 2619.960 2.400 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2635.640 -4.800 2636.760 2.400 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2652.440 -4.800 2653.560 2.400 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2669.240 -4.800 2670.360 2.400 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2686.040 -4.800 2687.160 2.400 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2702.840 -4.800 2703.960 2.400 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 888.440 -4.800 889.560 2.400 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2719.640 -4.800 2720.760 2.400 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2736.440 -4.800 2737.560 2.400 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2753.240 -4.800 2754.360 2.400 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2770.040 -4.800 2771.160 2.400 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2786.840 -4.800 2787.960 2.400 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2803.640 -4.800 2804.760 2.400 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2820.440 -4.800 2821.560 2.400 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2837.240 -4.800 2838.360 2.400 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 905.240 -4.800 906.360 2.400 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 922.040 -4.800 923.160 2.400 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 938.840 -4.800 939.960 2.400 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 955.640 -4.800 956.760 2.400 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 972.440 -4.800 973.560 2.400 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 989.240 -4.800 990.360 2.400 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1006.040 -4.800 1007.160 2.400 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1022.840 -4.800 1023.960 2.400 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 720.440 -4.800 721.560 2.400 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1039.640 -4.800 1040.760 2.400 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1056.440 -4.800 1057.560 2.400 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1073.240 -4.800 1074.360 2.400 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1090.040 -4.800 1091.160 2.400 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1106.840 -4.800 1107.960 2.400 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1123.640 -4.800 1124.760 2.400 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1140.440 -4.800 1141.560 2.400 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1157.240 -4.800 1158.360 2.400 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1174.040 -4.800 1175.160 2.400 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1190.840 -4.800 1191.960 2.400 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 737.240 -4.800 738.360 2.400 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1207.640 -4.800 1208.760 2.400 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1224.440 -4.800 1225.560 2.400 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1241.240 -4.800 1242.360 2.400 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1258.040 -4.800 1259.160 2.400 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1274.840 -4.800 1275.960 2.400 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1291.640 -4.800 1292.760 2.400 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1308.440 -4.800 1309.560 2.400 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1325.240 -4.800 1326.360 2.400 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1342.040 -4.800 1343.160 2.400 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1358.840 -4.800 1359.960 2.400 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 754.040 -4.800 755.160 2.400 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1375.640 -4.800 1376.760 2.400 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1392.440 -4.800 1393.560 2.400 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1409.240 -4.800 1410.360 2.400 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1426.040 -4.800 1427.160 2.400 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1442.840 -4.800 1443.960 2.400 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1459.640 -4.800 1460.760 2.400 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1476.440 -4.800 1477.560 2.400 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1493.240 -4.800 1494.360 2.400 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1510.040 -4.800 1511.160 2.400 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1526.840 -4.800 1527.960 2.400 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 770.840 -4.800 771.960 2.400 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1543.640 -4.800 1544.760 2.400 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1560.440 -4.800 1561.560 2.400 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1577.240 -4.800 1578.360 2.400 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1594.040 -4.800 1595.160 2.400 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1610.840 -4.800 1611.960 2.400 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1627.640 -4.800 1628.760 2.400 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1644.440 -4.800 1645.560 2.400 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1661.240 -4.800 1662.360 2.400 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1678.040 -4.800 1679.160 2.400 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1694.840 -4.800 1695.960 2.400 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 787.640 -4.800 788.760 2.400 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1711.640 -4.800 1712.760 2.400 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1728.440 -4.800 1729.560 2.400 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1745.240 -4.800 1746.360 2.400 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1762.040 -4.800 1763.160 2.400 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1778.840 -4.800 1779.960 2.400 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1795.640 -4.800 1796.760 2.400 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1812.440 -4.800 1813.560 2.400 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1829.240 -4.800 1830.360 2.400 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1846.040 -4.800 1847.160 2.400 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1862.840 -4.800 1863.960 2.400 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 804.440 -4.800 805.560 2.400 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1879.640 -4.800 1880.760 2.400 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1896.440 -4.800 1897.560 2.400 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1913.240 -4.800 1914.360 2.400 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1930.040 -4.800 1931.160 2.400 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1946.840 -4.800 1947.960 2.400 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1963.640 -4.800 1964.760 2.400 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1980.440 -4.800 1981.560 2.400 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1997.240 -4.800 1998.360 2.400 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2014.040 -4.800 2015.160 2.400 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2030.840 -4.800 2031.960 2.400 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 821.240 -4.800 822.360 2.400 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2047.640 -4.800 2048.760 2.400 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2064.440 -4.800 2065.560 2.400 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2081.240 -4.800 2082.360 2.400 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2098.040 -4.800 2099.160 2.400 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2114.840 -4.800 2115.960 2.400 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2131.640 -4.800 2132.760 2.400 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2148.440 -4.800 2149.560 2.400 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2165.240 -4.800 2166.360 2.400 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2182.040 -4.800 2183.160 2.400 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2198.840 -4.800 2199.960 2.400 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 838.040 -4.800 839.160 2.400 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2215.640 -4.800 2216.760 2.400 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2232.440 -4.800 2233.560 2.400 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2249.240 -4.800 2250.360 2.400 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2266.040 -4.800 2267.160 2.400 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2282.840 -4.800 2283.960 2.400 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2299.640 -4.800 2300.760 2.400 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2316.440 -4.800 2317.560 2.400 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2333.240 -4.800 2334.360 2.400 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2350.040 -4.800 2351.160 2.400 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2366.840 -4.800 2367.960 2.400 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 854.840 -4.800 855.960 2.400 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2842.840 -4.800 2843.960 2.400 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2848.440 -4.800 2849.560 2.400 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2854.040 -4.800 2855.160 2.400 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2859.640 -4.800 2860.760 2.400 ;
    END
  END user_irq[2]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT -4.780 -3.420 -1.680 2986.540 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.780 -3.420 2985.100 -0.320 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.780 2983.440 2985.100 2986.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2982.000 -3.420 2985.100 2986.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 15.770 -8.220 18.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 105.770 -8.220 108.870 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 105.770 2291.710 108.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 195.770 -8.220 198.870 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 195.770 2291.710 198.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 285.770 -8.220 288.870 387.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 285.770 556.190 288.870 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 285.770 2291.710 288.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 375.770 -8.220 378.870 387.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 375.770 556.190 378.870 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 375.770 2291.710 378.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 465.770 -8.220 468.870 387.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 465.770 556.190 468.870 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 465.770 2291.710 468.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 555.770 -8.220 558.870 387.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 555.770 556.190 558.870 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 555.770 2291.710 558.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 645.770 -8.220 648.870 387.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 645.770 556.190 648.870 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 645.770 2291.710 648.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 735.770 -8.220 738.870 387.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 735.770 556.190 738.870 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 735.770 2291.710 738.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 825.770 -8.220 828.870 387.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 825.770 556.190 828.870 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 825.770 2291.710 828.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 915.770 -8.220 918.870 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 915.770 2291.710 918.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1005.770 -8.220 1008.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1095.770 -8.220 1098.870 44.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1095.770 741.710 1098.870 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1095.770 2291.710 1098.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1185.770 -8.220 1188.870 44.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1185.770 741.710 1188.870 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1185.770 2291.710 1188.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1275.770 -8.220 1278.870 44.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1275.770 741.710 1278.870 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1275.770 2291.710 1278.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1365.770 -8.220 1368.870 44.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1365.770 741.710 1368.870 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1365.770 2291.710 1368.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1455.770 -8.220 1458.870 44.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1455.770 741.710 1458.870 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1455.770 2291.710 1458.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1545.770 -8.220 1548.870 44.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1545.770 741.710 1548.870 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1545.770 2291.710 1548.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1635.770 -8.220 1638.870 44.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1635.770 741.710 1638.870 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1635.770 2291.710 1638.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1725.770 -8.220 1728.870 44.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1725.770 741.710 1728.870 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1725.770 2291.710 1728.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1815.770 -8.220 1818.870 44.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1815.770 741.710 1818.870 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1815.770 2291.710 1818.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1905.770 -8.220 1908.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1995.770 -8.220 1998.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2085.770 -8.220 2088.870 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2085.770 2291.710 2088.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2175.770 -8.220 2178.870 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2175.770 2291.710 2178.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2265.770 -8.220 2268.870 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2265.770 2291.710 2268.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2355.770 -8.220 2358.870 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2355.770 2291.710 2358.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2445.770 -8.220 2448.870 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2445.770 2291.710 2448.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2535.770 -8.220 2538.870 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2535.770 2291.710 2538.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2625.770 -8.220 2628.870 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2625.770 2291.710 2628.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2715.770 -8.220 2718.870 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2715.770 2291.710 2718.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2805.770 -8.220 2808.870 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2805.770 2291.710 2808.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2895.770 -8.220 2898.870 2991.340 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 19.130 2989.900 22.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 109.130 2989.900 112.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 199.130 2989.900 202.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 289.130 2989.900 292.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 379.130 2989.900 382.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 469.130 2989.900 472.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 559.130 2989.900 562.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 649.130 2989.900 652.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 739.130 2989.900 742.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 829.130 2989.900 832.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 919.130 2989.900 922.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1009.130 2989.900 1012.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1099.130 2989.900 1102.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1189.130 2989.900 1192.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1279.130 2989.900 1282.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1369.130 2989.900 1372.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1459.130 2989.900 1462.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1549.130 2989.900 1552.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1639.130 2989.900 1642.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1729.130 2989.900 1732.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1819.130 2989.900 1822.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1909.130 2989.900 1912.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1999.130 2989.900 2002.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2089.130 2989.900 2092.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2179.130 2989.900 2182.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2269.130 2989.900 2272.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2359.130 2989.900 2362.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2449.130 2989.900 2452.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2539.130 2989.900 2542.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2629.130 2989.900 2632.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2719.130 2989.900 2722.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2809.130 2989.900 2812.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2899.130 2989.900 2902.230 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT -9.580 -8.220 -6.480 2991.340 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 -8.220 2989.900 -5.120 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2988.240 2989.900 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2986.800 -8.220 2989.900 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 34.370 -8.220 37.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 124.370 -8.220 127.470 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 124.370 1491.710 127.470 1594.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 124.370 2291.710 127.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 214.370 -8.220 217.470 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 214.370 1491.710 217.470 1594.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 214.370 2291.710 217.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 304.370 -8.220 307.470 387.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 304.370 556.190 307.470 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 304.370 1491.710 307.470 1594.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 304.370 2291.710 307.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 394.370 -8.220 397.470 387.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 394.370 556.190 397.470 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 394.370 1491.710 397.470 1594.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 394.370 2291.710 397.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 484.370 -8.220 487.470 387.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 484.370 556.190 487.470 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 484.370 1491.710 487.470 1594.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 484.370 2291.710 487.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 574.370 -8.220 577.470 387.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 574.370 556.190 577.470 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 574.370 1491.710 577.470 1594.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 574.370 2291.710 577.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 664.370 -8.220 667.470 387.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 664.370 556.190 667.470 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 664.370 1491.710 667.470 1594.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 664.370 2291.710 667.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 754.370 -8.220 757.470 387.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 754.370 556.190 757.470 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 754.370 1491.710 757.470 1594.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 754.370 2291.710 757.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 844.370 -8.220 847.470 387.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 844.370 556.190 847.470 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 844.370 1491.710 847.470 1594.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 844.370 2291.710 847.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 934.370 -8.220 937.470 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 934.370 1491.710 937.470 1594.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 934.370 2291.710 937.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1024.370 -8.220 1027.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1114.370 741.710 1117.470 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1114.370 1491.710 1117.470 1594.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1114.370 2291.710 1117.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1204.370 741.710 1207.470 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1204.370 1491.710 1207.470 1594.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1204.370 2291.710 1207.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1294.370 741.710 1297.470 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1294.370 1491.710 1297.470 1594.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1294.370 2291.710 1297.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1384.370 741.710 1387.470 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1384.370 1491.710 1387.470 1594.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1384.370 2291.710 1387.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1474.370 741.710 1477.470 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1474.370 1491.710 1477.470 1594.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1474.370 2291.710 1477.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1564.370 741.710 1567.470 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1564.370 1491.710 1567.470 1594.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1564.370 2291.710 1567.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1654.370 741.710 1657.470 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1654.370 1491.710 1657.470 1594.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1654.370 2291.710 1657.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1744.370 741.710 1747.470 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1744.370 1491.710 1747.470 1594.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1744.370 2291.710 1747.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1834.370 741.710 1837.470 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1834.370 1491.710 1837.470 1594.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1834.370 2291.710 1837.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1924.370 -8.220 1927.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2014.370 -8.220 2017.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2104.370 -8.220 2107.470 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2104.370 1491.710 2107.470 1594.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2104.370 2291.710 2107.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2194.370 -8.220 2197.470 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2194.370 1491.710 2197.470 1594.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2194.370 2291.710 2197.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2284.370 -8.220 2287.470 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2284.370 1491.710 2287.470 1594.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2284.370 2291.710 2287.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2374.370 -8.220 2377.470 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2374.370 1491.710 2377.470 1594.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2374.370 2291.710 2377.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2464.370 -8.220 2467.470 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2464.370 1491.710 2467.470 1594.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2464.370 2291.710 2467.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2554.370 -8.220 2557.470 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2554.370 1491.710 2557.470 1594.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2554.370 2291.710 2557.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2644.370 -8.220 2647.470 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2644.370 1491.710 2647.470 1594.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2644.370 2291.710 2647.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2734.370 -8.220 2737.470 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2734.370 1491.710 2737.470 1594.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2734.370 2291.710 2737.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2824.370 -8.220 2827.470 794.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2824.370 1491.710 2827.470 1594.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2824.370 2291.710 2827.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2914.370 -8.220 2917.470 2991.340 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 49.130 2989.900 52.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 139.130 2989.900 142.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 229.130 2989.900 232.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 319.130 2989.900 322.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 409.130 2989.900 412.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 499.130 2989.900 502.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 589.130 2989.900 592.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 679.130 2989.900 682.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 769.130 2989.900 772.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 859.130 2989.900 862.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 949.130 2989.900 952.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1039.130 2989.900 1042.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1129.130 2989.900 1132.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1219.130 2989.900 1222.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1309.130 2989.900 1312.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1399.130 2989.900 1402.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1489.130 2989.900 1492.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1579.130 2989.900 1582.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1669.130 2989.900 1672.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1759.130 2989.900 1762.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1849.130 2989.900 1852.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1939.130 2989.900 1942.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2029.130 2989.900 2032.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2119.130 2989.900 2122.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2209.130 2989.900 2212.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2299.130 2989.900 2302.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2389.130 2989.900 2392.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2479.130 2989.900 2482.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2569.130 2989.900 2572.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2659.130 2989.900 2662.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2749.130 2989.900 2752.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2839.130 2989.900 2842.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2929.130 2989.900 2932.230 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 98.840 -4.800 99.960 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 104.440 -4.800 105.560 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 110.040 -4.800 111.160 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 132.440 -4.800 133.560 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 322.840 -4.800 323.960 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 339.640 -4.800 340.760 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 356.440 -4.800 357.560 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 373.240 -4.800 374.360 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 390.040 -4.800 391.160 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 406.840 -4.800 407.960 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 423.640 -4.800 424.760 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 440.440 -4.800 441.560 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 457.240 -4.800 458.360 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 474.040 -4.800 475.160 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 154.840 -4.800 155.960 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 490.840 -4.800 491.960 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 507.640 -4.800 508.760 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 524.440 -4.800 525.560 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 541.240 -4.800 542.360 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 558.040 -4.800 559.160 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 574.840 -4.800 575.960 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 591.640 -4.800 592.760 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 608.440 -4.800 609.560 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 625.240 -4.800 626.360 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 642.040 -4.800 643.160 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 177.240 -4.800 178.360 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 658.840 -4.800 659.960 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 675.640 -4.800 676.760 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 199.640 -4.800 200.760 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 222.040 -4.800 223.160 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 238.840 -4.800 239.960 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 255.640 -4.800 256.760 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 272.440 -4.800 273.560 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 289.240 -4.800 290.360 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 306.040 -4.800 307.160 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 115.640 -4.800 116.760 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 138.040 -4.800 139.160 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 328.440 -4.800 329.560 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 345.240 -4.800 346.360 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 362.040 -4.800 363.160 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 378.840 -4.800 379.960 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 395.640 -4.800 396.760 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 412.440 -4.800 413.560 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 429.240 -4.800 430.360 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 446.040 -4.800 447.160 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 462.840 -4.800 463.960 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 479.640 -4.800 480.760 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 160.440 -4.800 161.560 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 496.440 -4.800 497.560 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 513.240 -4.800 514.360 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 530.040 -4.800 531.160 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 546.840 -4.800 547.960 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 563.640 -4.800 564.760 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 580.440 -4.800 581.560 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 597.240 -4.800 598.360 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 614.040 -4.800 615.160 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 630.840 -4.800 631.960 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 647.640 -4.800 648.760 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 182.840 -4.800 183.960 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 664.440 -4.800 665.560 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 681.240 -4.800 682.360 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 205.240 -4.800 206.360 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 227.640 -4.800 228.760 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 244.440 -4.800 245.560 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 261.240 -4.800 262.360 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 278.040 -4.800 279.160 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 294.840 -4.800 295.960 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 311.640 -4.800 312.760 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 143.640 -4.800 144.760 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 334.040 -4.800 335.160 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 350.840 -4.800 351.960 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 367.640 -4.800 368.760 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 384.440 -4.800 385.560 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 401.240 -4.800 402.360 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 418.040 -4.800 419.160 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 434.840 -4.800 435.960 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 451.640 -4.800 452.760 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 468.440 -4.800 469.560 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 485.240 -4.800 486.360 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 166.040 -4.800 167.160 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 502.040 -4.800 503.160 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 518.840 -4.800 519.960 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 535.640 -4.800 536.760 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 552.440 -4.800 553.560 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 569.240 -4.800 570.360 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 586.040 -4.800 587.160 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 602.840 -4.800 603.960 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 619.640 -4.800 620.760 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 636.440 -4.800 637.560 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 653.240 -4.800 654.360 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 188.440 -4.800 189.560 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 670.040 -4.800 671.160 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 686.840 -4.800 687.960 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 210.840 -4.800 211.960 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 233.240 -4.800 234.360 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 250.040 -4.800 251.160 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 266.840 -4.800 267.960 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 283.640 -4.800 284.760 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 300.440 -4.800 301.560 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 317.240 -4.800 318.360 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 149.240 -4.800 150.360 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 171.640 -4.800 172.760 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 194.040 -4.800 195.160 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 216.440 -4.800 217.560 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 121.240 -4.800 122.360 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 126.840 -4.800 127.960 2.400 ;
    END
  END wbs_we_i
  OBS
      LAYER Metal1 ;
        RECT 51.720 65.380 2888.200 2301.980 ;
      LAYER Metal2 ;
        RECT 0.140 2957.500 48.140 2958.340 ;
        RECT 49.860 2957.500 129.900 2958.340 ;
        RECT 131.620 2957.500 211.660 2958.340 ;
        RECT 213.380 2957.500 293.420 2958.340 ;
        RECT 295.140 2957.500 375.180 2958.340 ;
        RECT 376.900 2957.500 456.940 2958.340 ;
        RECT 458.660 2957.500 538.700 2958.340 ;
        RECT 540.420 2957.500 620.460 2958.340 ;
        RECT 622.180 2957.500 702.220 2958.340 ;
        RECT 703.940 2957.500 783.980 2958.340 ;
        RECT 785.700 2957.500 865.740 2958.340 ;
        RECT 867.460 2957.500 947.500 2958.340 ;
        RECT 949.220 2957.500 1029.260 2958.340 ;
        RECT 1030.980 2957.500 1111.020 2958.340 ;
        RECT 1112.740 2957.500 1192.780 2958.340 ;
        RECT 1194.500 2957.500 1274.540 2958.340 ;
        RECT 1276.260 2957.500 1356.300 2958.340 ;
        RECT 1358.020 2957.500 1438.060 2958.340 ;
        RECT 1439.780 2957.500 1519.820 2958.340 ;
        RECT 1521.540 2957.500 1601.580 2958.340 ;
        RECT 1603.300 2957.500 1683.340 2958.340 ;
        RECT 1685.060 2957.500 1765.100 2958.340 ;
        RECT 1766.820 2957.500 1846.860 2958.340 ;
        RECT 1848.580 2957.500 1928.620 2958.340 ;
        RECT 1930.340 2957.500 2010.380 2958.340 ;
        RECT 2012.100 2957.500 2092.140 2958.340 ;
        RECT 2093.860 2957.500 2173.900 2958.340 ;
        RECT 2175.620 2957.500 2255.660 2958.340 ;
        RECT 2257.380 2957.500 2337.420 2958.340 ;
        RECT 2339.140 2957.500 2419.180 2958.340 ;
        RECT 2420.900 2957.500 2500.940 2958.340 ;
        RECT 2502.660 2957.500 2582.700 2958.340 ;
        RECT 2584.420 2957.500 2664.460 2958.340 ;
        RECT 2666.180 2957.500 2746.220 2958.340 ;
        RECT 2747.940 2957.500 2827.980 2958.340 ;
        RECT 2829.700 2957.500 2909.740 2958.340 ;
        RECT 2911.460 2957.500 2950.500 2958.340 ;
        RECT 0.140 2.700 2950.500 2957.500 ;
        RECT 0.140 1.820 98.540 2.700 ;
        RECT 100.260 1.820 104.140 2.700 ;
        RECT 105.860 1.820 109.740 2.700 ;
        RECT 111.460 1.820 115.340 2.700 ;
        RECT 117.060 1.820 120.940 2.700 ;
        RECT 122.660 1.820 126.540 2.700 ;
        RECT 128.260 1.820 132.140 2.700 ;
        RECT 133.860 1.820 137.740 2.700 ;
        RECT 139.460 1.820 143.340 2.700 ;
        RECT 145.060 1.820 148.940 2.700 ;
        RECT 150.660 1.820 154.540 2.700 ;
        RECT 156.260 1.820 160.140 2.700 ;
        RECT 161.860 1.820 165.740 2.700 ;
        RECT 167.460 1.820 171.340 2.700 ;
        RECT 173.060 1.820 176.940 2.700 ;
        RECT 178.660 1.820 182.540 2.700 ;
        RECT 184.260 1.820 188.140 2.700 ;
        RECT 189.860 1.820 193.740 2.700 ;
        RECT 195.460 1.820 199.340 2.700 ;
        RECT 201.060 1.820 204.940 2.700 ;
        RECT 206.660 1.820 210.540 2.700 ;
        RECT 212.260 1.820 216.140 2.700 ;
        RECT 217.860 1.820 221.740 2.700 ;
        RECT 223.460 1.820 227.340 2.700 ;
        RECT 229.060 1.820 232.940 2.700 ;
        RECT 234.660 1.820 238.540 2.700 ;
        RECT 240.260 1.820 244.140 2.700 ;
        RECT 245.860 1.820 249.740 2.700 ;
        RECT 251.460 1.820 255.340 2.700 ;
        RECT 257.060 1.820 260.940 2.700 ;
        RECT 262.660 1.820 266.540 2.700 ;
        RECT 268.260 1.820 272.140 2.700 ;
        RECT 273.860 1.820 277.740 2.700 ;
        RECT 279.460 1.820 283.340 2.700 ;
        RECT 285.060 1.820 288.940 2.700 ;
        RECT 290.660 1.820 294.540 2.700 ;
        RECT 296.260 1.820 300.140 2.700 ;
        RECT 301.860 1.820 305.740 2.700 ;
        RECT 307.460 1.820 311.340 2.700 ;
        RECT 313.060 1.820 316.940 2.700 ;
        RECT 318.660 1.820 322.540 2.700 ;
        RECT 324.260 1.820 328.140 2.700 ;
        RECT 329.860 1.820 333.740 2.700 ;
        RECT 335.460 1.820 339.340 2.700 ;
        RECT 341.060 1.820 344.940 2.700 ;
        RECT 346.660 1.820 350.540 2.700 ;
        RECT 352.260 1.820 356.140 2.700 ;
        RECT 357.860 1.820 361.740 2.700 ;
        RECT 363.460 1.820 367.340 2.700 ;
        RECT 369.060 1.820 372.940 2.700 ;
        RECT 374.660 1.820 378.540 2.700 ;
        RECT 380.260 1.820 384.140 2.700 ;
        RECT 385.860 1.820 389.740 2.700 ;
        RECT 391.460 1.820 395.340 2.700 ;
        RECT 397.060 1.820 400.940 2.700 ;
        RECT 402.660 1.820 406.540 2.700 ;
        RECT 408.260 1.820 412.140 2.700 ;
        RECT 413.860 1.820 417.740 2.700 ;
        RECT 419.460 1.820 423.340 2.700 ;
        RECT 425.060 1.820 428.940 2.700 ;
        RECT 430.660 1.820 434.540 2.700 ;
        RECT 436.260 1.820 440.140 2.700 ;
        RECT 441.860 1.820 445.740 2.700 ;
        RECT 447.460 1.820 451.340 2.700 ;
        RECT 453.060 1.820 456.940 2.700 ;
        RECT 458.660 1.820 462.540 2.700 ;
        RECT 464.260 1.820 468.140 2.700 ;
        RECT 469.860 1.820 473.740 2.700 ;
        RECT 475.460 1.820 479.340 2.700 ;
        RECT 481.060 1.820 484.940 2.700 ;
        RECT 486.660 1.820 490.540 2.700 ;
        RECT 492.260 1.820 496.140 2.700 ;
        RECT 497.860 1.820 501.740 2.700 ;
        RECT 503.460 1.820 507.340 2.700 ;
        RECT 509.060 1.820 512.940 2.700 ;
        RECT 514.660 1.820 518.540 2.700 ;
        RECT 520.260 1.820 524.140 2.700 ;
        RECT 525.860 1.820 529.740 2.700 ;
        RECT 531.460 1.820 535.340 2.700 ;
        RECT 537.060 1.820 540.940 2.700 ;
        RECT 542.660 1.820 546.540 2.700 ;
        RECT 548.260 1.820 552.140 2.700 ;
        RECT 553.860 1.820 557.740 2.700 ;
        RECT 559.460 1.820 563.340 2.700 ;
        RECT 565.060 1.820 568.940 2.700 ;
        RECT 570.660 1.820 574.540 2.700 ;
        RECT 576.260 1.820 580.140 2.700 ;
        RECT 581.860 1.820 585.740 2.700 ;
        RECT 587.460 1.820 591.340 2.700 ;
        RECT 593.060 1.820 596.940 2.700 ;
        RECT 598.660 1.820 602.540 2.700 ;
        RECT 604.260 1.820 608.140 2.700 ;
        RECT 609.860 1.820 613.740 2.700 ;
        RECT 615.460 1.820 619.340 2.700 ;
        RECT 621.060 1.820 624.940 2.700 ;
        RECT 626.660 1.820 630.540 2.700 ;
        RECT 632.260 1.820 636.140 2.700 ;
        RECT 637.860 1.820 641.740 2.700 ;
        RECT 643.460 1.820 647.340 2.700 ;
        RECT 649.060 1.820 652.940 2.700 ;
        RECT 654.660 1.820 658.540 2.700 ;
        RECT 660.260 1.820 664.140 2.700 ;
        RECT 665.860 1.820 669.740 2.700 ;
        RECT 671.460 1.820 675.340 2.700 ;
        RECT 677.060 1.820 680.940 2.700 ;
        RECT 682.660 1.820 686.540 2.700 ;
        RECT 688.260 1.820 692.140 2.700 ;
        RECT 693.860 1.820 697.740 2.700 ;
        RECT 699.460 1.820 703.340 2.700 ;
        RECT 705.060 1.820 708.940 2.700 ;
        RECT 710.660 1.820 714.540 2.700 ;
        RECT 716.260 1.820 720.140 2.700 ;
        RECT 721.860 1.820 725.740 2.700 ;
        RECT 727.460 1.820 731.340 2.700 ;
        RECT 733.060 1.820 736.940 2.700 ;
        RECT 738.660 1.820 742.540 2.700 ;
        RECT 744.260 1.820 748.140 2.700 ;
        RECT 749.860 1.820 753.740 2.700 ;
        RECT 755.460 1.820 759.340 2.700 ;
        RECT 761.060 1.820 764.940 2.700 ;
        RECT 766.660 1.820 770.540 2.700 ;
        RECT 772.260 1.820 776.140 2.700 ;
        RECT 777.860 1.820 781.740 2.700 ;
        RECT 783.460 1.820 787.340 2.700 ;
        RECT 789.060 1.820 792.940 2.700 ;
        RECT 794.660 1.820 798.540 2.700 ;
        RECT 800.260 1.820 804.140 2.700 ;
        RECT 805.860 1.820 809.740 2.700 ;
        RECT 811.460 1.820 815.340 2.700 ;
        RECT 817.060 1.820 820.940 2.700 ;
        RECT 822.660 1.820 826.540 2.700 ;
        RECT 828.260 1.820 832.140 2.700 ;
        RECT 833.860 1.820 837.740 2.700 ;
        RECT 839.460 1.820 843.340 2.700 ;
        RECT 845.060 1.820 848.940 2.700 ;
        RECT 850.660 1.820 854.540 2.700 ;
        RECT 856.260 1.820 860.140 2.700 ;
        RECT 861.860 1.820 865.740 2.700 ;
        RECT 867.460 1.820 871.340 2.700 ;
        RECT 873.060 1.820 876.940 2.700 ;
        RECT 878.660 1.820 882.540 2.700 ;
        RECT 884.260 1.820 888.140 2.700 ;
        RECT 889.860 1.820 893.740 2.700 ;
        RECT 895.460 1.820 899.340 2.700 ;
        RECT 901.060 1.820 904.940 2.700 ;
        RECT 906.660 1.820 910.540 2.700 ;
        RECT 912.260 1.820 916.140 2.700 ;
        RECT 917.860 1.820 921.740 2.700 ;
        RECT 923.460 1.820 927.340 2.700 ;
        RECT 929.060 1.820 932.940 2.700 ;
        RECT 934.660 1.820 938.540 2.700 ;
        RECT 940.260 1.820 944.140 2.700 ;
        RECT 945.860 1.820 949.740 2.700 ;
        RECT 951.460 1.820 955.340 2.700 ;
        RECT 957.060 1.820 960.940 2.700 ;
        RECT 962.660 1.820 966.540 2.700 ;
        RECT 968.260 1.820 972.140 2.700 ;
        RECT 973.860 1.820 977.740 2.700 ;
        RECT 979.460 1.820 983.340 2.700 ;
        RECT 985.060 1.820 988.940 2.700 ;
        RECT 990.660 1.820 994.540 2.700 ;
        RECT 996.260 1.820 1000.140 2.700 ;
        RECT 1001.860 1.820 1005.740 2.700 ;
        RECT 1007.460 1.820 1011.340 2.700 ;
        RECT 1013.060 1.820 1016.940 2.700 ;
        RECT 1018.660 1.820 1022.540 2.700 ;
        RECT 1024.260 1.820 1028.140 2.700 ;
        RECT 1029.860 1.820 1033.740 2.700 ;
        RECT 1035.460 1.820 1039.340 2.700 ;
        RECT 1041.060 1.820 1044.940 2.700 ;
        RECT 1046.660 1.820 1050.540 2.700 ;
        RECT 1052.260 1.820 1056.140 2.700 ;
        RECT 1057.860 1.820 1061.740 2.700 ;
        RECT 1063.460 1.820 1067.340 2.700 ;
        RECT 1069.060 1.820 1072.940 2.700 ;
        RECT 1074.660 1.820 1078.540 2.700 ;
        RECT 1080.260 1.820 1084.140 2.700 ;
        RECT 1085.860 1.820 1089.740 2.700 ;
        RECT 1091.460 1.820 1095.340 2.700 ;
        RECT 1097.060 1.820 1100.940 2.700 ;
        RECT 1102.660 1.820 1106.540 2.700 ;
        RECT 1108.260 1.820 1112.140 2.700 ;
        RECT 1113.860 1.820 1117.740 2.700 ;
        RECT 1119.460 1.820 1123.340 2.700 ;
        RECT 1125.060 1.820 1128.940 2.700 ;
        RECT 1130.660 1.820 1134.540 2.700 ;
        RECT 1136.260 1.820 1140.140 2.700 ;
        RECT 1141.860 1.820 1145.740 2.700 ;
        RECT 1147.460 1.820 1151.340 2.700 ;
        RECT 1153.060 1.820 1156.940 2.700 ;
        RECT 1158.660 1.820 1162.540 2.700 ;
        RECT 1164.260 1.820 1168.140 2.700 ;
        RECT 1169.860 1.820 1173.740 2.700 ;
        RECT 1175.460 1.820 1179.340 2.700 ;
        RECT 1181.060 1.820 1184.940 2.700 ;
        RECT 1186.660 1.820 1190.540 2.700 ;
        RECT 1192.260 1.820 1196.140 2.700 ;
        RECT 1197.860 1.820 1201.740 2.700 ;
        RECT 1203.460 1.820 1207.340 2.700 ;
        RECT 1209.060 1.820 1212.940 2.700 ;
        RECT 1214.660 1.820 1218.540 2.700 ;
        RECT 1220.260 1.820 1224.140 2.700 ;
        RECT 1225.860 1.820 1229.740 2.700 ;
        RECT 1231.460 1.820 1235.340 2.700 ;
        RECT 1237.060 1.820 1240.940 2.700 ;
        RECT 1242.660 1.820 1246.540 2.700 ;
        RECT 1248.260 1.820 1252.140 2.700 ;
        RECT 1253.860 1.820 1257.740 2.700 ;
        RECT 1259.460 1.820 1263.340 2.700 ;
        RECT 1265.060 1.820 1268.940 2.700 ;
        RECT 1270.660 1.820 1274.540 2.700 ;
        RECT 1276.260 1.820 1280.140 2.700 ;
        RECT 1281.860 1.820 1285.740 2.700 ;
        RECT 1287.460 1.820 1291.340 2.700 ;
        RECT 1293.060 1.820 1296.940 2.700 ;
        RECT 1298.660 1.820 1302.540 2.700 ;
        RECT 1304.260 1.820 1308.140 2.700 ;
        RECT 1309.860 1.820 1313.740 2.700 ;
        RECT 1315.460 1.820 1319.340 2.700 ;
        RECT 1321.060 1.820 1324.940 2.700 ;
        RECT 1326.660 1.820 1330.540 2.700 ;
        RECT 1332.260 1.820 1336.140 2.700 ;
        RECT 1337.860 1.820 1341.740 2.700 ;
        RECT 1343.460 1.820 1347.340 2.700 ;
        RECT 1349.060 1.820 1352.940 2.700 ;
        RECT 1354.660 1.820 1358.540 2.700 ;
        RECT 1360.260 1.820 1364.140 2.700 ;
        RECT 1365.860 1.820 1369.740 2.700 ;
        RECT 1371.460 1.820 1375.340 2.700 ;
        RECT 1377.060 1.820 1380.940 2.700 ;
        RECT 1382.660 1.820 1386.540 2.700 ;
        RECT 1388.260 1.820 1392.140 2.700 ;
        RECT 1393.860 1.820 1397.740 2.700 ;
        RECT 1399.460 1.820 1403.340 2.700 ;
        RECT 1405.060 1.820 1408.940 2.700 ;
        RECT 1410.660 1.820 1414.540 2.700 ;
        RECT 1416.260 1.820 1420.140 2.700 ;
        RECT 1421.860 1.820 1425.740 2.700 ;
        RECT 1427.460 1.820 1431.340 2.700 ;
        RECT 1433.060 1.820 1436.940 2.700 ;
        RECT 1438.660 1.820 1442.540 2.700 ;
        RECT 1444.260 1.820 1448.140 2.700 ;
        RECT 1449.860 1.820 1453.740 2.700 ;
        RECT 1455.460 1.820 1459.340 2.700 ;
        RECT 1461.060 1.820 1464.940 2.700 ;
        RECT 1466.660 1.820 1470.540 2.700 ;
        RECT 1472.260 1.820 1476.140 2.700 ;
        RECT 1477.860 1.820 1481.740 2.700 ;
        RECT 1483.460 1.820 1487.340 2.700 ;
        RECT 1489.060 1.820 1492.940 2.700 ;
        RECT 1494.660 1.820 1498.540 2.700 ;
        RECT 1500.260 1.820 1504.140 2.700 ;
        RECT 1505.860 1.820 1509.740 2.700 ;
        RECT 1511.460 1.820 1515.340 2.700 ;
        RECT 1517.060 1.820 1520.940 2.700 ;
        RECT 1522.660 1.820 1526.540 2.700 ;
        RECT 1528.260 1.820 1532.140 2.700 ;
        RECT 1533.860 1.820 1537.740 2.700 ;
        RECT 1539.460 1.820 1543.340 2.700 ;
        RECT 1545.060 1.820 1548.940 2.700 ;
        RECT 1550.660 1.820 1554.540 2.700 ;
        RECT 1556.260 1.820 1560.140 2.700 ;
        RECT 1561.860 1.820 1565.740 2.700 ;
        RECT 1567.460 1.820 1571.340 2.700 ;
        RECT 1573.060 1.820 1576.940 2.700 ;
        RECT 1578.660 1.820 1582.540 2.700 ;
        RECT 1584.260 1.820 1588.140 2.700 ;
        RECT 1589.860 1.820 1593.740 2.700 ;
        RECT 1595.460 1.820 1599.340 2.700 ;
        RECT 1601.060 1.820 1604.940 2.700 ;
        RECT 1606.660 1.820 1610.540 2.700 ;
        RECT 1612.260 1.820 1616.140 2.700 ;
        RECT 1617.860 1.820 1621.740 2.700 ;
        RECT 1623.460 1.820 1627.340 2.700 ;
        RECT 1629.060 1.820 1632.940 2.700 ;
        RECT 1634.660 1.820 1638.540 2.700 ;
        RECT 1640.260 1.820 1644.140 2.700 ;
        RECT 1645.860 1.820 1649.740 2.700 ;
        RECT 1651.460 1.820 1655.340 2.700 ;
        RECT 1657.060 1.820 1660.940 2.700 ;
        RECT 1662.660 1.820 1666.540 2.700 ;
        RECT 1668.260 1.820 1672.140 2.700 ;
        RECT 1673.860 1.820 1677.740 2.700 ;
        RECT 1679.460 1.820 1683.340 2.700 ;
        RECT 1685.060 1.820 1688.940 2.700 ;
        RECT 1690.660 1.820 1694.540 2.700 ;
        RECT 1696.260 1.820 1700.140 2.700 ;
        RECT 1701.860 1.820 1705.740 2.700 ;
        RECT 1707.460 1.820 1711.340 2.700 ;
        RECT 1713.060 1.820 1716.940 2.700 ;
        RECT 1718.660 1.820 1722.540 2.700 ;
        RECT 1724.260 1.820 1728.140 2.700 ;
        RECT 1729.860 1.820 1733.740 2.700 ;
        RECT 1735.460 1.820 1739.340 2.700 ;
        RECT 1741.060 1.820 1744.940 2.700 ;
        RECT 1746.660 1.820 1750.540 2.700 ;
        RECT 1752.260 1.820 1756.140 2.700 ;
        RECT 1757.860 1.820 1761.740 2.700 ;
        RECT 1763.460 1.820 1767.340 2.700 ;
        RECT 1769.060 1.820 1772.940 2.700 ;
        RECT 1774.660 1.820 1778.540 2.700 ;
        RECT 1780.260 1.820 1784.140 2.700 ;
        RECT 1785.860 1.820 1789.740 2.700 ;
        RECT 1791.460 1.820 1795.340 2.700 ;
        RECT 1797.060 1.820 1800.940 2.700 ;
        RECT 1802.660 1.820 1806.540 2.700 ;
        RECT 1808.260 1.820 1812.140 2.700 ;
        RECT 1813.860 1.820 1817.740 2.700 ;
        RECT 1819.460 1.820 1823.340 2.700 ;
        RECT 1825.060 1.820 1828.940 2.700 ;
        RECT 1830.660 1.820 1834.540 2.700 ;
        RECT 1836.260 1.820 1840.140 2.700 ;
        RECT 1841.860 1.820 1845.740 2.700 ;
        RECT 1847.460 1.820 1851.340 2.700 ;
        RECT 1853.060 1.820 1856.940 2.700 ;
        RECT 1858.660 1.820 1862.540 2.700 ;
        RECT 1864.260 1.820 1868.140 2.700 ;
        RECT 1869.860 1.820 1873.740 2.700 ;
        RECT 1875.460 1.820 1879.340 2.700 ;
        RECT 1881.060 1.820 1884.940 2.700 ;
        RECT 1886.660 1.820 1890.540 2.700 ;
        RECT 1892.260 1.820 1896.140 2.700 ;
        RECT 1897.860 1.820 1901.740 2.700 ;
        RECT 1903.460 1.820 1907.340 2.700 ;
        RECT 1909.060 1.820 1912.940 2.700 ;
        RECT 1914.660 1.820 1918.540 2.700 ;
        RECT 1920.260 1.820 1924.140 2.700 ;
        RECT 1925.860 1.820 1929.740 2.700 ;
        RECT 1931.460 1.820 1935.340 2.700 ;
        RECT 1937.060 1.820 1940.940 2.700 ;
        RECT 1942.660 1.820 1946.540 2.700 ;
        RECT 1948.260 1.820 1952.140 2.700 ;
        RECT 1953.860 1.820 1957.740 2.700 ;
        RECT 1959.460 1.820 1963.340 2.700 ;
        RECT 1965.060 1.820 1968.940 2.700 ;
        RECT 1970.660 1.820 1974.540 2.700 ;
        RECT 1976.260 1.820 1980.140 2.700 ;
        RECT 1981.860 1.820 1985.740 2.700 ;
        RECT 1987.460 1.820 1991.340 2.700 ;
        RECT 1993.060 1.820 1996.940 2.700 ;
        RECT 1998.660 1.820 2002.540 2.700 ;
        RECT 2004.260 1.820 2008.140 2.700 ;
        RECT 2009.860 1.820 2013.740 2.700 ;
        RECT 2015.460 1.820 2019.340 2.700 ;
        RECT 2021.060 1.820 2024.940 2.700 ;
        RECT 2026.660 1.820 2030.540 2.700 ;
        RECT 2032.260 1.820 2036.140 2.700 ;
        RECT 2037.860 1.820 2041.740 2.700 ;
        RECT 2043.460 1.820 2047.340 2.700 ;
        RECT 2049.060 1.820 2052.940 2.700 ;
        RECT 2054.660 1.820 2058.540 2.700 ;
        RECT 2060.260 1.820 2064.140 2.700 ;
        RECT 2065.860 1.820 2069.740 2.700 ;
        RECT 2071.460 1.820 2075.340 2.700 ;
        RECT 2077.060 1.820 2080.940 2.700 ;
        RECT 2082.660 1.820 2086.540 2.700 ;
        RECT 2088.260 1.820 2092.140 2.700 ;
        RECT 2093.860 1.820 2097.740 2.700 ;
        RECT 2099.460 1.820 2103.340 2.700 ;
        RECT 2105.060 1.820 2108.940 2.700 ;
        RECT 2110.660 1.820 2114.540 2.700 ;
        RECT 2116.260 1.820 2120.140 2.700 ;
        RECT 2121.860 1.820 2125.740 2.700 ;
        RECT 2127.460 1.820 2131.340 2.700 ;
        RECT 2133.060 1.820 2136.940 2.700 ;
        RECT 2138.660 1.820 2142.540 2.700 ;
        RECT 2144.260 1.820 2148.140 2.700 ;
        RECT 2149.860 1.820 2153.740 2.700 ;
        RECT 2155.460 1.820 2159.340 2.700 ;
        RECT 2161.060 1.820 2164.940 2.700 ;
        RECT 2166.660 1.820 2170.540 2.700 ;
        RECT 2172.260 1.820 2176.140 2.700 ;
        RECT 2177.860 1.820 2181.740 2.700 ;
        RECT 2183.460 1.820 2187.340 2.700 ;
        RECT 2189.060 1.820 2192.940 2.700 ;
        RECT 2194.660 1.820 2198.540 2.700 ;
        RECT 2200.260 1.820 2204.140 2.700 ;
        RECT 2205.860 1.820 2209.740 2.700 ;
        RECT 2211.460 1.820 2215.340 2.700 ;
        RECT 2217.060 1.820 2220.940 2.700 ;
        RECT 2222.660 1.820 2226.540 2.700 ;
        RECT 2228.260 1.820 2232.140 2.700 ;
        RECT 2233.860 1.820 2237.740 2.700 ;
        RECT 2239.460 1.820 2243.340 2.700 ;
        RECT 2245.060 1.820 2248.940 2.700 ;
        RECT 2250.660 1.820 2254.540 2.700 ;
        RECT 2256.260 1.820 2260.140 2.700 ;
        RECT 2261.860 1.820 2265.740 2.700 ;
        RECT 2267.460 1.820 2271.340 2.700 ;
        RECT 2273.060 1.820 2276.940 2.700 ;
        RECT 2278.660 1.820 2282.540 2.700 ;
        RECT 2284.260 1.820 2288.140 2.700 ;
        RECT 2289.860 1.820 2293.740 2.700 ;
        RECT 2295.460 1.820 2299.340 2.700 ;
        RECT 2301.060 1.820 2304.940 2.700 ;
        RECT 2306.660 1.820 2310.540 2.700 ;
        RECT 2312.260 1.820 2316.140 2.700 ;
        RECT 2317.860 1.820 2321.740 2.700 ;
        RECT 2323.460 1.820 2327.340 2.700 ;
        RECT 2329.060 1.820 2332.940 2.700 ;
        RECT 2334.660 1.820 2338.540 2.700 ;
        RECT 2340.260 1.820 2344.140 2.700 ;
        RECT 2345.860 1.820 2349.740 2.700 ;
        RECT 2351.460 1.820 2355.340 2.700 ;
        RECT 2357.060 1.820 2360.940 2.700 ;
        RECT 2362.660 1.820 2366.540 2.700 ;
        RECT 2368.260 1.820 2372.140 2.700 ;
        RECT 2373.860 1.820 2377.740 2.700 ;
        RECT 2379.460 1.820 2383.340 2.700 ;
        RECT 2385.060 1.820 2388.940 2.700 ;
        RECT 2390.660 1.820 2394.540 2.700 ;
        RECT 2396.260 1.820 2400.140 2.700 ;
        RECT 2401.860 1.820 2405.740 2.700 ;
        RECT 2407.460 1.820 2411.340 2.700 ;
        RECT 2413.060 1.820 2416.940 2.700 ;
        RECT 2418.660 1.820 2422.540 2.700 ;
        RECT 2424.260 1.820 2428.140 2.700 ;
        RECT 2429.860 1.820 2433.740 2.700 ;
        RECT 2435.460 1.820 2439.340 2.700 ;
        RECT 2441.060 1.820 2444.940 2.700 ;
        RECT 2446.660 1.820 2450.540 2.700 ;
        RECT 2452.260 1.820 2456.140 2.700 ;
        RECT 2457.860 1.820 2461.740 2.700 ;
        RECT 2463.460 1.820 2467.340 2.700 ;
        RECT 2469.060 1.820 2472.940 2.700 ;
        RECT 2474.660 1.820 2478.540 2.700 ;
        RECT 2480.260 1.820 2484.140 2.700 ;
        RECT 2485.860 1.820 2489.740 2.700 ;
        RECT 2491.460 1.820 2495.340 2.700 ;
        RECT 2497.060 1.820 2500.940 2.700 ;
        RECT 2502.660 1.820 2506.540 2.700 ;
        RECT 2508.260 1.820 2512.140 2.700 ;
        RECT 2513.860 1.820 2517.740 2.700 ;
        RECT 2519.460 1.820 2523.340 2.700 ;
        RECT 2525.060 1.820 2528.940 2.700 ;
        RECT 2530.660 1.820 2534.540 2.700 ;
        RECT 2536.260 1.820 2540.140 2.700 ;
        RECT 2541.860 1.820 2545.740 2.700 ;
        RECT 2547.460 1.820 2551.340 2.700 ;
        RECT 2553.060 1.820 2556.940 2.700 ;
        RECT 2558.660 1.820 2562.540 2.700 ;
        RECT 2564.260 1.820 2568.140 2.700 ;
        RECT 2569.860 1.820 2573.740 2.700 ;
        RECT 2575.460 1.820 2579.340 2.700 ;
        RECT 2581.060 1.820 2584.940 2.700 ;
        RECT 2586.660 1.820 2590.540 2.700 ;
        RECT 2592.260 1.820 2596.140 2.700 ;
        RECT 2597.860 1.820 2601.740 2.700 ;
        RECT 2603.460 1.820 2607.340 2.700 ;
        RECT 2609.060 1.820 2612.940 2.700 ;
        RECT 2614.660 1.820 2618.540 2.700 ;
        RECT 2620.260 1.820 2624.140 2.700 ;
        RECT 2625.860 1.820 2629.740 2.700 ;
        RECT 2631.460 1.820 2635.340 2.700 ;
        RECT 2637.060 1.820 2640.940 2.700 ;
        RECT 2642.660 1.820 2646.540 2.700 ;
        RECT 2648.260 1.820 2652.140 2.700 ;
        RECT 2653.860 1.820 2657.740 2.700 ;
        RECT 2659.460 1.820 2663.340 2.700 ;
        RECT 2665.060 1.820 2668.940 2.700 ;
        RECT 2670.660 1.820 2674.540 2.700 ;
        RECT 2676.260 1.820 2680.140 2.700 ;
        RECT 2681.860 1.820 2685.740 2.700 ;
        RECT 2687.460 1.820 2691.340 2.700 ;
        RECT 2693.060 1.820 2696.940 2.700 ;
        RECT 2698.660 1.820 2702.540 2.700 ;
        RECT 2704.260 1.820 2708.140 2.700 ;
        RECT 2709.860 1.820 2713.740 2.700 ;
        RECT 2715.460 1.820 2719.340 2.700 ;
        RECT 2721.060 1.820 2724.940 2.700 ;
        RECT 2726.660 1.820 2730.540 2.700 ;
        RECT 2732.260 1.820 2736.140 2.700 ;
        RECT 2737.860 1.820 2741.740 2.700 ;
        RECT 2743.460 1.820 2747.340 2.700 ;
        RECT 2749.060 1.820 2752.940 2.700 ;
        RECT 2754.660 1.820 2758.540 2.700 ;
        RECT 2760.260 1.820 2764.140 2.700 ;
        RECT 2765.860 1.820 2769.740 2.700 ;
        RECT 2771.460 1.820 2775.340 2.700 ;
        RECT 2777.060 1.820 2780.940 2.700 ;
        RECT 2782.660 1.820 2786.540 2.700 ;
        RECT 2788.260 1.820 2792.140 2.700 ;
        RECT 2793.860 1.820 2797.740 2.700 ;
        RECT 2799.460 1.820 2803.340 2.700 ;
        RECT 2805.060 1.820 2808.940 2.700 ;
        RECT 2810.660 1.820 2814.540 2.700 ;
        RECT 2816.260 1.820 2820.140 2.700 ;
        RECT 2821.860 1.820 2825.740 2.700 ;
        RECT 2827.460 1.820 2831.340 2.700 ;
        RECT 2833.060 1.820 2836.940 2.700 ;
        RECT 2838.660 1.820 2842.540 2.700 ;
        RECT 2844.260 1.820 2848.140 2.700 ;
        RECT 2849.860 1.820 2853.740 2.700 ;
        RECT 2855.460 1.820 2859.340 2.700 ;
        RECT 2861.060 1.820 2950.500 2.700 ;
      LAYER Metal3 ;
        RECT 0.090 2922.100 2958.340 2939.860 ;
        RECT 0.090 2920.420 2957.500 2922.100 ;
        RECT 2.700 2920.380 2957.500 2920.420 ;
        RECT 2.700 2918.700 2958.340 2920.380 ;
        RECT 0.090 2866.660 2958.340 2918.700 ;
        RECT 0.090 2866.100 2957.500 2866.660 ;
        RECT 2.700 2864.940 2957.500 2866.100 ;
        RECT 2.700 2864.380 2958.340 2864.940 ;
        RECT 0.090 2811.780 2958.340 2864.380 ;
        RECT 2.700 2811.220 2958.340 2811.780 ;
        RECT 2.700 2810.060 2957.500 2811.220 ;
        RECT 0.090 2809.500 2957.500 2810.060 ;
        RECT 0.090 2757.460 2958.340 2809.500 ;
        RECT 2.700 2755.780 2958.340 2757.460 ;
        RECT 2.700 2755.740 2957.500 2755.780 ;
        RECT 0.090 2754.060 2957.500 2755.740 ;
        RECT 0.090 2703.140 2958.340 2754.060 ;
        RECT 2.700 2701.420 2958.340 2703.140 ;
        RECT 0.090 2700.340 2958.340 2701.420 ;
        RECT 0.090 2698.620 2957.500 2700.340 ;
        RECT 0.090 2648.820 2958.340 2698.620 ;
        RECT 2.700 2647.100 2958.340 2648.820 ;
        RECT 0.090 2644.900 2958.340 2647.100 ;
        RECT 0.090 2643.180 2957.500 2644.900 ;
        RECT 0.090 2594.500 2958.340 2643.180 ;
        RECT 2.700 2592.780 2958.340 2594.500 ;
        RECT 0.090 2589.460 2958.340 2592.780 ;
        RECT 0.090 2587.740 2957.500 2589.460 ;
        RECT 0.090 2540.180 2958.340 2587.740 ;
        RECT 2.700 2538.460 2958.340 2540.180 ;
        RECT 0.090 2534.020 2958.340 2538.460 ;
        RECT 0.090 2532.300 2957.500 2534.020 ;
        RECT 0.090 2485.860 2958.340 2532.300 ;
        RECT 2.700 2484.140 2958.340 2485.860 ;
        RECT 0.090 2478.580 2958.340 2484.140 ;
        RECT 0.090 2476.860 2957.500 2478.580 ;
        RECT 0.090 2431.540 2958.340 2476.860 ;
        RECT 2.700 2429.820 2958.340 2431.540 ;
        RECT 0.090 2423.140 2958.340 2429.820 ;
        RECT 0.090 2421.420 2957.500 2423.140 ;
        RECT 0.090 2377.220 2958.340 2421.420 ;
        RECT 2.700 2375.500 2958.340 2377.220 ;
        RECT 0.090 2367.700 2958.340 2375.500 ;
        RECT 0.090 2365.980 2957.500 2367.700 ;
        RECT 0.090 2322.900 2958.340 2365.980 ;
        RECT 2.700 2321.180 2958.340 2322.900 ;
        RECT 0.090 2312.260 2958.340 2321.180 ;
        RECT 0.090 2310.540 2957.500 2312.260 ;
        RECT 0.090 2268.580 2958.340 2310.540 ;
        RECT 2.700 2266.860 2958.340 2268.580 ;
        RECT 0.090 2256.820 2958.340 2266.860 ;
        RECT 0.090 2255.100 2957.500 2256.820 ;
        RECT 0.090 2214.260 2958.340 2255.100 ;
        RECT 2.700 2212.540 2958.340 2214.260 ;
        RECT 0.090 2201.380 2958.340 2212.540 ;
        RECT 0.090 2199.660 2957.500 2201.380 ;
        RECT 0.090 2159.940 2958.340 2199.660 ;
        RECT 2.700 2158.220 2958.340 2159.940 ;
        RECT 0.090 2145.940 2958.340 2158.220 ;
        RECT 0.090 2144.220 2957.500 2145.940 ;
        RECT 0.090 2105.620 2958.340 2144.220 ;
        RECT 2.700 2103.900 2958.340 2105.620 ;
        RECT 0.090 2090.500 2958.340 2103.900 ;
        RECT 0.090 2088.780 2957.500 2090.500 ;
        RECT 0.090 2051.300 2958.340 2088.780 ;
        RECT 2.700 2049.580 2958.340 2051.300 ;
        RECT 0.090 2035.060 2958.340 2049.580 ;
        RECT 0.090 2033.340 2957.500 2035.060 ;
        RECT 0.090 1996.980 2958.340 2033.340 ;
        RECT 2.700 1995.260 2958.340 1996.980 ;
        RECT 0.090 1979.620 2958.340 1995.260 ;
        RECT 0.090 1977.900 2957.500 1979.620 ;
        RECT 0.090 1942.660 2958.340 1977.900 ;
        RECT 2.700 1940.940 2958.340 1942.660 ;
        RECT 0.090 1924.180 2958.340 1940.940 ;
        RECT 0.090 1922.460 2957.500 1924.180 ;
        RECT 0.090 1888.340 2958.340 1922.460 ;
        RECT 2.700 1886.620 2958.340 1888.340 ;
        RECT 0.090 1868.740 2958.340 1886.620 ;
        RECT 0.090 1867.020 2957.500 1868.740 ;
        RECT 0.090 1834.020 2958.340 1867.020 ;
        RECT 2.700 1832.300 2958.340 1834.020 ;
        RECT 0.090 1813.300 2958.340 1832.300 ;
        RECT 0.090 1811.580 2957.500 1813.300 ;
        RECT 0.090 1779.700 2958.340 1811.580 ;
        RECT 2.700 1777.980 2958.340 1779.700 ;
        RECT 0.090 1757.860 2958.340 1777.980 ;
        RECT 0.090 1756.140 2957.500 1757.860 ;
        RECT 0.090 1725.380 2958.340 1756.140 ;
        RECT 2.700 1723.660 2958.340 1725.380 ;
        RECT 0.090 1702.420 2958.340 1723.660 ;
        RECT 0.090 1700.700 2957.500 1702.420 ;
        RECT 0.090 1671.060 2958.340 1700.700 ;
        RECT 2.700 1669.340 2958.340 1671.060 ;
        RECT 0.090 1646.980 2958.340 1669.340 ;
        RECT 0.090 1645.260 2957.500 1646.980 ;
        RECT 0.090 1616.740 2958.340 1645.260 ;
        RECT 2.700 1615.020 2958.340 1616.740 ;
        RECT 0.090 1591.540 2958.340 1615.020 ;
        RECT 0.090 1589.820 2957.500 1591.540 ;
        RECT 0.090 1562.420 2958.340 1589.820 ;
        RECT 2.700 1560.700 2958.340 1562.420 ;
        RECT 0.090 1536.100 2958.340 1560.700 ;
        RECT 0.090 1534.380 2957.500 1536.100 ;
        RECT 0.090 1508.100 2958.340 1534.380 ;
        RECT 2.700 1506.380 2958.340 1508.100 ;
        RECT 0.090 1480.660 2958.340 1506.380 ;
        RECT 0.090 1478.940 2957.500 1480.660 ;
        RECT 0.090 1453.780 2958.340 1478.940 ;
        RECT 2.700 1452.060 2958.340 1453.780 ;
        RECT 0.090 1425.220 2958.340 1452.060 ;
        RECT 0.090 1423.500 2957.500 1425.220 ;
        RECT 0.090 1399.460 2958.340 1423.500 ;
        RECT 2.700 1397.740 2958.340 1399.460 ;
        RECT 0.090 1369.780 2958.340 1397.740 ;
        RECT 0.090 1368.060 2957.500 1369.780 ;
        RECT 0.090 1345.140 2958.340 1368.060 ;
        RECT 2.700 1343.420 2958.340 1345.140 ;
        RECT 0.090 1314.340 2958.340 1343.420 ;
        RECT 0.090 1312.620 2957.500 1314.340 ;
        RECT 0.090 1290.820 2958.340 1312.620 ;
        RECT 2.700 1289.100 2958.340 1290.820 ;
        RECT 0.090 1258.900 2958.340 1289.100 ;
        RECT 0.090 1257.180 2957.500 1258.900 ;
        RECT 0.090 1236.500 2958.340 1257.180 ;
        RECT 2.700 1234.780 2958.340 1236.500 ;
        RECT 0.090 1203.460 2958.340 1234.780 ;
        RECT 0.090 1201.740 2957.500 1203.460 ;
        RECT 0.090 1182.180 2958.340 1201.740 ;
        RECT 2.700 1180.460 2958.340 1182.180 ;
        RECT 0.090 1148.020 2958.340 1180.460 ;
        RECT 0.090 1146.300 2957.500 1148.020 ;
        RECT 0.090 1127.860 2958.340 1146.300 ;
        RECT 2.700 1126.140 2958.340 1127.860 ;
        RECT 0.090 1092.580 2958.340 1126.140 ;
        RECT 0.090 1090.860 2957.500 1092.580 ;
        RECT 0.090 1073.540 2958.340 1090.860 ;
        RECT 2.700 1071.820 2958.340 1073.540 ;
        RECT 0.090 1037.140 2958.340 1071.820 ;
        RECT 0.090 1035.420 2957.500 1037.140 ;
        RECT 0.090 1019.220 2958.340 1035.420 ;
        RECT 2.700 1017.500 2958.340 1019.220 ;
        RECT 0.090 981.700 2958.340 1017.500 ;
        RECT 0.090 979.980 2957.500 981.700 ;
        RECT 0.090 964.900 2958.340 979.980 ;
        RECT 2.700 963.180 2958.340 964.900 ;
        RECT 0.090 926.260 2958.340 963.180 ;
        RECT 0.090 924.540 2957.500 926.260 ;
        RECT 0.090 910.580 2958.340 924.540 ;
        RECT 2.700 908.860 2958.340 910.580 ;
        RECT 0.090 870.820 2958.340 908.860 ;
        RECT 0.090 869.100 2957.500 870.820 ;
        RECT 0.090 856.260 2958.340 869.100 ;
        RECT 2.700 854.540 2958.340 856.260 ;
        RECT 0.090 815.380 2958.340 854.540 ;
        RECT 0.090 813.660 2957.500 815.380 ;
        RECT 0.090 801.940 2958.340 813.660 ;
        RECT 2.700 800.220 2958.340 801.940 ;
        RECT 0.090 759.940 2958.340 800.220 ;
        RECT 0.090 758.220 2957.500 759.940 ;
        RECT 0.090 747.620 2958.340 758.220 ;
        RECT 2.700 745.900 2958.340 747.620 ;
        RECT 0.090 704.500 2958.340 745.900 ;
        RECT 0.090 702.780 2957.500 704.500 ;
        RECT 0.090 693.300 2958.340 702.780 ;
        RECT 2.700 691.580 2958.340 693.300 ;
        RECT 0.090 649.060 2958.340 691.580 ;
        RECT 0.090 647.340 2957.500 649.060 ;
        RECT 0.090 638.980 2958.340 647.340 ;
        RECT 2.700 637.260 2958.340 638.980 ;
        RECT 0.090 593.620 2958.340 637.260 ;
        RECT 0.090 591.900 2957.500 593.620 ;
        RECT 0.090 584.660 2958.340 591.900 ;
        RECT 2.700 582.940 2958.340 584.660 ;
        RECT 0.090 538.180 2958.340 582.940 ;
        RECT 0.090 536.460 2957.500 538.180 ;
        RECT 0.090 530.340 2958.340 536.460 ;
        RECT 2.700 528.620 2958.340 530.340 ;
        RECT 0.090 482.740 2958.340 528.620 ;
        RECT 0.090 481.020 2957.500 482.740 ;
        RECT 0.090 476.020 2958.340 481.020 ;
        RECT 2.700 474.300 2958.340 476.020 ;
        RECT 0.090 427.300 2958.340 474.300 ;
        RECT 0.090 425.580 2957.500 427.300 ;
        RECT 0.090 421.700 2958.340 425.580 ;
        RECT 2.700 419.980 2958.340 421.700 ;
        RECT 0.090 371.860 2958.340 419.980 ;
        RECT 0.090 370.140 2957.500 371.860 ;
        RECT 0.090 367.380 2958.340 370.140 ;
        RECT 2.700 365.660 2958.340 367.380 ;
        RECT 0.090 316.420 2958.340 365.660 ;
        RECT 0.090 314.700 2957.500 316.420 ;
        RECT 0.090 313.060 2958.340 314.700 ;
        RECT 2.700 311.340 2958.340 313.060 ;
        RECT 0.090 260.980 2958.340 311.340 ;
        RECT 0.090 259.260 2957.500 260.980 ;
        RECT 0.090 258.740 2958.340 259.260 ;
        RECT 2.700 257.020 2958.340 258.740 ;
        RECT 0.090 205.540 2958.340 257.020 ;
        RECT 0.090 204.420 2957.500 205.540 ;
        RECT 2.700 203.820 2957.500 204.420 ;
        RECT 2.700 202.700 2958.340 203.820 ;
        RECT 0.090 150.100 2958.340 202.700 ;
        RECT 2.700 148.380 2957.500 150.100 ;
        RECT 0.090 95.780 2958.340 148.380 ;
        RECT 2.700 94.660 2958.340 95.780 ;
        RECT 2.700 94.060 2957.500 94.660 ;
        RECT 0.090 92.940 2957.500 94.060 ;
        RECT 0.090 41.460 2958.340 92.940 ;
        RECT 2.700 39.740 2958.340 41.460 ;
        RECT 0.090 39.220 2958.340 39.740 ;
        RECT 0.090 37.500 2957.500 39.220 ;
        RECT 0.090 3.500 2958.340 37.500 ;
      LAYER Metal4 ;
        RECT 38.220 2291.410 105.470 2939.910 ;
        RECT 109.170 2291.410 124.070 2939.910 ;
        RECT 127.770 2291.410 195.470 2939.910 ;
        RECT 199.170 2291.410 214.070 2939.910 ;
        RECT 217.770 2291.410 285.470 2939.910 ;
        RECT 289.170 2291.410 304.070 2939.910 ;
        RECT 307.770 2291.410 375.470 2939.910 ;
        RECT 379.170 2291.410 394.070 2939.910 ;
        RECT 397.770 2291.410 465.470 2939.910 ;
        RECT 469.170 2291.410 484.070 2939.910 ;
        RECT 487.770 2291.410 555.470 2939.910 ;
        RECT 559.170 2291.410 574.070 2939.910 ;
        RECT 577.770 2291.410 645.470 2939.910 ;
        RECT 649.170 2291.410 664.070 2939.910 ;
        RECT 667.770 2291.410 735.470 2939.910 ;
        RECT 739.170 2291.410 754.070 2939.910 ;
        RECT 757.770 2291.410 825.470 2939.910 ;
        RECT 829.170 2291.410 844.070 2939.910 ;
        RECT 847.770 2291.410 915.470 2939.910 ;
        RECT 919.170 2291.410 934.070 2939.910 ;
        RECT 937.770 2291.410 1005.470 2939.910 ;
        RECT 38.220 1594.590 1005.470 2291.410 ;
        RECT 38.220 1491.410 124.070 1594.590 ;
        RECT 127.770 1491.410 214.070 1594.590 ;
        RECT 217.770 1491.410 304.070 1594.590 ;
        RECT 307.770 1491.410 394.070 1594.590 ;
        RECT 397.770 1491.410 484.070 1594.590 ;
        RECT 487.770 1491.410 574.070 1594.590 ;
        RECT 577.770 1491.410 664.070 1594.590 ;
        RECT 667.770 1491.410 754.070 1594.590 ;
        RECT 757.770 1491.410 844.070 1594.590 ;
        RECT 847.770 1491.410 934.070 1594.590 ;
        RECT 937.770 1491.410 1005.470 1594.590 ;
        RECT 38.220 794.590 1005.470 1491.410 ;
        RECT 38.220 3.450 105.470 794.590 ;
        RECT 109.170 3.450 124.070 794.590 ;
        RECT 127.770 3.450 195.470 794.590 ;
        RECT 199.170 3.450 214.070 794.590 ;
        RECT 217.770 555.890 285.470 794.590 ;
        RECT 289.170 555.890 304.070 794.590 ;
        RECT 307.770 555.890 375.470 794.590 ;
        RECT 379.170 555.890 394.070 794.590 ;
        RECT 397.770 555.890 465.470 794.590 ;
        RECT 469.170 555.890 484.070 794.590 ;
        RECT 487.770 555.890 555.470 794.590 ;
        RECT 559.170 555.890 574.070 794.590 ;
        RECT 577.770 555.890 645.470 794.590 ;
        RECT 649.170 555.890 664.070 794.590 ;
        RECT 667.770 555.890 735.470 794.590 ;
        RECT 739.170 555.890 754.070 794.590 ;
        RECT 757.770 555.890 825.470 794.590 ;
        RECT 829.170 555.890 844.070 794.590 ;
        RECT 847.770 555.890 915.470 794.590 ;
        RECT 217.770 388.270 915.470 555.890 ;
        RECT 217.770 3.450 285.470 388.270 ;
        RECT 289.170 3.450 304.070 388.270 ;
        RECT 307.770 3.450 375.470 388.270 ;
        RECT 379.170 3.450 394.070 388.270 ;
        RECT 397.770 3.450 465.470 388.270 ;
        RECT 469.170 3.450 484.070 388.270 ;
        RECT 487.770 3.450 555.470 388.270 ;
        RECT 559.170 3.450 574.070 388.270 ;
        RECT 577.770 3.450 645.470 388.270 ;
        RECT 649.170 3.450 664.070 388.270 ;
        RECT 667.770 3.450 735.470 388.270 ;
        RECT 739.170 3.450 754.070 388.270 ;
        RECT 757.770 3.450 825.470 388.270 ;
        RECT 829.170 3.450 844.070 388.270 ;
        RECT 847.770 3.450 915.470 388.270 ;
        RECT 919.170 3.450 934.070 794.590 ;
        RECT 937.770 3.450 1005.470 794.590 ;
        RECT 1009.170 3.450 1024.070 2939.910 ;
        RECT 1027.770 2291.410 1095.470 2939.910 ;
        RECT 1099.170 2291.410 1114.070 2939.910 ;
        RECT 1117.770 2291.410 1185.470 2939.910 ;
        RECT 1189.170 2291.410 1204.070 2939.910 ;
        RECT 1207.770 2291.410 1275.470 2939.910 ;
        RECT 1279.170 2291.410 1294.070 2939.910 ;
        RECT 1297.770 2291.410 1365.470 2939.910 ;
        RECT 1369.170 2291.410 1384.070 2939.910 ;
        RECT 1387.770 2291.410 1455.470 2939.910 ;
        RECT 1459.170 2291.410 1474.070 2939.910 ;
        RECT 1477.770 2291.410 1545.470 2939.910 ;
        RECT 1549.170 2291.410 1564.070 2939.910 ;
        RECT 1567.770 2291.410 1635.470 2939.910 ;
        RECT 1639.170 2291.410 1654.070 2939.910 ;
        RECT 1657.770 2291.410 1725.470 2939.910 ;
        RECT 1729.170 2291.410 1744.070 2939.910 ;
        RECT 1747.770 2291.410 1815.470 2939.910 ;
        RECT 1819.170 2291.410 1834.070 2939.910 ;
        RECT 1837.770 2291.410 1905.470 2939.910 ;
        RECT 1027.770 1594.590 1905.470 2291.410 ;
        RECT 1027.770 1491.410 1114.070 1594.590 ;
        RECT 1117.770 1491.410 1204.070 1594.590 ;
        RECT 1207.770 1491.410 1294.070 1594.590 ;
        RECT 1297.770 1491.410 1384.070 1594.590 ;
        RECT 1387.770 1491.410 1474.070 1594.590 ;
        RECT 1477.770 1491.410 1564.070 1594.590 ;
        RECT 1567.770 1491.410 1654.070 1594.590 ;
        RECT 1657.770 1491.410 1744.070 1594.590 ;
        RECT 1747.770 1491.410 1834.070 1594.590 ;
        RECT 1837.770 1491.410 1905.470 1594.590 ;
        RECT 1027.770 794.590 1905.470 1491.410 ;
        RECT 1027.770 741.410 1095.470 794.590 ;
        RECT 1099.170 741.410 1114.070 794.590 ;
        RECT 1117.770 741.410 1185.470 794.590 ;
        RECT 1189.170 741.410 1204.070 794.590 ;
        RECT 1207.770 741.410 1275.470 794.590 ;
        RECT 1279.170 741.410 1294.070 794.590 ;
        RECT 1297.770 741.410 1365.470 794.590 ;
        RECT 1369.170 741.410 1384.070 794.590 ;
        RECT 1387.770 741.410 1455.470 794.590 ;
        RECT 1459.170 741.410 1474.070 794.590 ;
        RECT 1477.770 741.410 1545.470 794.590 ;
        RECT 1549.170 741.410 1564.070 794.590 ;
        RECT 1567.770 741.410 1635.470 794.590 ;
        RECT 1639.170 741.410 1654.070 794.590 ;
        RECT 1657.770 741.410 1725.470 794.590 ;
        RECT 1729.170 741.410 1744.070 794.590 ;
        RECT 1747.770 741.410 1815.470 794.590 ;
        RECT 1819.170 741.410 1834.070 794.590 ;
        RECT 1837.770 741.410 1905.470 794.590 ;
        RECT 1027.770 44.590 1905.470 741.410 ;
        RECT 1027.770 3.450 1095.470 44.590 ;
        RECT 1099.170 3.450 1185.470 44.590 ;
        RECT 1189.170 3.450 1275.470 44.590 ;
        RECT 1279.170 3.450 1365.470 44.590 ;
        RECT 1369.170 3.450 1455.470 44.590 ;
        RECT 1459.170 3.450 1545.470 44.590 ;
        RECT 1549.170 3.450 1635.470 44.590 ;
        RECT 1639.170 3.450 1725.470 44.590 ;
        RECT 1729.170 3.450 1815.470 44.590 ;
        RECT 1819.170 3.450 1905.470 44.590 ;
        RECT 1909.170 3.450 1924.070 2939.910 ;
        RECT 1927.770 3.450 1995.470 2939.910 ;
        RECT 1999.170 3.450 2014.070 2939.910 ;
        RECT 2017.770 2291.410 2085.470 2939.910 ;
        RECT 2089.170 2291.410 2104.070 2939.910 ;
        RECT 2107.770 2291.410 2175.470 2939.910 ;
        RECT 2179.170 2291.410 2194.070 2939.910 ;
        RECT 2197.770 2291.410 2265.470 2939.910 ;
        RECT 2269.170 2291.410 2284.070 2939.910 ;
        RECT 2287.770 2291.410 2355.470 2939.910 ;
        RECT 2359.170 2291.410 2374.070 2939.910 ;
        RECT 2377.770 2291.410 2445.470 2939.910 ;
        RECT 2449.170 2291.410 2464.070 2939.910 ;
        RECT 2467.770 2291.410 2535.470 2939.910 ;
        RECT 2539.170 2291.410 2554.070 2939.910 ;
        RECT 2557.770 2291.410 2625.470 2939.910 ;
        RECT 2629.170 2291.410 2644.070 2939.910 ;
        RECT 2647.770 2291.410 2715.470 2939.910 ;
        RECT 2719.170 2291.410 2734.070 2939.910 ;
        RECT 2737.770 2291.410 2805.470 2939.910 ;
        RECT 2809.170 2291.410 2824.070 2939.910 ;
        RECT 2827.770 2291.410 2879.660 2939.910 ;
        RECT 2017.770 1594.590 2879.660 2291.410 ;
        RECT 2017.770 1491.410 2104.070 1594.590 ;
        RECT 2107.770 1491.410 2194.070 1594.590 ;
        RECT 2197.770 1491.410 2284.070 1594.590 ;
        RECT 2287.770 1491.410 2374.070 1594.590 ;
        RECT 2377.770 1491.410 2464.070 1594.590 ;
        RECT 2467.770 1491.410 2554.070 1594.590 ;
        RECT 2557.770 1491.410 2644.070 1594.590 ;
        RECT 2647.770 1491.410 2734.070 1594.590 ;
        RECT 2737.770 1491.410 2824.070 1594.590 ;
        RECT 2827.770 1491.410 2879.660 1594.590 ;
        RECT 2017.770 794.590 2879.660 1491.410 ;
        RECT 2017.770 3.450 2085.470 794.590 ;
        RECT 2089.170 3.450 2104.070 794.590 ;
        RECT 2107.770 3.450 2175.470 794.590 ;
        RECT 2179.170 3.450 2194.070 794.590 ;
        RECT 2197.770 3.450 2265.470 794.590 ;
        RECT 2269.170 3.450 2284.070 794.590 ;
        RECT 2287.770 3.450 2355.470 794.590 ;
        RECT 2359.170 3.450 2374.070 794.590 ;
        RECT 2377.770 3.450 2445.470 794.590 ;
        RECT 2449.170 3.450 2464.070 794.590 ;
        RECT 2467.770 3.450 2535.470 794.590 ;
        RECT 2539.170 3.450 2554.070 794.590 ;
        RECT 2557.770 3.450 2625.470 794.590 ;
        RECT 2629.170 3.450 2644.070 794.590 ;
        RECT 2647.770 3.450 2715.470 794.590 ;
        RECT 2719.170 3.450 2734.070 794.590 ;
        RECT 2737.770 3.450 2805.470 794.590 ;
        RECT 2809.170 3.450 2824.070 794.590 ;
        RECT 2827.770 3.450 2879.660 794.590 ;
  END
END user_project_wrapper
END LIBRARY

